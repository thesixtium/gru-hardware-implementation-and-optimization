`timescale 1ns / 1ps

module gru_tb;

// Parameters
parameter int D          = 64;
parameter int H          = 16;
parameter int DATA_WIDTH = 11;
parameter int FRAC_BITS  = 5;
parameter int NUM_PARALLEL = 1;
parameter real CLK_PERIOD = 10.0;

// Clock and reset
logic clk;
logic rst_n;
logic start;
logic done;

// Cycle counter
int cycle_count = 0;
int test_start_cycle = 0;
int test_cycles = 0;
int total_cycles = 0;
bit test_timeout = 0;

// Input arrays
logic signed [DATA_WIDTH-1:0] x_t [D-1:0];
logic signed [DATA_WIDTH-1:0] h_t_prev [H-1:0];
logic signed [DATA_WIDTH-1:0] h_t [H-1:0];

// Weight matrices
logic signed [DATA_WIDTH-1:0] W_ir [H-1:0][D-1:0];
logic signed [DATA_WIDTH-1:0] W_hr [H-1:0][H-1:0];
logic signed [DATA_WIDTH-1:0] b_ir [H-1:0];
logic signed [DATA_WIDTH-1:0] b_hr [H-1:0];

logic signed [DATA_WIDTH-1:0] W_iz [H-1:0][D-1:0];
logic signed [DATA_WIDTH-1:0] W_hz [H-1:0][H-1:0];
logic signed [DATA_WIDTH-1:0] b_iz [H-1:0];
logic signed [DATA_WIDTH-1:0] b_hz [H-1:0];

logic signed [DATA_WIDTH-1:0] W_in [H-1:0][D-1:0];
logic signed [DATA_WIDTH-1:0] W_hn [H-1:0][H-1:0];
logic signed [DATA_WIDTH-1:0] b_in [H-1:0];
logic signed [DATA_WIDTH-1:0] b_hn [H-1:0];

// DUT instantiation
gru_cell_parallel #(
    .D(D),
    .H(H),
    .DATA_WIDTH(DATA_WIDTH),
    .FRAC_BITS(FRAC_BITS),
    .NUM_PARALLEL(NUM_PARALLEL)
) dut (
    .clk(clk),
    .rst_n(rst_n),
    .start(start),
    .x_t(x_t),
    .h_t_prev(h_t_prev),
    .W_ir(W_ir),
    .W_hr(W_hr),
    .b_ir(b_ir),
    .b_hr(b_hr),
    .W_iz(W_iz),
    .W_hz(W_hz),
    .b_iz(b_iz),
    .b_hz(b_hz),
    .W_in(W_in),
    .W_hn(W_hn),
    .b_in(b_in),
    .b_hn(b_hn),
    .h_t(h_t),
    .done(done)
);

// Clock generation
initial begin
    clk = 0;
    forever #5 clk = ~clk; // 100MHz clock
end

// Cycle counter
always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        cycle_count <= 0;
    end else begin
        cycle_count <= cycle_count + 1;
    end
end

initial begin
    // Open files for writing
    integer fd_output;
    integer fd_cycles;
    
    fd_output = $fopen("../../../../../output_d64_h16_dw11_fb5_np1.txt", "w+");
    if (fd_output == 0) begin
        $display("ERROR: Failed to open output file!");
        $finish;
    end
    
    fd_cycles = $fopen("../../../../../cycles_d64_h16_dw11_fb5_np1.txt", "w+");
    if (fd_cycles == 0) begin
        $display("ERROR: Failed to open cycles file!");
        $fclose(fd_output);
        $finish;
    end
    
    // Write header to cycles file
    $fdisplay(fd_cycles, "==========================================================");
    $fdisplay(fd_cycles, "GRU Cell Parallel Cycle Count Results");
    $fdisplay(fd_cycles, "==========================================================");
    $fdisplay(fd_cycles, "Parameters:");
    $fdisplay(fd_cycles, "  D (Input Dimension):     64");
    $fdisplay(fd_cycles, "  H (Hidden Dimension):    16");
    $fdisplay(fd_cycles, "  DATA_WIDTH:              11");
    $fdisplay(fd_cycles, "  FRAC_BITS:               5");
    $fdisplay(fd_cycles, "  NUM_PARALLEL:            1");
    $fdisplay(fd_cycles, "  Total Test Vectors:      100");
    $fdisplay(fd_cycles, "==========================================================");
    $fdisplay(fd_cycles, "");
    
    // Initialize weights
    // Initialize W_ir weights
    W_ir[0][0] = 11'b00000000011;
    W_ir[0][1] = 11'b00000000101;
    W_ir[0][2] = 11'b00000000100;
    W_ir[0][3] = 11'b00000000100;
    W_ir[0][4] = 11'b11111111110;
    W_ir[0][5] = 11'b11111111011;
    W_ir[0][6] = 11'b00000000100;
    W_ir[0][7] = 11'b00000000010;
    W_ir[0][8] = 11'b11111111001;
    W_ir[0][9] = 11'b00000000001;
    W_ir[0][10] = 11'b00000001000;
    W_ir[0][11] = 11'b00000000000;
    W_ir[0][12] = 11'b00000000101;
    W_ir[0][13] = 11'b00000000001;
    W_ir[0][14] = 11'b00000000001;
    W_ir[0][15] = 11'b00000000110;
    W_ir[0][16] = 11'b11111111111;
    W_ir[0][17] = 11'b00000000111;
    W_ir[0][18] = 11'b11111111111;
    W_ir[0][19] = 11'b00000000101;
    W_ir[0][20] = 11'b11111111111;
    W_ir[0][21] = 11'b00000000100;
    W_ir[0][22] = 11'b00000000011;
    W_ir[0][23] = 11'b00000000011;
    W_ir[0][24] = 11'b11111111011;
    W_ir[0][25] = 11'b00000000100;
    W_ir[0][26] = 11'b00000000100;
    W_ir[0][27] = 11'b00000000011;
    W_ir[0][28] = 11'b00000000111;
    W_ir[0][29] = 11'b11111111001;
    W_ir[0][30] = 11'b11111111110;
    W_ir[0][31] = 11'b00000000011;
    W_ir[0][32] = 11'b00000000010;
    W_ir[0][33] = 11'b00000000100;
    W_ir[0][34] = 11'b00000000100;
    W_ir[0][35] = 11'b00000000001;
    W_ir[0][36] = 11'b00000001000;
    W_ir[0][37] = 11'b00000000011;
    W_ir[0][38] = 11'b11111111110;
    W_ir[0][39] = 11'b00000000010;
    W_ir[0][40] = 11'b00000000101;
    W_ir[0][41] = 11'b11111111010;
    W_ir[0][42] = 11'b00000000010;
    W_ir[0][43] = 11'b11111111101;
    W_ir[0][44] = 11'b00000000000;
    W_ir[0][45] = 11'b11111111100;
    W_ir[0][46] = 11'b11111111010;
    W_ir[0][47] = 11'b00000000111;
    W_ir[0][48] = 11'b11111111110;
    W_ir[0][49] = 11'b11111111101;
    W_ir[0][50] = 11'b11111111111;
    W_ir[0][51] = 11'b00000000000;
    W_ir[0][52] = 11'b11111111001;
    W_ir[0][53] = 11'b11111111101;
    W_ir[0][54] = 11'b00000000010;
    W_ir[0][55] = 11'b11111111101;
    W_ir[0][56] = 11'b00000000101;
    W_ir[0][57] = 11'b11111111101;
    W_ir[0][58] = 11'b11111111101;
    W_ir[0][59] = 11'b00000000100;
    W_ir[0][60] = 11'b11111111011;
    W_ir[0][61] = 11'b11111111010;
    W_ir[0][62] = 11'b11111111010;
    W_ir[0][63] = 11'b00000000100;
    W_ir[1][0] = 11'b11111111100;
    W_ir[1][1] = 11'b11111111101;
    W_ir[1][2] = 11'b00000000110;
    W_ir[1][3] = 11'b00000000101;
    W_ir[1][4] = 11'b00000000001;
    W_ir[1][5] = 11'b00000000010;
    W_ir[1][6] = 11'b00000000010;
    W_ir[1][7] = 11'b00000000001;
    W_ir[1][8] = 11'b00000000001;
    W_ir[1][9] = 11'b00000000001;
    W_ir[1][10] = 11'b11111111111;
    W_ir[1][11] = 11'b00000000000;
    W_ir[1][12] = 11'b00000000001;
    W_ir[1][13] = 11'b00000000100;
    W_ir[1][14] = 11'b11111111011;
    W_ir[1][15] = 11'b00000000001;
    W_ir[1][16] = 11'b00000000000;
    W_ir[1][17] = 11'b00000000000;
    W_ir[1][18] = 11'b00000000000;
    W_ir[1][19] = 11'b11111111101;
    W_ir[1][20] = 11'b00000000000;
    W_ir[1][21] = 11'b00000000001;
    W_ir[1][22] = 11'b11111111110;
    W_ir[1][23] = 11'b11111111101;
    W_ir[1][24] = 11'b00000000000;
    W_ir[1][25] = 11'b00000000110;
    W_ir[1][26] = 11'b11111111010;
    W_ir[1][27] = 11'b11111111010;
    W_ir[1][28] = 11'b00000000111;
    W_ir[1][29] = 11'b00000000010;
    W_ir[1][30] = 11'b00000000000;
    W_ir[1][31] = 11'b00000000000;
    W_ir[1][32] = 11'b11111111100;
    W_ir[1][33] = 11'b00000000000;
    W_ir[1][34] = 11'b11111111111;
    W_ir[1][35] = 11'b00000000000;
    W_ir[1][36] = 11'b00000000010;
    W_ir[1][37] = 11'b00000000001;
    W_ir[1][38] = 11'b00000000010;
    W_ir[1][39] = 11'b00000000100;
    W_ir[1][40] = 11'b00000000010;
    W_ir[1][41] = 11'b00000000000;
    W_ir[1][42] = 11'b00000000000;
    W_ir[1][43] = 11'b00000000010;
    W_ir[1][44] = 11'b00000000001;
    W_ir[1][45] = 11'b00000000010;
    W_ir[1][46] = 11'b00000000000;
    W_ir[1][47] = 11'b11111111111;
    W_ir[1][48] = 11'b11111111111;
    W_ir[1][49] = 11'b11111111001;
    W_ir[1][50] = 11'b00000000100;
    W_ir[1][51] = 11'b00000000101;
    W_ir[1][52] = 11'b11111111110;
    W_ir[1][53] = 11'b11111111101;
    W_ir[1][54] = 11'b11111111101;
    W_ir[1][55] = 11'b11111111101;
    W_ir[1][56] = 11'b11111111110;
    W_ir[1][57] = 11'b00000000110;
    W_ir[1][58] = 11'b00000000100;
    W_ir[1][59] = 11'b11111111100;
    W_ir[1][60] = 11'b11111111111;
    W_ir[1][61] = 11'b11111111110;
    W_ir[1][62] = 11'b00000000101;
    W_ir[1][63] = 11'b11111111101;
    W_ir[2][0] = 11'b11111111101;
    W_ir[2][1] = 11'b11111111110;
    W_ir[2][2] = 11'b11111111001;
    W_ir[2][3] = 11'b11111111100;
    W_ir[2][4] = 11'b11111111110;
    W_ir[2][5] = 11'b11111111111;
    W_ir[2][6] = 11'b00000000001;
    W_ir[2][7] = 11'b11111111011;
    W_ir[2][8] = 11'b11111111111;
    W_ir[2][9] = 11'b11111111111;
    W_ir[2][10] = 11'b11111111111;
    W_ir[2][11] = 11'b11111111001;
    W_ir[2][12] = 11'b11111111111;
    W_ir[2][13] = 11'b00000000010;
    W_ir[2][14] = 11'b11111111111;
    W_ir[2][15] = 11'b00000000011;
    W_ir[2][16] = 11'b11111111011;
    W_ir[2][17] = 11'b00000000111;
    W_ir[2][18] = 11'b00000000000;
    W_ir[2][19] = 11'b00000000010;
    W_ir[2][20] = 11'b00000000010;
    W_ir[2][21] = 11'b11111111110;
    W_ir[2][22] = 11'b00000000100;
    W_ir[2][23] = 11'b00000000111;
    W_ir[2][24] = 11'b00000000011;
    W_ir[2][25] = 11'b00000000001;
    W_ir[2][26] = 11'b00000000000;
    W_ir[2][27] = 11'b11111111001;
    W_ir[2][28] = 11'b11111111110;
    W_ir[2][29] = 11'b00000001000;
    W_ir[2][30] = 11'b11111111101;
    W_ir[2][31] = 11'b11111111101;
    W_ir[2][32] = 11'b00000000000;
    W_ir[2][33] = 11'b00000000011;
    W_ir[2][34] = 11'b11111111111;
    W_ir[2][35] = 11'b11111111110;
    W_ir[2][36] = 11'b00000000000;
    W_ir[2][37] = 11'b00000000001;
    W_ir[2][38] = 11'b00000000100;
    W_ir[2][39] = 11'b00000000000;
    W_ir[2][40] = 11'b00000000100;
    W_ir[2][41] = 11'b11111111110;
    W_ir[2][42] = 11'b00000000100;
    W_ir[2][43] = 11'b00000000000;
    W_ir[2][44] = 11'b00000000001;
    W_ir[2][45] = 11'b00000000010;
    W_ir[2][46] = 11'b00000000010;
    W_ir[2][47] = 11'b00000000001;
    W_ir[2][48] = 11'b00000000010;
    W_ir[2][49] = 11'b00000000001;
    W_ir[2][50] = 11'b11111111100;
    W_ir[2][51] = 11'b00000000011;
    W_ir[2][52] = 11'b00000000011;
    W_ir[2][53] = 11'b00000000010;
    W_ir[2][54] = 11'b11111111001;
    W_ir[2][55] = 11'b00000000010;
    W_ir[2][56] = 11'b00000000010;
    W_ir[2][57] = 11'b11111111011;
    W_ir[2][58] = 11'b11111111100;
    W_ir[2][59] = 11'b11111111101;
    W_ir[2][60] = 11'b00000000101;
    W_ir[2][61] = 11'b00000000010;
    W_ir[2][62] = 11'b00000000101;
    W_ir[2][63] = 11'b00000001001;
    W_ir[3][0] = 11'b00000000000;
    W_ir[3][1] = 11'b00000001000;
    W_ir[3][2] = 11'b00000000000;
    W_ir[3][3] = 11'b00000000110;
    W_ir[3][4] = 11'b11111111010;
    W_ir[3][5] = 11'b00000000001;
    W_ir[3][6] = 11'b00000000001;
    W_ir[3][7] = 11'b11111111110;
    W_ir[3][8] = 11'b11111111111;
    W_ir[3][9] = 11'b00000000101;
    W_ir[3][10] = 11'b11111111100;
    W_ir[3][11] = 11'b11111111111;
    W_ir[3][12] = 11'b11111111100;
    W_ir[3][13] = 11'b11111111111;
    W_ir[3][14] = 11'b11111111110;
    W_ir[3][15] = 11'b11111111111;
    W_ir[3][16] = 11'b00000000000;
    W_ir[3][17] = 11'b00000000001;
    W_ir[3][18] = 11'b11111111101;
    W_ir[3][19] = 11'b00000000100;
    W_ir[3][20] = 11'b11111111110;
    W_ir[3][21] = 11'b00000000010;
    W_ir[3][22] = 11'b00000000011;
    W_ir[3][23] = 11'b00000000010;
    W_ir[3][24] = 11'b00000000111;
    W_ir[3][25] = 11'b00000000001;
    W_ir[3][26] = 11'b11111111111;
    W_ir[3][27] = 11'b11111111110;
    W_ir[3][28] = 11'b00000000001;
    W_ir[3][29] = 11'b00000000001;
    W_ir[3][30] = 11'b11111111100;
    W_ir[3][31] = 11'b00000001000;
    W_ir[3][32] = 11'b00000000100;
    W_ir[3][33] = 11'b11111111011;
    W_ir[3][34] = 11'b00000000010;
    W_ir[3][35] = 11'b00000000001;
    W_ir[3][36] = 11'b00000000001;
    W_ir[3][37] = 11'b11111111001;
    W_ir[3][38] = 11'b00000000011;
    W_ir[3][39] = 11'b00000000000;
    W_ir[3][40] = 11'b00000000000;
    W_ir[3][41] = 11'b00000000101;
    W_ir[3][42] = 11'b11111111011;
    W_ir[3][43] = 11'b00000000001;
    W_ir[3][44] = 11'b11111111101;
    W_ir[3][45] = 11'b11111111110;
    W_ir[3][46] = 11'b00000000110;
    W_ir[3][47] = 11'b11111111101;
    W_ir[3][48] = 11'b11111111110;
    W_ir[3][49] = 11'b11111111111;
    W_ir[3][50] = 11'b11111111100;
    W_ir[3][51] = 11'b11111111101;
    W_ir[3][52] = 11'b11111111101;
    W_ir[3][53] = 11'b11111111100;
    W_ir[3][54] = 11'b11111111110;
    W_ir[3][55] = 11'b11111111001;
    W_ir[3][56] = 11'b11111111101;
    W_ir[3][57] = 11'b00000000100;
    W_ir[3][58] = 11'b11111111100;
    W_ir[3][59] = 11'b11111111101;
    W_ir[3][60] = 11'b11111111101;
    W_ir[3][61] = 11'b11111111101;
    W_ir[3][62] = 11'b11111111010;
    W_ir[3][63] = 11'b11111111110;
    W_ir[4][0] = 11'b00000000000;
    W_ir[4][1] = 11'b11111111110;
    W_ir[4][2] = 11'b11111111111;
    W_ir[4][3] = 11'b11111111101;
    W_ir[4][4] = 11'b00000000000;
    W_ir[4][5] = 11'b00000000011;
    W_ir[4][6] = 11'b11111111100;
    W_ir[4][7] = 11'b11111111011;
    W_ir[4][8] = 11'b11111111001;
    W_ir[4][9] = 11'b11111111101;
    W_ir[4][10] = 11'b11111111001;
    W_ir[4][11] = 11'b11111111110;
    W_ir[4][12] = 11'b11111111111;
    W_ir[4][13] = 11'b00000000011;
    W_ir[4][14] = 11'b00000000001;
    W_ir[4][15] = 11'b11111111111;
    W_ir[4][16] = 11'b11111111100;
    W_ir[4][17] = 11'b11111111101;
    W_ir[4][18] = 11'b11111111100;
    W_ir[4][19] = 11'b11111111011;
    W_ir[4][20] = 11'b11111111111;
    W_ir[4][21] = 11'b00000000011;
    W_ir[4][22] = 11'b00000001000;
    W_ir[4][23] = 11'b00000000101;
    W_ir[4][24] = 11'b11111111001;
    W_ir[4][25] = 11'b11111111010;
    W_ir[4][26] = 11'b00000000000;
    W_ir[4][27] = 11'b11111111001;
    W_ir[4][28] = 11'b00000000110;
    W_ir[4][29] = 11'b00000000000;
    W_ir[4][30] = 11'b00000000110;
    W_ir[4][31] = 11'b11111111100;
    W_ir[4][32] = 11'b11111111001;
    W_ir[4][33] = 11'b11111111010;
    W_ir[4][34] = 11'b11111111100;
    W_ir[4][35] = 11'b11111111100;
    W_ir[4][36] = 11'b11111111010;
    W_ir[4][37] = 11'b11111111011;
    W_ir[4][38] = 11'b11111111101;
    W_ir[4][39] = 11'b00000000010;
    W_ir[4][40] = 11'b00000000001;
    W_ir[4][41] = 11'b11111111100;
    W_ir[4][42] = 11'b11111111111;
    W_ir[4][43] = 11'b11111111101;
    W_ir[4][44] = 11'b11111111000;
    W_ir[4][45] = 11'b11111111111;
    W_ir[4][46] = 11'b11111111111;
    W_ir[4][47] = 11'b11111111111;
    W_ir[4][48] = 11'b00000000000;
    W_ir[4][49] = 11'b11111111110;
    W_ir[4][50] = 11'b00000000101;
    W_ir[4][51] = 11'b11111111101;
    W_ir[4][52] = 11'b00000000111;
    W_ir[4][53] = 11'b00000000100;
    W_ir[4][54] = 11'b00000001000;
    W_ir[4][55] = 11'b00000000110;
    W_ir[4][56] = 11'b00000000011;
    W_ir[4][57] = 11'b11111111001;
    W_ir[4][58] = 11'b00000000100;
    W_ir[4][59] = 11'b00000001110;
    W_ir[4][60] = 11'b00000001010;
    W_ir[4][61] = 11'b00000001011;
    W_ir[4][62] = 11'b00000001101;
    W_ir[4][63] = 11'b00000001100;
    W_ir[5][0] = 11'b00000000001;
    W_ir[5][1] = 11'b00000000001;
    W_ir[5][2] = 11'b00000000010;
    W_ir[5][3] = 11'b11111111111;
    W_ir[5][4] = 11'b11111111111;
    W_ir[5][5] = 11'b11111111011;
    W_ir[5][6] = 11'b00000000110;
    W_ir[5][7] = 11'b11111111001;
    W_ir[5][8] = 11'b11111111010;
    W_ir[5][9] = 11'b11111111110;
    W_ir[5][10] = 11'b00000000000;
    W_ir[5][11] = 11'b11111111111;
    W_ir[5][12] = 11'b11111111100;
    W_ir[5][13] = 11'b11111111111;
    W_ir[5][14] = 11'b11111111100;
    W_ir[5][15] = 11'b11111111100;
    W_ir[5][16] = 11'b00000000101;
    W_ir[5][17] = 11'b11111111011;
    W_ir[5][18] = 11'b00000000001;
    W_ir[5][19] = 11'b11111111010;
    W_ir[5][20] = 11'b11111111111;
    W_ir[5][21] = 11'b00000000000;
    W_ir[5][22] = 11'b00000000011;
    W_ir[5][23] = 11'b00000000010;
    W_ir[5][24] = 11'b11111111111;
    W_ir[5][25] = 11'b11111111101;
    W_ir[5][26] = 11'b11111111111;
    W_ir[5][27] = 11'b00000000011;
    W_ir[5][28] = 11'b00000000001;
    W_ir[5][29] = 11'b11111111100;
    W_ir[5][30] = 11'b11111111110;
    W_ir[5][31] = 11'b11111111001;
    W_ir[5][32] = 11'b00000000000;
    W_ir[5][33] = 11'b11111111000;
    W_ir[5][34] = 11'b11111111110;
    W_ir[5][35] = 11'b00000000100;
    W_ir[5][36] = 11'b11111111100;
    W_ir[5][37] = 11'b11111111010;
    W_ir[5][38] = 11'b11111110111;
    W_ir[5][39] = 11'b00000000101;
    W_ir[5][40] = 11'b11111111101;
    W_ir[5][41] = 11'b11111111111;
    W_ir[5][42] = 11'b00000000000;
    W_ir[5][43] = 11'b11111111101;
    W_ir[5][44] = 11'b00000000001;
    W_ir[5][45] = 11'b11111111101;
    W_ir[5][46] = 11'b11111111111;
    W_ir[5][47] = 11'b00000000100;
    W_ir[5][48] = 11'b00000000010;
    W_ir[5][49] = 11'b00000000010;
    W_ir[5][50] = 11'b00000000001;
    W_ir[5][51] = 11'b00000000001;
    W_ir[5][52] = 11'b11111111110;
    W_ir[5][53] = 11'b11111111101;
    W_ir[5][54] = 11'b00000000010;
    W_ir[5][55] = 11'b00000000000;
    W_ir[5][56] = 11'b00000000001;
    W_ir[5][57] = 11'b11111111011;
    W_ir[5][58] = 11'b11111111100;
    W_ir[5][59] = 11'b11111111110;
    W_ir[5][60] = 11'b00000000111;
    W_ir[5][61] = 11'b00000000101;
    W_ir[5][62] = 11'b11111111110;
    W_ir[5][63] = 11'b00000000101;
    W_ir[6][0] = 11'b00000000110;
    W_ir[6][1] = 11'b11111111110;
    W_ir[6][2] = 11'b00000001001;
    W_ir[6][3] = 11'b11111111110;
    W_ir[6][4] = 11'b00000000101;
    W_ir[6][5] = 11'b00000000001;
    W_ir[6][6] = 11'b11111111001;
    W_ir[6][7] = 11'b00000001001;
    W_ir[6][8] = 11'b00000001011;
    W_ir[6][9] = 11'b00000000110;
    W_ir[6][10] = 11'b00000001000;
    W_ir[6][11] = 11'b00000000000;
    W_ir[6][12] = 11'b00000000000;
    W_ir[6][13] = 11'b00000000010;
    W_ir[6][14] = 11'b11111111110;
    W_ir[6][15] = 11'b11111111001;
    W_ir[6][16] = 11'b11111111101;
    W_ir[6][17] = 11'b00000000101;
    W_ir[6][18] = 11'b00000000000;
    W_ir[6][19] = 11'b00000000000;
    W_ir[6][20] = 11'b11111111111;
    W_ir[6][21] = 11'b11111111011;
    W_ir[6][22] = 11'b00000001001;
    W_ir[6][23] = 11'b00000000000;
    W_ir[6][24] = 11'b11111111011;
    W_ir[6][25] = 11'b00000000011;
    W_ir[6][26] = 11'b11111111010;
    W_ir[6][27] = 11'b11111111100;
    W_ir[6][28] = 11'b00000000110;
    W_ir[6][29] = 11'b00000000101;
    W_ir[6][30] = 11'b11111111011;
    W_ir[6][31] = 11'b00000000101;
    W_ir[6][32] = 11'b00000000000;
    W_ir[6][33] = 11'b00000000011;
    W_ir[6][34] = 11'b00000000111;
    W_ir[6][35] = 11'b00000001000;
    W_ir[6][36] = 11'b11111111111;
    W_ir[6][37] = 11'b00000000010;
    W_ir[6][38] = 11'b11111111000;
    W_ir[6][39] = 11'b11111111111;
    W_ir[6][40] = 11'b00000000100;
    W_ir[6][41] = 11'b11111111101;
    W_ir[6][42] = 11'b00000001001;
    W_ir[6][43] = 11'b00000000010;
    W_ir[6][44] = 11'b00000000100;
    W_ir[6][45] = 11'b11111111100;
    W_ir[6][46] = 11'b11111111001;
    W_ir[6][47] = 11'b00000001000;
    W_ir[6][48] = 11'b11111111010;
    W_ir[6][49] = 11'b11111111100;
    W_ir[6][50] = 11'b00000000100;
    W_ir[6][51] = 11'b11111111111;
    W_ir[6][52] = 11'b00000000100;
    W_ir[6][53] = 11'b11111110010;
    W_ir[6][54] = 11'b11111111110;
    W_ir[6][55] = 11'b00000000001;
    W_ir[6][56] = 11'b11111111011;
    W_ir[6][57] = 11'b11111111110;
    W_ir[6][58] = 11'b11111111011;
    W_ir[6][59] = 11'b11111111010;
    W_ir[6][60] = 11'b11111111110;
    W_ir[6][61] = 11'b11111110100;
    W_ir[6][62] = 11'b11111110001;
    W_ir[6][63] = 11'b11111110000;
    W_ir[7][0] = 11'b11111110101;
    W_ir[7][1] = 11'b11111110101;
    W_ir[7][2] = 11'b00000000011;
    W_ir[7][3] = 11'b11111111110;
    W_ir[7][4] = 11'b00000000110;
    W_ir[7][5] = 11'b00000001000;
    W_ir[7][6] = 11'b11111111001;
    W_ir[7][7] = 11'b00000000010;
    W_ir[7][8] = 11'b11111111011;
    W_ir[7][9] = 11'b11111110100;
    W_ir[7][10] = 11'b11111111100;
    W_ir[7][11] = 11'b00000000101;
    W_ir[7][12] = 11'b00000000110;
    W_ir[7][13] = 11'b11111111010;
    W_ir[7][14] = 11'b00000000110;
    W_ir[7][15] = 11'b00000000000;
    W_ir[7][16] = 11'b00000000001;
    W_ir[7][17] = 11'b11111111101;
    W_ir[7][18] = 11'b00000000001;
    W_ir[7][19] = 11'b00000000111;
    W_ir[7][20] = 11'b11111111100;
    W_ir[7][21] = 11'b11111111101;
    W_ir[7][22] = 11'b00000001000;
    W_ir[7][23] = 11'b11111111101;
    W_ir[7][24] = 11'b00000000111;
    W_ir[7][25] = 11'b00000000011;
    W_ir[7][26] = 11'b00000000100;
    W_ir[7][27] = 11'b11111111110;
    W_ir[7][28] = 11'b00000000110;
    W_ir[7][29] = 11'b00000001001;
    W_ir[7][30] = 11'b00000000110;
    W_ir[7][31] = 11'b00000000011;
    W_ir[7][32] = 11'b11111111011;
    W_ir[7][33] = 11'b11111111101;
    W_ir[7][34] = 11'b11111110100;
    W_ir[7][35] = 11'b11111111010;
    W_ir[7][36] = 11'b00000001000;
    W_ir[7][37] = 11'b00000000000;
    W_ir[7][38] = 11'b00000000110;
    W_ir[7][39] = 11'b11111110111;
    W_ir[7][40] = 11'b00000000000;
    W_ir[7][41] = 11'b11111111000;
    W_ir[7][42] = 11'b11111110111;
    W_ir[7][43] = 11'b11111110111;
    W_ir[7][44] = 11'b11111111011;
    W_ir[7][45] = 11'b00000000001;
    W_ir[7][46] = 11'b00000010010;
    W_ir[7][47] = 11'b11111111011;
    W_ir[7][48] = 11'b11111111111;
    W_ir[7][49] = 11'b11111111011;
    W_ir[7][50] = 11'b11111111000;
    W_ir[7][51] = 11'b00000001100;
    W_ir[7][52] = 11'b11111110111;
    W_ir[7][53] = 11'b00000000011;
    W_ir[7][54] = 11'b00000001001;
    W_ir[7][55] = 11'b00000000001;
    W_ir[7][56] = 11'b00000010010;
    W_ir[7][57] = 11'b00000000010;
    W_ir[7][58] = 11'b00000010011;
    W_ir[7][59] = 11'b00000000011;
    W_ir[7][60] = 11'b11111111000;
    W_ir[7][61] = 11'b00000001001;
    W_ir[7][62] = 11'b00000001100;
    W_ir[7][63] = 11'b11111111000;
    W_ir[8][0] = 11'b11111111100;
    W_ir[8][1] = 11'b00000000010;
    W_ir[8][2] = 11'b11111111110;
    W_ir[8][3] = 11'b00000000100;
    W_ir[8][4] = 11'b11111111111;
    W_ir[8][5] = 11'b11111111110;
    W_ir[8][6] = 11'b11111111001;
    W_ir[8][7] = 11'b11111111100;
    W_ir[8][8] = 11'b11111111110;
    W_ir[8][9] = 11'b00000000101;
    W_ir[8][10] = 11'b00000000010;
    W_ir[8][11] = 11'b00000000111;
    W_ir[8][12] = 11'b11111111110;
    W_ir[8][13] = 11'b00000000100;
    W_ir[8][14] = 11'b00000000100;
    W_ir[8][15] = 11'b00000000010;
    W_ir[8][16] = 11'b11111111111;
    W_ir[8][17] = 11'b00000000101;
    W_ir[8][18] = 11'b00000001000;
    W_ir[8][19] = 11'b00000000100;
    W_ir[8][20] = 11'b11111111111;
    W_ir[8][21] = 11'b00000000001;
    W_ir[8][22] = 11'b00000000110;
    W_ir[8][23] = 11'b00000000001;
    W_ir[8][24] = 11'b00000000000;
    W_ir[8][25] = 11'b11111111111;
    W_ir[8][26] = 11'b11111111001;
    W_ir[8][27] = 11'b00000000010;
    W_ir[8][28] = 11'b00000000100;
    W_ir[8][29] = 11'b00000000000;
    W_ir[8][30] = 11'b00000000101;
    W_ir[8][31] = 11'b00000000100;
    W_ir[8][32] = 11'b11111111111;
    W_ir[8][33] = 11'b11111111011;
    W_ir[8][34] = 11'b11111111010;
    W_ir[8][35] = 11'b11111111101;
    W_ir[8][36] = 11'b11111111101;
    W_ir[8][37] = 11'b11111110110;
    W_ir[8][38] = 11'b00000000010;
    W_ir[8][39] = 11'b11111111111;
    W_ir[8][40] = 11'b11111111111;
    W_ir[8][41] = 11'b00000000111;
    W_ir[8][42] = 11'b11111111011;
    W_ir[8][43] = 11'b00000000100;
    W_ir[8][44] = 11'b00000000000;
    W_ir[8][45] = 11'b11111111100;
    W_ir[8][46] = 11'b11111111011;
    W_ir[8][47] = 11'b00000000101;
    W_ir[8][48] = 11'b00000000010;
    W_ir[8][49] = 11'b00000001001;
    W_ir[8][50] = 11'b00000000000;
    W_ir[8][51] = 11'b00000000010;
    W_ir[8][52] = 11'b11111111110;
    W_ir[8][53] = 11'b11111111010;
    W_ir[8][54] = 11'b11111111001;
    W_ir[8][55] = 11'b11111111101;
    W_ir[8][56] = 11'b00000000111;
    W_ir[8][57] = 11'b11111111110;
    W_ir[8][58] = 11'b00000001000;
    W_ir[8][59] = 11'b11111111110;
    W_ir[8][60] = 11'b11111110111;
    W_ir[8][61] = 11'b11111110010;
    W_ir[8][62] = 11'b11111110000;
    W_ir[8][63] = 11'b00000000011;
    W_ir[9][0] = 11'b00000000110;
    W_ir[9][1] = 11'b00000000010;
    W_ir[9][2] = 11'b00000000001;
    W_ir[9][3] = 11'b00000000000;
    W_ir[9][4] = 11'b00000000001;
    W_ir[9][5] = 11'b00000000101;
    W_ir[9][6] = 11'b11111111010;
    W_ir[9][7] = 11'b11111111011;
    W_ir[9][8] = 11'b00000000000;
    W_ir[9][9] = 11'b00000001000;
    W_ir[9][10] = 11'b00000000100;
    W_ir[9][11] = 11'b11111111000;
    W_ir[9][12] = 11'b11111111011;
    W_ir[9][13] = 11'b00000000101;
    W_ir[9][14] = 11'b11111111110;
    W_ir[9][15] = 11'b00000000110;
    W_ir[9][16] = 11'b11111111000;
    W_ir[9][17] = 11'b00000000100;
    W_ir[9][18] = 11'b00000001001;
    W_ir[9][19] = 11'b11111111011;
    W_ir[9][20] = 11'b11111111011;
    W_ir[9][21] = 11'b11111111001;
    W_ir[9][22] = 11'b00000000100;
    W_ir[9][23] = 11'b00000001010;
    W_ir[9][24] = 11'b00000000100;
    W_ir[9][25] = 11'b11111111100;
    W_ir[9][26] = 11'b11111111101;
    W_ir[9][27] = 11'b11111111100;
    W_ir[9][28] = 11'b11111111101;
    W_ir[9][29] = 11'b11111111010;
    W_ir[9][30] = 11'b11111111110;
    W_ir[9][31] = 11'b11111111010;
    W_ir[9][32] = 11'b00000000101;
    W_ir[9][33] = 11'b11111111110;
    W_ir[9][34] = 11'b11111111100;
    W_ir[9][35] = 11'b00000000101;
    W_ir[9][36] = 11'b11111110111;
    W_ir[9][37] = 11'b00000000001;
    W_ir[9][38] = 11'b00000000000;
    W_ir[9][39] = 11'b11111111100;
    W_ir[9][40] = 11'b00000000110;
    W_ir[9][41] = 11'b00000000011;
    W_ir[9][42] = 11'b00000000111;
    W_ir[9][43] = 11'b00000000110;
    W_ir[9][44] = 11'b00000000000;
    W_ir[9][45] = 11'b00000000111;
    W_ir[9][46] = 11'b00000000010;
    W_ir[9][47] = 11'b11111111110;
    W_ir[9][48] = 11'b11111111010;
    W_ir[9][49] = 11'b11111111111;
    W_ir[9][50] = 11'b11111111101;
    W_ir[9][51] = 11'b00000000100;
    W_ir[9][52] = 11'b00000000101;
    W_ir[9][53] = 11'b00000000011;
    W_ir[9][54] = 11'b11111111000;
    W_ir[9][55] = 11'b00000001010;
    W_ir[9][56] = 11'b00000000101;
    W_ir[9][57] = 11'b11111111110;
    W_ir[9][58] = 11'b11111111111;
    W_ir[9][59] = 11'b00000000111;
    W_ir[9][60] = 11'b11111110111;
    W_ir[9][61] = 11'b00000000000;
    W_ir[9][62] = 11'b11111111101;
    W_ir[9][63] = 11'b11111111101;
    W_ir[10][0] = 11'b00000000011;
    W_ir[10][1] = 11'b00000000100;
    W_ir[10][2] = 11'b11111111111;
    W_ir[10][3] = 11'b00000000010;
    W_ir[10][4] = 11'b00000000110;
    W_ir[10][5] = 11'b00000000011;
    W_ir[10][6] = 11'b11111110111;
    W_ir[10][7] = 11'b00000000011;
    W_ir[10][8] = 11'b11111110100;
    W_ir[10][9] = 11'b11111111110;
    W_ir[10][10] = 11'b00000000000;
    W_ir[10][11] = 11'b11111111100;
    W_ir[10][12] = 11'b11111111001;
    W_ir[10][13] = 11'b00000000011;
    W_ir[10][14] = 11'b00000000000;
    W_ir[10][15] = 11'b11111110101;
    W_ir[10][16] = 11'b00000000100;
    W_ir[10][17] = 11'b00000000101;
    W_ir[10][18] = 11'b11111110100;
    W_ir[10][19] = 11'b11111111000;
    W_ir[10][20] = 11'b00000000111;
    W_ir[10][21] = 11'b11111111010;
    W_ir[10][22] = 11'b00000000011;
    W_ir[10][23] = 11'b11111111010;
    W_ir[10][24] = 11'b00000000011;
    W_ir[10][25] = 11'b11111111011;
    W_ir[10][26] = 11'b00000001001;
    W_ir[10][27] = 11'b11111111110;
    W_ir[10][28] = 11'b00000000110;
    W_ir[10][29] = 11'b00000001001;
    W_ir[10][30] = 11'b11111111111;
    W_ir[10][31] = 11'b00000000000;
    W_ir[10][32] = 11'b00000001011;
    W_ir[10][33] = 11'b11111111000;
    W_ir[10][34] = 11'b11111111000;
    W_ir[10][35] = 11'b11111111100;
    W_ir[10][36] = 11'b00000001010;
    W_ir[10][37] = 11'b00000001000;
    W_ir[10][38] = 11'b11111111011;
    W_ir[10][39] = 11'b11111110101;
    W_ir[10][40] = 11'b00000000100;
    W_ir[10][41] = 11'b11111111111;
    W_ir[10][42] = 11'b11111111000;
    W_ir[10][43] = 11'b00000000001;
    W_ir[10][44] = 11'b11111111101;
    W_ir[10][45] = 11'b00000000101;
    W_ir[10][46] = 11'b11111111110;
    W_ir[10][47] = 11'b11111111110;
    W_ir[10][48] = 11'b11111111101;
    W_ir[10][49] = 11'b00000000000;
    W_ir[10][50] = 11'b11111111000;
    W_ir[10][51] = 11'b11111111101;
    W_ir[10][52] = 11'b11111111000;
    W_ir[10][53] = 11'b00000000111;
    W_ir[10][54] = 11'b11111111111;
    W_ir[10][55] = 11'b11111111100;
    W_ir[10][56] = 11'b11111111101;
    W_ir[10][57] = 11'b00000000111;
    W_ir[10][58] = 11'b00000001000;
    W_ir[10][59] = 11'b00000001010;
    W_ir[10][60] = 11'b00000001111;
    W_ir[10][61] = 11'b00000001010;
    W_ir[10][62] = 11'b00000010001;
    W_ir[10][63] = 11'b00000001101;
    W_ir[11][0] = 11'b11111110101;
    W_ir[11][1] = 11'b00000001000;
    W_ir[11][2] = 11'b00000000001;
    W_ir[11][3] = 11'b00000001001;
    W_ir[11][4] = 11'b11111110110;
    W_ir[11][5] = 11'b00000000010;
    W_ir[11][6] = 11'b11111110111;
    W_ir[11][7] = 11'b00000000101;
    W_ir[11][8] = 11'b11111110010;
    W_ir[11][9] = 11'b11111110101;
    W_ir[11][10] = 11'b00000001001;
    W_ir[11][11] = 11'b11111110101;
    W_ir[11][12] = 11'b11111110101;
    W_ir[11][13] = 11'b00000000101;
    W_ir[11][14] = 11'b00000000100;
    W_ir[11][15] = 11'b00000000100;
    W_ir[11][16] = 11'b00000001011;
    W_ir[11][17] = 11'b11111111110;
    W_ir[11][18] = 11'b00000000000;
    W_ir[11][19] = 11'b00000001101;
    W_ir[11][20] = 11'b11111111110;
    W_ir[11][21] = 11'b11111111000;
    W_ir[11][22] = 11'b11111111101;
    W_ir[11][23] = 11'b11111111100;
    W_ir[11][24] = 11'b11111110110;
    W_ir[11][25] = 11'b11111111110;
    W_ir[11][26] = 11'b11111111000;
    W_ir[11][27] = 11'b11111110110;
    W_ir[11][28] = 11'b00000001101;
    W_ir[11][29] = 11'b00000000100;
    W_ir[11][30] = 11'b00000000001;
    W_ir[11][31] = 11'b00000000111;
    W_ir[11][32] = 11'b00000000100;
    W_ir[11][33] = 11'b11111111110;
    W_ir[11][34] = 11'b00000000111;
    W_ir[11][35] = 11'b00000000100;
    W_ir[11][36] = 11'b11111110111;
    W_ir[11][37] = 11'b11111110110;
    W_ir[11][38] = 11'b00000000100;
    W_ir[11][39] = 11'b00000000000;
    W_ir[11][40] = 11'b11111110100;
    W_ir[11][41] = 11'b11111110110;
    W_ir[11][42] = 11'b00000001000;
    W_ir[11][43] = 11'b00000000001;
    W_ir[11][44] = 11'b00000000011;
    W_ir[11][45] = 11'b00000001100;
    W_ir[11][46] = 11'b11111111111;
    W_ir[11][47] = 11'b00000001010;
    W_ir[11][48] = 11'b00000000001;
    W_ir[11][49] = 11'b11111111111;
    W_ir[11][50] = 11'b11111111011;
    W_ir[11][51] = 11'b00000000110;
    W_ir[11][52] = 11'b11111111110;
    W_ir[11][53] = 11'b11111110110;
    W_ir[11][54] = 11'b00000001100;
    W_ir[11][55] = 11'b00000000010;
    W_ir[11][56] = 11'b11111111010;
    W_ir[11][57] = 11'b00000000110;
    W_ir[11][58] = 11'b11111111011;
    W_ir[11][59] = 11'b00000001011;
    W_ir[11][60] = 11'b00000001011;
    W_ir[11][61] = 11'b00000000011;
    W_ir[11][62] = 11'b00000000001;
    W_ir[11][63] = 11'b00000001001;
    W_ir[12][0] = 11'b00000000011;
    W_ir[12][1] = 11'b00000000101;
    W_ir[12][2] = 11'b00000000100;
    W_ir[12][3] = 11'b00000000100;
    W_ir[12][4] = 11'b11111111110;
    W_ir[12][5] = 11'b11111111011;
    W_ir[12][6] = 11'b00000000100;
    W_ir[12][7] = 11'b00000000010;
    W_ir[12][8] = 11'b11111111001;
    W_ir[12][9] = 11'b00000000001;
    W_ir[12][10] = 11'b00000001000;
    W_ir[12][11] = 11'b00000000000;
    W_ir[12][12] = 11'b00000000101;
    W_ir[12][13] = 11'b00000000001;
    W_ir[12][14] = 11'b00000000001;
    W_ir[12][15] = 11'b00000000110;
    W_ir[12][16] = 11'b11111111111;
    W_ir[12][17] = 11'b00000000111;
    W_ir[12][18] = 11'b11111111111;
    W_ir[12][19] = 11'b00000000101;
    W_ir[12][20] = 11'b11111111111;
    W_ir[12][21] = 11'b00000000100;
    W_ir[12][22] = 11'b00000000011;
    W_ir[12][23] = 11'b00000000011;
    W_ir[12][24] = 11'b11111111011;
    W_ir[12][25] = 11'b00000000100;
    W_ir[12][26] = 11'b00000000100;
    W_ir[12][27] = 11'b00000000011;
    W_ir[12][28] = 11'b00000000111;
    W_ir[12][29] = 11'b11111111001;
    W_ir[12][30] = 11'b11111111110;
    W_ir[12][31] = 11'b00000000011;
    W_ir[12][32] = 11'b00000000010;
    W_ir[12][33] = 11'b00000000100;
    W_ir[12][34] = 11'b00000000100;
    W_ir[12][35] = 11'b00000000001;
    W_ir[12][36] = 11'b00000001000;
    W_ir[12][37] = 11'b00000000011;
    W_ir[12][38] = 11'b11111111110;
    W_ir[12][39] = 11'b00000000010;
    W_ir[12][40] = 11'b00000000101;
    W_ir[12][41] = 11'b11111111010;
    W_ir[12][42] = 11'b00000000010;
    W_ir[12][43] = 11'b11111111101;
    W_ir[12][44] = 11'b00000000000;
    W_ir[12][45] = 11'b11111111100;
    W_ir[12][46] = 11'b11111111010;
    W_ir[12][47] = 11'b00000000111;
    W_ir[12][48] = 11'b11111111110;
    W_ir[12][49] = 11'b11111111101;
    W_ir[12][50] = 11'b11111111111;
    W_ir[12][51] = 11'b00000000000;
    W_ir[12][52] = 11'b11111111001;
    W_ir[12][53] = 11'b11111111101;
    W_ir[12][54] = 11'b00000000010;
    W_ir[12][55] = 11'b11111111101;
    W_ir[12][56] = 11'b00000000101;
    W_ir[12][57] = 11'b11111111101;
    W_ir[12][58] = 11'b11111111101;
    W_ir[12][59] = 11'b00000000100;
    W_ir[12][60] = 11'b11111111011;
    W_ir[12][61] = 11'b11111111010;
    W_ir[12][62] = 11'b11111111010;
    W_ir[12][63] = 11'b00000000100;
    W_ir[13][0] = 11'b11111111100;
    W_ir[13][1] = 11'b11111111101;
    W_ir[13][2] = 11'b00000000110;
    W_ir[13][3] = 11'b00000000101;
    W_ir[13][4] = 11'b00000000001;
    W_ir[13][5] = 11'b00000000010;
    W_ir[13][6] = 11'b00000000010;
    W_ir[13][7] = 11'b00000000001;
    W_ir[13][8] = 11'b00000000001;
    W_ir[13][9] = 11'b00000000001;
    W_ir[13][10] = 11'b11111111111;
    W_ir[13][11] = 11'b00000000000;
    W_ir[13][12] = 11'b00000000001;
    W_ir[13][13] = 11'b00000000100;
    W_ir[13][14] = 11'b11111111011;
    W_ir[13][15] = 11'b00000000001;
    W_ir[13][16] = 11'b00000000000;
    W_ir[13][17] = 11'b00000000000;
    W_ir[13][18] = 11'b00000000000;
    W_ir[13][19] = 11'b11111111101;
    W_ir[13][20] = 11'b00000000000;
    W_ir[13][21] = 11'b00000000001;
    W_ir[13][22] = 11'b11111111110;
    W_ir[13][23] = 11'b11111111101;
    W_ir[13][24] = 11'b00000000000;
    W_ir[13][25] = 11'b00000000110;
    W_ir[13][26] = 11'b11111111010;
    W_ir[13][27] = 11'b11111111010;
    W_ir[13][28] = 11'b00000000111;
    W_ir[13][29] = 11'b00000000010;
    W_ir[13][30] = 11'b00000000000;
    W_ir[13][31] = 11'b00000000000;
    W_ir[13][32] = 11'b11111111100;
    W_ir[13][33] = 11'b00000000000;
    W_ir[13][34] = 11'b11111111111;
    W_ir[13][35] = 11'b00000000000;
    W_ir[13][36] = 11'b00000000010;
    W_ir[13][37] = 11'b00000000001;
    W_ir[13][38] = 11'b00000000010;
    W_ir[13][39] = 11'b00000000100;
    W_ir[13][40] = 11'b00000000010;
    W_ir[13][41] = 11'b00000000000;
    W_ir[13][42] = 11'b00000000000;
    W_ir[13][43] = 11'b00000000010;
    W_ir[13][44] = 11'b00000000001;
    W_ir[13][45] = 11'b00000000010;
    W_ir[13][46] = 11'b00000000000;
    W_ir[13][47] = 11'b11111111111;
    W_ir[13][48] = 11'b11111111111;
    W_ir[13][49] = 11'b11111111001;
    W_ir[13][50] = 11'b00000000100;
    W_ir[13][51] = 11'b00000000101;
    W_ir[13][52] = 11'b11111111110;
    W_ir[13][53] = 11'b11111111101;
    W_ir[13][54] = 11'b11111111101;
    W_ir[13][55] = 11'b11111111101;
    W_ir[13][56] = 11'b11111111110;
    W_ir[13][57] = 11'b00000000110;
    W_ir[13][58] = 11'b00000000100;
    W_ir[13][59] = 11'b11111111100;
    W_ir[13][60] = 11'b11111111111;
    W_ir[13][61] = 11'b11111111110;
    W_ir[13][62] = 11'b00000000101;
    W_ir[13][63] = 11'b11111111101;
    W_ir[14][0] = 11'b11111111101;
    W_ir[14][1] = 11'b11111111110;
    W_ir[14][2] = 11'b11111111001;
    W_ir[14][3] = 11'b11111111100;
    W_ir[14][4] = 11'b11111111110;
    W_ir[14][5] = 11'b11111111111;
    W_ir[14][6] = 11'b00000000001;
    W_ir[14][7] = 11'b11111111011;
    W_ir[14][8] = 11'b11111111111;
    W_ir[14][9] = 11'b11111111111;
    W_ir[14][10] = 11'b11111111111;
    W_ir[14][11] = 11'b11111111001;
    W_ir[14][12] = 11'b11111111111;
    W_ir[14][13] = 11'b00000000010;
    W_ir[14][14] = 11'b11111111111;
    W_ir[14][15] = 11'b00000000011;
    W_ir[14][16] = 11'b11111111011;
    W_ir[14][17] = 11'b00000000111;
    W_ir[14][18] = 11'b00000000000;
    W_ir[14][19] = 11'b00000000010;
    W_ir[14][20] = 11'b00000000010;
    W_ir[14][21] = 11'b11111111110;
    W_ir[14][22] = 11'b00000000100;
    W_ir[14][23] = 11'b00000000111;
    W_ir[14][24] = 11'b00000000011;
    W_ir[14][25] = 11'b00000000001;
    W_ir[14][26] = 11'b00000000000;
    W_ir[14][27] = 11'b11111111001;
    W_ir[14][28] = 11'b11111111110;
    W_ir[14][29] = 11'b00000001000;
    W_ir[14][30] = 11'b11111111101;
    W_ir[14][31] = 11'b11111111101;
    W_ir[14][32] = 11'b00000000000;
    W_ir[14][33] = 11'b00000000011;
    W_ir[14][34] = 11'b11111111111;
    W_ir[14][35] = 11'b11111111110;
    W_ir[14][36] = 11'b00000000000;
    W_ir[14][37] = 11'b00000000001;
    W_ir[14][38] = 11'b00000000100;
    W_ir[14][39] = 11'b00000000000;
    W_ir[14][40] = 11'b00000000100;
    W_ir[14][41] = 11'b11111111110;
    W_ir[14][42] = 11'b00000000100;
    W_ir[14][43] = 11'b00000000000;
    W_ir[14][44] = 11'b00000000001;
    W_ir[14][45] = 11'b00000000010;
    W_ir[14][46] = 11'b00000000010;
    W_ir[14][47] = 11'b00000000001;
    W_ir[14][48] = 11'b00000000010;
    W_ir[14][49] = 11'b00000000001;
    W_ir[14][50] = 11'b11111111100;
    W_ir[14][51] = 11'b00000000011;
    W_ir[14][52] = 11'b00000000011;
    W_ir[14][53] = 11'b00000000010;
    W_ir[14][54] = 11'b11111111001;
    W_ir[14][55] = 11'b00000000010;
    W_ir[14][56] = 11'b00000000010;
    W_ir[14][57] = 11'b11111111011;
    W_ir[14][58] = 11'b11111111100;
    W_ir[14][59] = 11'b11111111101;
    W_ir[14][60] = 11'b00000000101;
    W_ir[14][61] = 11'b00000000010;
    W_ir[14][62] = 11'b00000000101;
    W_ir[14][63] = 11'b00000001001;
    W_ir[15][0] = 11'b00000000000;
    W_ir[15][1] = 11'b00000001000;
    W_ir[15][2] = 11'b00000000000;
    W_ir[15][3] = 11'b00000000110;
    W_ir[15][4] = 11'b11111111010;
    W_ir[15][5] = 11'b00000000001;
    W_ir[15][6] = 11'b00000000001;
    W_ir[15][7] = 11'b11111111110;
    W_ir[15][8] = 11'b11111111111;
    W_ir[15][9] = 11'b00000000101;
    W_ir[15][10] = 11'b11111111100;
    W_ir[15][11] = 11'b11111111111;
    W_ir[15][12] = 11'b11111111100;
    W_ir[15][13] = 11'b11111111111;
    W_ir[15][14] = 11'b11111111110;
    W_ir[15][15] = 11'b11111111111;
    W_ir[15][16] = 11'b00000000000;
    W_ir[15][17] = 11'b00000000001;
    W_ir[15][18] = 11'b11111111101;
    W_ir[15][19] = 11'b00000000100;
    W_ir[15][20] = 11'b11111111110;
    W_ir[15][21] = 11'b00000000010;
    W_ir[15][22] = 11'b00000000011;
    W_ir[15][23] = 11'b00000000010;
    W_ir[15][24] = 11'b00000000111;
    W_ir[15][25] = 11'b00000000001;
    W_ir[15][26] = 11'b11111111111;
    W_ir[15][27] = 11'b11111111110;
    W_ir[15][28] = 11'b00000000001;
    W_ir[15][29] = 11'b00000000001;
    W_ir[15][30] = 11'b11111111100;
    W_ir[15][31] = 11'b00000001000;
    W_ir[15][32] = 11'b00000000100;
    W_ir[15][33] = 11'b11111111011;
    W_ir[15][34] = 11'b00000000010;
    W_ir[15][35] = 11'b00000000001;
    W_ir[15][36] = 11'b00000000001;
    W_ir[15][37] = 11'b11111111001;
    W_ir[15][38] = 11'b00000000011;
    W_ir[15][39] = 11'b00000000000;
    W_ir[15][40] = 11'b00000000000;
    W_ir[15][41] = 11'b00000000101;
    W_ir[15][42] = 11'b11111111011;
    W_ir[15][43] = 11'b00000000001;
    W_ir[15][44] = 11'b11111111101;
    W_ir[15][45] = 11'b11111111110;
    W_ir[15][46] = 11'b00000000110;
    W_ir[15][47] = 11'b11111111101;
    W_ir[15][48] = 11'b11111111110;
    W_ir[15][49] = 11'b11111111111;
    W_ir[15][50] = 11'b11111111100;
    W_ir[15][51] = 11'b11111111101;
    W_ir[15][52] = 11'b11111111101;
    W_ir[15][53] = 11'b11111111100;
    W_ir[15][54] = 11'b11111111110;
    W_ir[15][55] = 11'b11111111001;
    W_ir[15][56] = 11'b11111111101;
    W_ir[15][57] = 11'b00000000100;
    W_ir[15][58] = 11'b11111111100;
    W_ir[15][59] = 11'b11111111101;
    W_ir[15][60] = 11'b11111111101;
    W_ir[15][61] = 11'b11111111101;
    W_ir[15][62] = 11'b11111111010;
    W_ir[15][63] = 11'b11111111110;

    // Initialize W_iz weights
    W_iz[0][0] = 11'b00000000000;
    W_iz[0][1] = 11'b11111111110;
    W_iz[0][2] = 11'b11111111111;
    W_iz[0][3] = 11'b11111111101;
    W_iz[0][4] = 11'b00000000000;
    W_iz[0][5] = 11'b00000000011;
    W_iz[0][6] = 11'b11111111100;
    W_iz[0][7] = 11'b11111111011;
    W_iz[0][8] = 11'b11111111001;
    W_iz[0][9] = 11'b11111111101;
    W_iz[0][10] = 11'b11111111001;
    W_iz[0][11] = 11'b11111111110;
    W_iz[0][12] = 11'b11111111111;
    W_iz[0][13] = 11'b00000000011;
    W_iz[0][14] = 11'b00000000001;
    W_iz[0][15] = 11'b11111111111;
    W_iz[0][16] = 11'b11111111100;
    W_iz[0][17] = 11'b11111111101;
    W_iz[0][18] = 11'b11111111100;
    W_iz[0][19] = 11'b11111111011;
    W_iz[0][20] = 11'b11111111111;
    W_iz[0][21] = 11'b00000000011;
    W_iz[0][22] = 11'b00000001000;
    W_iz[0][23] = 11'b00000000101;
    W_iz[0][24] = 11'b11111111001;
    W_iz[0][25] = 11'b11111111010;
    W_iz[0][26] = 11'b00000000000;
    W_iz[0][27] = 11'b11111111001;
    W_iz[0][28] = 11'b00000000110;
    W_iz[0][29] = 11'b00000000000;
    W_iz[0][30] = 11'b00000000110;
    W_iz[0][31] = 11'b11111111100;
    W_iz[0][32] = 11'b11111111001;
    W_iz[0][33] = 11'b11111111010;
    W_iz[0][34] = 11'b11111111100;
    W_iz[0][35] = 11'b11111111100;
    W_iz[0][36] = 11'b11111111010;
    W_iz[0][37] = 11'b11111111011;
    W_iz[0][38] = 11'b11111111101;
    W_iz[0][39] = 11'b00000000010;
    W_iz[0][40] = 11'b00000000001;
    W_iz[0][41] = 11'b11111111100;
    W_iz[0][42] = 11'b11111111111;
    W_iz[0][43] = 11'b11111111101;
    W_iz[0][44] = 11'b11111111000;
    W_iz[0][45] = 11'b11111111111;
    W_iz[0][46] = 11'b11111111111;
    W_iz[0][47] = 11'b11111111111;
    W_iz[0][48] = 11'b00000000000;
    W_iz[0][49] = 11'b11111111110;
    W_iz[0][50] = 11'b00000000101;
    W_iz[0][51] = 11'b11111111101;
    W_iz[0][52] = 11'b00000000111;
    W_iz[0][53] = 11'b00000000100;
    W_iz[0][54] = 11'b00000001000;
    W_iz[0][55] = 11'b00000000110;
    W_iz[0][56] = 11'b00000000011;
    W_iz[0][57] = 11'b11111111001;
    W_iz[0][58] = 11'b00000000100;
    W_iz[0][59] = 11'b00000001110;
    W_iz[0][60] = 11'b00000001010;
    W_iz[0][61] = 11'b00000001011;
    W_iz[0][62] = 11'b00000001101;
    W_iz[0][63] = 11'b00000001100;
    W_iz[1][0] = 11'b00000000001;
    W_iz[1][1] = 11'b00000000001;
    W_iz[1][2] = 11'b00000000010;
    W_iz[1][3] = 11'b11111111111;
    W_iz[1][4] = 11'b11111111111;
    W_iz[1][5] = 11'b11111111011;
    W_iz[1][6] = 11'b00000000110;
    W_iz[1][7] = 11'b11111111001;
    W_iz[1][8] = 11'b11111111010;
    W_iz[1][9] = 11'b11111111110;
    W_iz[1][10] = 11'b00000000000;
    W_iz[1][11] = 11'b11111111111;
    W_iz[1][12] = 11'b11111111100;
    W_iz[1][13] = 11'b11111111111;
    W_iz[1][14] = 11'b11111111100;
    W_iz[1][15] = 11'b11111111100;
    W_iz[1][16] = 11'b00000000101;
    W_iz[1][17] = 11'b11111111011;
    W_iz[1][18] = 11'b00000000001;
    W_iz[1][19] = 11'b11111111010;
    W_iz[1][20] = 11'b11111111111;
    W_iz[1][21] = 11'b00000000000;
    W_iz[1][22] = 11'b00000000011;
    W_iz[1][23] = 11'b00000000010;
    W_iz[1][24] = 11'b11111111111;
    W_iz[1][25] = 11'b11111111101;
    W_iz[1][26] = 11'b11111111111;
    W_iz[1][27] = 11'b00000000011;
    W_iz[1][28] = 11'b00000000001;
    W_iz[1][29] = 11'b11111111100;
    W_iz[1][30] = 11'b11111111110;
    W_iz[1][31] = 11'b11111111001;
    W_iz[1][32] = 11'b00000000000;
    W_iz[1][33] = 11'b11111111000;
    W_iz[1][34] = 11'b11111111110;
    W_iz[1][35] = 11'b00000000100;
    W_iz[1][36] = 11'b11111111100;
    W_iz[1][37] = 11'b11111111010;
    W_iz[1][38] = 11'b11111110111;
    W_iz[1][39] = 11'b00000000101;
    W_iz[1][40] = 11'b11111111101;
    W_iz[1][41] = 11'b11111111111;
    W_iz[1][42] = 11'b00000000000;
    W_iz[1][43] = 11'b11111111101;
    W_iz[1][44] = 11'b00000000001;
    W_iz[1][45] = 11'b11111111101;
    W_iz[1][46] = 11'b11111111111;
    W_iz[1][47] = 11'b00000000100;
    W_iz[1][48] = 11'b00000000010;
    W_iz[1][49] = 11'b00000000010;
    W_iz[1][50] = 11'b00000000001;
    W_iz[1][51] = 11'b00000000001;
    W_iz[1][52] = 11'b11111111110;
    W_iz[1][53] = 11'b11111111101;
    W_iz[1][54] = 11'b00000000010;
    W_iz[1][55] = 11'b00000000000;
    W_iz[1][56] = 11'b00000000001;
    W_iz[1][57] = 11'b11111111011;
    W_iz[1][58] = 11'b11111111100;
    W_iz[1][59] = 11'b11111111110;
    W_iz[1][60] = 11'b00000000111;
    W_iz[1][61] = 11'b00000000101;
    W_iz[1][62] = 11'b11111111110;
    W_iz[1][63] = 11'b00000000101;
    W_iz[2][0] = 11'b00000000110;
    W_iz[2][1] = 11'b11111111110;
    W_iz[2][2] = 11'b00000001001;
    W_iz[2][3] = 11'b11111111110;
    W_iz[2][4] = 11'b00000000101;
    W_iz[2][5] = 11'b00000000001;
    W_iz[2][6] = 11'b11111111001;
    W_iz[2][7] = 11'b00000001001;
    W_iz[2][8] = 11'b00000001011;
    W_iz[2][9] = 11'b00000000110;
    W_iz[2][10] = 11'b00000001000;
    W_iz[2][11] = 11'b00000000000;
    W_iz[2][12] = 11'b00000000000;
    W_iz[2][13] = 11'b00000000010;
    W_iz[2][14] = 11'b11111111110;
    W_iz[2][15] = 11'b11111111001;
    W_iz[2][16] = 11'b11111111101;
    W_iz[2][17] = 11'b00000000101;
    W_iz[2][18] = 11'b00000000000;
    W_iz[2][19] = 11'b00000000000;
    W_iz[2][20] = 11'b11111111111;
    W_iz[2][21] = 11'b11111111011;
    W_iz[2][22] = 11'b00000001001;
    W_iz[2][23] = 11'b00000000000;
    W_iz[2][24] = 11'b11111111011;
    W_iz[2][25] = 11'b00000000011;
    W_iz[2][26] = 11'b11111111010;
    W_iz[2][27] = 11'b11111111100;
    W_iz[2][28] = 11'b00000000110;
    W_iz[2][29] = 11'b00000000101;
    W_iz[2][30] = 11'b11111111011;
    W_iz[2][31] = 11'b00000000101;
    W_iz[2][32] = 11'b00000000000;
    W_iz[2][33] = 11'b00000000011;
    W_iz[2][34] = 11'b00000000111;
    W_iz[2][35] = 11'b00000001000;
    W_iz[2][36] = 11'b11111111111;
    W_iz[2][37] = 11'b00000000010;
    W_iz[2][38] = 11'b11111111000;
    W_iz[2][39] = 11'b11111111111;
    W_iz[2][40] = 11'b00000000100;
    W_iz[2][41] = 11'b11111111101;
    W_iz[2][42] = 11'b00000001001;
    W_iz[2][43] = 11'b00000000010;
    W_iz[2][44] = 11'b00000000100;
    W_iz[2][45] = 11'b11111111100;
    W_iz[2][46] = 11'b11111111001;
    W_iz[2][47] = 11'b00000001000;
    W_iz[2][48] = 11'b11111111010;
    W_iz[2][49] = 11'b11111111100;
    W_iz[2][50] = 11'b00000000100;
    W_iz[2][51] = 11'b11111111111;
    W_iz[2][52] = 11'b00000000100;
    W_iz[2][53] = 11'b11111110010;
    W_iz[2][54] = 11'b11111111110;
    W_iz[2][55] = 11'b00000000001;
    W_iz[2][56] = 11'b11111111011;
    W_iz[2][57] = 11'b11111111110;
    W_iz[2][58] = 11'b11111111011;
    W_iz[2][59] = 11'b11111111010;
    W_iz[2][60] = 11'b11111111110;
    W_iz[2][61] = 11'b11111110100;
    W_iz[2][62] = 11'b11111110001;
    W_iz[2][63] = 11'b11111110000;
    W_iz[3][0] = 11'b11111110101;
    W_iz[3][1] = 11'b11111110101;
    W_iz[3][2] = 11'b00000000011;
    W_iz[3][3] = 11'b11111111110;
    W_iz[3][4] = 11'b00000000110;
    W_iz[3][5] = 11'b00000001000;
    W_iz[3][6] = 11'b11111111001;
    W_iz[3][7] = 11'b00000000010;
    W_iz[3][8] = 11'b11111111011;
    W_iz[3][9] = 11'b11111110100;
    W_iz[3][10] = 11'b11111111100;
    W_iz[3][11] = 11'b00000000101;
    W_iz[3][12] = 11'b00000000110;
    W_iz[3][13] = 11'b11111111010;
    W_iz[3][14] = 11'b00000000110;
    W_iz[3][15] = 11'b00000000000;
    W_iz[3][16] = 11'b00000000001;
    W_iz[3][17] = 11'b11111111101;
    W_iz[3][18] = 11'b00000000001;
    W_iz[3][19] = 11'b00000000111;
    W_iz[3][20] = 11'b11111111100;
    W_iz[3][21] = 11'b11111111101;
    W_iz[3][22] = 11'b00000001000;
    W_iz[3][23] = 11'b11111111101;
    W_iz[3][24] = 11'b00000000111;
    W_iz[3][25] = 11'b00000000011;
    W_iz[3][26] = 11'b00000000100;
    W_iz[3][27] = 11'b11111111110;
    W_iz[3][28] = 11'b00000000110;
    W_iz[3][29] = 11'b00000001001;
    W_iz[3][30] = 11'b00000000110;
    W_iz[3][31] = 11'b00000000011;
    W_iz[3][32] = 11'b11111111011;
    W_iz[3][33] = 11'b11111111101;
    W_iz[3][34] = 11'b11111110100;
    W_iz[3][35] = 11'b11111111010;
    W_iz[3][36] = 11'b00000001000;
    W_iz[3][37] = 11'b00000000000;
    W_iz[3][38] = 11'b00000000110;
    W_iz[3][39] = 11'b11111110111;
    W_iz[3][40] = 11'b00000000000;
    W_iz[3][41] = 11'b11111111000;
    W_iz[3][42] = 11'b11111110111;
    W_iz[3][43] = 11'b11111110111;
    W_iz[3][44] = 11'b11111111011;
    W_iz[3][45] = 11'b00000000001;
    W_iz[3][46] = 11'b00000010010;
    W_iz[3][47] = 11'b11111111011;
    W_iz[3][48] = 11'b11111111111;
    W_iz[3][49] = 11'b11111111011;
    W_iz[3][50] = 11'b11111111000;
    W_iz[3][51] = 11'b00000001100;
    W_iz[3][52] = 11'b11111110111;
    W_iz[3][53] = 11'b00000000011;
    W_iz[3][54] = 11'b00000001001;
    W_iz[3][55] = 11'b00000000001;
    W_iz[3][56] = 11'b00000010010;
    W_iz[3][57] = 11'b00000000010;
    W_iz[3][58] = 11'b00000010011;
    W_iz[3][59] = 11'b00000000011;
    W_iz[3][60] = 11'b11111111000;
    W_iz[3][61] = 11'b00000001001;
    W_iz[3][62] = 11'b00000001100;
    W_iz[3][63] = 11'b11111111000;
    W_iz[4][0] = 11'b11111111100;
    W_iz[4][1] = 11'b00000000010;
    W_iz[4][2] = 11'b11111111110;
    W_iz[4][3] = 11'b00000000100;
    W_iz[4][4] = 11'b11111111111;
    W_iz[4][5] = 11'b11111111110;
    W_iz[4][6] = 11'b11111111001;
    W_iz[4][7] = 11'b11111111100;
    W_iz[4][8] = 11'b11111111110;
    W_iz[4][9] = 11'b00000000101;
    W_iz[4][10] = 11'b00000000010;
    W_iz[4][11] = 11'b00000000111;
    W_iz[4][12] = 11'b11111111110;
    W_iz[4][13] = 11'b00000000100;
    W_iz[4][14] = 11'b00000000100;
    W_iz[4][15] = 11'b00000000010;
    W_iz[4][16] = 11'b11111111111;
    W_iz[4][17] = 11'b00000000101;
    W_iz[4][18] = 11'b00000001000;
    W_iz[4][19] = 11'b00000000100;
    W_iz[4][20] = 11'b11111111111;
    W_iz[4][21] = 11'b00000000001;
    W_iz[4][22] = 11'b00000000110;
    W_iz[4][23] = 11'b00000000001;
    W_iz[4][24] = 11'b00000000000;
    W_iz[4][25] = 11'b11111111111;
    W_iz[4][26] = 11'b11111111001;
    W_iz[4][27] = 11'b00000000010;
    W_iz[4][28] = 11'b00000000100;
    W_iz[4][29] = 11'b00000000000;
    W_iz[4][30] = 11'b00000000101;
    W_iz[4][31] = 11'b00000000100;
    W_iz[4][32] = 11'b11111111111;
    W_iz[4][33] = 11'b11111111011;
    W_iz[4][34] = 11'b11111111010;
    W_iz[4][35] = 11'b11111111101;
    W_iz[4][36] = 11'b11111111101;
    W_iz[4][37] = 11'b11111110110;
    W_iz[4][38] = 11'b00000000010;
    W_iz[4][39] = 11'b11111111111;
    W_iz[4][40] = 11'b11111111111;
    W_iz[4][41] = 11'b00000000111;
    W_iz[4][42] = 11'b11111111011;
    W_iz[4][43] = 11'b00000000100;
    W_iz[4][44] = 11'b00000000000;
    W_iz[4][45] = 11'b11111111100;
    W_iz[4][46] = 11'b11111111011;
    W_iz[4][47] = 11'b00000000101;
    W_iz[4][48] = 11'b00000000010;
    W_iz[4][49] = 11'b00000001001;
    W_iz[4][50] = 11'b00000000000;
    W_iz[4][51] = 11'b00000000010;
    W_iz[4][52] = 11'b11111111110;
    W_iz[4][53] = 11'b11111111010;
    W_iz[4][54] = 11'b11111111001;
    W_iz[4][55] = 11'b11111111101;
    W_iz[4][56] = 11'b00000000111;
    W_iz[4][57] = 11'b11111111110;
    W_iz[4][58] = 11'b00000001000;
    W_iz[4][59] = 11'b11111111110;
    W_iz[4][60] = 11'b11111110111;
    W_iz[4][61] = 11'b11111110010;
    W_iz[4][62] = 11'b11111110000;
    W_iz[4][63] = 11'b00000000011;
    W_iz[5][0] = 11'b00000000110;
    W_iz[5][1] = 11'b00000000010;
    W_iz[5][2] = 11'b00000000001;
    W_iz[5][3] = 11'b00000000000;
    W_iz[5][4] = 11'b00000000001;
    W_iz[5][5] = 11'b00000000101;
    W_iz[5][6] = 11'b11111111010;
    W_iz[5][7] = 11'b11111111011;
    W_iz[5][8] = 11'b00000000000;
    W_iz[5][9] = 11'b00000001000;
    W_iz[5][10] = 11'b00000000100;
    W_iz[5][11] = 11'b11111111000;
    W_iz[5][12] = 11'b11111111011;
    W_iz[5][13] = 11'b00000000101;
    W_iz[5][14] = 11'b11111111110;
    W_iz[5][15] = 11'b00000000110;
    W_iz[5][16] = 11'b11111111000;
    W_iz[5][17] = 11'b00000000100;
    W_iz[5][18] = 11'b00000001001;
    W_iz[5][19] = 11'b11111111011;
    W_iz[5][20] = 11'b11111111011;
    W_iz[5][21] = 11'b11111111001;
    W_iz[5][22] = 11'b00000000100;
    W_iz[5][23] = 11'b00000001010;
    W_iz[5][24] = 11'b00000000100;
    W_iz[5][25] = 11'b11111111100;
    W_iz[5][26] = 11'b11111111101;
    W_iz[5][27] = 11'b11111111100;
    W_iz[5][28] = 11'b11111111101;
    W_iz[5][29] = 11'b11111111010;
    W_iz[5][30] = 11'b11111111110;
    W_iz[5][31] = 11'b11111111010;
    W_iz[5][32] = 11'b00000000101;
    W_iz[5][33] = 11'b11111111110;
    W_iz[5][34] = 11'b11111111100;
    W_iz[5][35] = 11'b00000000101;
    W_iz[5][36] = 11'b11111110111;
    W_iz[5][37] = 11'b00000000001;
    W_iz[5][38] = 11'b00000000000;
    W_iz[5][39] = 11'b11111111100;
    W_iz[5][40] = 11'b00000000110;
    W_iz[5][41] = 11'b00000000011;
    W_iz[5][42] = 11'b00000000111;
    W_iz[5][43] = 11'b00000000110;
    W_iz[5][44] = 11'b00000000000;
    W_iz[5][45] = 11'b00000000111;
    W_iz[5][46] = 11'b00000000010;
    W_iz[5][47] = 11'b11111111110;
    W_iz[5][48] = 11'b11111111010;
    W_iz[5][49] = 11'b11111111111;
    W_iz[5][50] = 11'b11111111101;
    W_iz[5][51] = 11'b00000000100;
    W_iz[5][52] = 11'b00000000101;
    W_iz[5][53] = 11'b00000000011;
    W_iz[5][54] = 11'b11111111000;
    W_iz[5][55] = 11'b00000001010;
    W_iz[5][56] = 11'b00000000101;
    W_iz[5][57] = 11'b11111111110;
    W_iz[5][58] = 11'b11111111111;
    W_iz[5][59] = 11'b00000000111;
    W_iz[5][60] = 11'b11111110111;
    W_iz[5][61] = 11'b00000000000;
    W_iz[5][62] = 11'b11111111101;
    W_iz[5][63] = 11'b11111111101;
    W_iz[6][0] = 11'b00000000011;
    W_iz[6][1] = 11'b00000000100;
    W_iz[6][2] = 11'b11111111111;
    W_iz[6][3] = 11'b00000000010;
    W_iz[6][4] = 11'b00000000110;
    W_iz[6][5] = 11'b00000000011;
    W_iz[6][6] = 11'b11111110111;
    W_iz[6][7] = 11'b00000000011;
    W_iz[6][8] = 11'b11111110100;
    W_iz[6][9] = 11'b11111111110;
    W_iz[6][10] = 11'b00000000000;
    W_iz[6][11] = 11'b11111111100;
    W_iz[6][12] = 11'b11111111001;
    W_iz[6][13] = 11'b00000000011;
    W_iz[6][14] = 11'b00000000000;
    W_iz[6][15] = 11'b11111110101;
    W_iz[6][16] = 11'b00000000100;
    W_iz[6][17] = 11'b00000000101;
    W_iz[6][18] = 11'b11111110100;
    W_iz[6][19] = 11'b11111111000;
    W_iz[6][20] = 11'b00000000111;
    W_iz[6][21] = 11'b11111111010;
    W_iz[6][22] = 11'b00000000011;
    W_iz[6][23] = 11'b11111111010;
    W_iz[6][24] = 11'b00000000011;
    W_iz[6][25] = 11'b11111111011;
    W_iz[6][26] = 11'b00000001001;
    W_iz[6][27] = 11'b11111111110;
    W_iz[6][28] = 11'b00000000110;
    W_iz[6][29] = 11'b00000001001;
    W_iz[6][30] = 11'b11111111111;
    W_iz[6][31] = 11'b00000000000;
    W_iz[6][32] = 11'b00000001011;
    W_iz[6][33] = 11'b11111111000;
    W_iz[6][34] = 11'b11111111000;
    W_iz[6][35] = 11'b11111111100;
    W_iz[6][36] = 11'b00000001010;
    W_iz[6][37] = 11'b00000001000;
    W_iz[6][38] = 11'b11111111011;
    W_iz[6][39] = 11'b11111110101;
    W_iz[6][40] = 11'b00000000100;
    W_iz[6][41] = 11'b11111111111;
    W_iz[6][42] = 11'b11111111000;
    W_iz[6][43] = 11'b00000000001;
    W_iz[6][44] = 11'b11111111101;
    W_iz[6][45] = 11'b00000000101;
    W_iz[6][46] = 11'b11111111110;
    W_iz[6][47] = 11'b11111111110;
    W_iz[6][48] = 11'b11111111101;
    W_iz[6][49] = 11'b00000000000;
    W_iz[6][50] = 11'b11111111000;
    W_iz[6][51] = 11'b11111111101;
    W_iz[6][52] = 11'b11111111000;
    W_iz[6][53] = 11'b00000000111;
    W_iz[6][54] = 11'b11111111111;
    W_iz[6][55] = 11'b11111111100;
    W_iz[6][56] = 11'b11111111101;
    W_iz[6][57] = 11'b00000000111;
    W_iz[6][58] = 11'b00000001000;
    W_iz[6][59] = 11'b00000001010;
    W_iz[6][60] = 11'b00000001111;
    W_iz[6][61] = 11'b00000001010;
    W_iz[6][62] = 11'b00000010001;
    W_iz[6][63] = 11'b00000001101;
    W_iz[7][0] = 11'b11111110101;
    W_iz[7][1] = 11'b00000001000;
    W_iz[7][2] = 11'b00000000001;
    W_iz[7][3] = 11'b00000001001;
    W_iz[7][4] = 11'b11111110110;
    W_iz[7][5] = 11'b00000000010;
    W_iz[7][6] = 11'b11111110111;
    W_iz[7][7] = 11'b00000000101;
    W_iz[7][8] = 11'b11111110010;
    W_iz[7][9] = 11'b11111110101;
    W_iz[7][10] = 11'b00000001001;
    W_iz[7][11] = 11'b11111110101;
    W_iz[7][12] = 11'b11111110101;
    W_iz[7][13] = 11'b00000000101;
    W_iz[7][14] = 11'b00000000100;
    W_iz[7][15] = 11'b00000000100;
    W_iz[7][16] = 11'b00000001011;
    W_iz[7][17] = 11'b11111111110;
    W_iz[7][18] = 11'b00000000000;
    W_iz[7][19] = 11'b00000001101;
    W_iz[7][20] = 11'b11111111110;
    W_iz[7][21] = 11'b11111111000;
    W_iz[7][22] = 11'b11111111101;
    W_iz[7][23] = 11'b11111111100;
    W_iz[7][24] = 11'b11111110110;
    W_iz[7][25] = 11'b11111111110;
    W_iz[7][26] = 11'b11111111000;
    W_iz[7][27] = 11'b11111110110;
    W_iz[7][28] = 11'b00000001101;
    W_iz[7][29] = 11'b00000000100;
    W_iz[7][30] = 11'b00000000001;
    W_iz[7][31] = 11'b00000000111;
    W_iz[7][32] = 11'b00000000100;
    W_iz[7][33] = 11'b11111111110;
    W_iz[7][34] = 11'b00000000111;
    W_iz[7][35] = 11'b00000000100;
    W_iz[7][36] = 11'b11111110111;
    W_iz[7][37] = 11'b11111110110;
    W_iz[7][38] = 11'b00000000100;
    W_iz[7][39] = 11'b00000000000;
    W_iz[7][40] = 11'b11111110100;
    W_iz[7][41] = 11'b11111110110;
    W_iz[7][42] = 11'b00000001000;
    W_iz[7][43] = 11'b00000000001;
    W_iz[7][44] = 11'b00000000011;
    W_iz[7][45] = 11'b00000001100;
    W_iz[7][46] = 11'b11111111111;
    W_iz[7][47] = 11'b00000001010;
    W_iz[7][48] = 11'b00000000001;
    W_iz[7][49] = 11'b11111111111;
    W_iz[7][50] = 11'b11111111011;
    W_iz[7][51] = 11'b00000000110;
    W_iz[7][52] = 11'b11111111110;
    W_iz[7][53] = 11'b11111110110;
    W_iz[7][54] = 11'b00000001100;
    W_iz[7][55] = 11'b00000000010;
    W_iz[7][56] = 11'b11111111010;
    W_iz[7][57] = 11'b00000000110;
    W_iz[7][58] = 11'b11111111011;
    W_iz[7][59] = 11'b00000001011;
    W_iz[7][60] = 11'b00000001011;
    W_iz[7][61] = 11'b00000000011;
    W_iz[7][62] = 11'b00000000001;
    W_iz[7][63] = 11'b00000001001;
    W_iz[8][0] = 11'b00000000011;
    W_iz[8][1] = 11'b00000000101;
    W_iz[8][2] = 11'b00000000100;
    W_iz[8][3] = 11'b00000000100;
    W_iz[8][4] = 11'b11111111110;
    W_iz[8][5] = 11'b11111111011;
    W_iz[8][6] = 11'b00000000100;
    W_iz[8][7] = 11'b00000000010;
    W_iz[8][8] = 11'b11111111001;
    W_iz[8][9] = 11'b00000000001;
    W_iz[8][10] = 11'b00000001000;
    W_iz[8][11] = 11'b00000000000;
    W_iz[8][12] = 11'b00000000101;
    W_iz[8][13] = 11'b00000000001;
    W_iz[8][14] = 11'b00000000001;
    W_iz[8][15] = 11'b00000000110;
    W_iz[8][16] = 11'b11111111111;
    W_iz[8][17] = 11'b00000000111;
    W_iz[8][18] = 11'b11111111111;
    W_iz[8][19] = 11'b00000000101;
    W_iz[8][20] = 11'b11111111111;
    W_iz[8][21] = 11'b00000000100;
    W_iz[8][22] = 11'b00000000011;
    W_iz[8][23] = 11'b00000000011;
    W_iz[8][24] = 11'b11111111011;
    W_iz[8][25] = 11'b00000000100;
    W_iz[8][26] = 11'b00000000100;
    W_iz[8][27] = 11'b00000000011;
    W_iz[8][28] = 11'b00000000111;
    W_iz[8][29] = 11'b11111111001;
    W_iz[8][30] = 11'b11111111110;
    W_iz[8][31] = 11'b00000000011;
    W_iz[8][32] = 11'b00000000010;
    W_iz[8][33] = 11'b00000000100;
    W_iz[8][34] = 11'b00000000100;
    W_iz[8][35] = 11'b00000000001;
    W_iz[8][36] = 11'b00000001000;
    W_iz[8][37] = 11'b00000000011;
    W_iz[8][38] = 11'b11111111110;
    W_iz[8][39] = 11'b00000000010;
    W_iz[8][40] = 11'b00000000101;
    W_iz[8][41] = 11'b11111111010;
    W_iz[8][42] = 11'b00000000010;
    W_iz[8][43] = 11'b11111111101;
    W_iz[8][44] = 11'b00000000000;
    W_iz[8][45] = 11'b11111111100;
    W_iz[8][46] = 11'b11111111010;
    W_iz[8][47] = 11'b00000000111;
    W_iz[8][48] = 11'b11111111110;
    W_iz[8][49] = 11'b11111111101;
    W_iz[8][50] = 11'b11111111111;
    W_iz[8][51] = 11'b00000000000;
    W_iz[8][52] = 11'b11111111001;
    W_iz[8][53] = 11'b11111111101;
    W_iz[8][54] = 11'b00000000010;
    W_iz[8][55] = 11'b11111111101;
    W_iz[8][56] = 11'b00000000101;
    W_iz[8][57] = 11'b11111111101;
    W_iz[8][58] = 11'b11111111101;
    W_iz[8][59] = 11'b00000000100;
    W_iz[8][60] = 11'b11111111011;
    W_iz[8][61] = 11'b11111111010;
    W_iz[8][62] = 11'b11111111010;
    W_iz[8][63] = 11'b00000000100;
    W_iz[9][0] = 11'b11111111100;
    W_iz[9][1] = 11'b11111111101;
    W_iz[9][2] = 11'b00000000110;
    W_iz[9][3] = 11'b00000000101;
    W_iz[9][4] = 11'b00000000001;
    W_iz[9][5] = 11'b00000000010;
    W_iz[9][6] = 11'b00000000010;
    W_iz[9][7] = 11'b00000000001;
    W_iz[9][8] = 11'b00000000001;
    W_iz[9][9] = 11'b00000000001;
    W_iz[9][10] = 11'b11111111111;
    W_iz[9][11] = 11'b00000000000;
    W_iz[9][12] = 11'b00000000001;
    W_iz[9][13] = 11'b00000000100;
    W_iz[9][14] = 11'b11111111011;
    W_iz[9][15] = 11'b00000000001;
    W_iz[9][16] = 11'b00000000000;
    W_iz[9][17] = 11'b00000000000;
    W_iz[9][18] = 11'b00000000000;
    W_iz[9][19] = 11'b11111111101;
    W_iz[9][20] = 11'b00000000000;
    W_iz[9][21] = 11'b00000000001;
    W_iz[9][22] = 11'b11111111110;
    W_iz[9][23] = 11'b11111111101;
    W_iz[9][24] = 11'b00000000000;
    W_iz[9][25] = 11'b00000000110;
    W_iz[9][26] = 11'b11111111010;
    W_iz[9][27] = 11'b11111111010;
    W_iz[9][28] = 11'b00000000111;
    W_iz[9][29] = 11'b00000000010;
    W_iz[9][30] = 11'b00000000000;
    W_iz[9][31] = 11'b00000000000;
    W_iz[9][32] = 11'b11111111100;
    W_iz[9][33] = 11'b00000000000;
    W_iz[9][34] = 11'b11111111111;
    W_iz[9][35] = 11'b00000000000;
    W_iz[9][36] = 11'b00000000010;
    W_iz[9][37] = 11'b00000000001;
    W_iz[9][38] = 11'b00000000010;
    W_iz[9][39] = 11'b00000000100;
    W_iz[9][40] = 11'b00000000010;
    W_iz[9][41] = 11'b00000000000;
    W_iz[9][42] = 11'b00000000000;
    W_iz[9][43] = 11'b00000000010;
    W_iz[9][44] = 11'b00000000001;
    W_iz[9][45] = 11'b00000000010;
    W_iz[9][46] = 11'b00000000000;
    W_iz[9][47] = 11'b11111111111;
    W_iz[9][48] = 11'b11111111111;
    W_iz[9][49] = 11'b11111111001;
    W_iz[9][50] = 11'b00000000100;
    W_iz[9][51] = 11'b00000000101;
    W_iz[9][52] = 11'b11111111110;
    W_iz[9][53] = 11'b11111111101;
    W_iz[9][54] = 11'b11111111101;
    W_iz[9][55] = 11'b11111111101;
    W_iz[9][56] = 11'b11111111110;
    W_iz[9][57] = 11'b00000000110;
    W_iz[9][58] = 11'b00000000100;
    W_iz[9][59] = 11'b11111111100;
    W_iz[9][60] = 11'b11111111111;
    W_iz[9][61] = 11'b11111111110;
    W_iz[9][62] = 11'b00000000101;
    W_iz[9][63] = 11'b11111111101;
    W_iz[10][0] = 11'b11111111101;
    W_iz[10][1] = 11'b11111111110;
    W_iz[10][2] = 11'b11111111001;
    W_iz[10][3] = 11'b11111111100;
    W_iz[10][4] = 11'b11111111110;
    W_iz[10][5] = 11'b11111111111;
    W_iz[10][6] = 11'b00000000001;
    W_iz[10][7] = 11'b11111111011;
    W_iz[10][8] = 11'b11111111111;
    W_iz[10][9] = 11'b11111111111;
    W_iz[10][10] = 11'b11111111111;
    W_iz[10][11] = 11'b11111111001;
    W_iz[10][12] = 11'b11111111111;
    W_iz[10][13] = 11'b00000000010;
    W_iz[10][14] = 11'b11111111111;
    W_iz[10][15] = 11'b00000000011;
    W_iz[10][16] = 11'b11111111011;
    W_iz[10][17] = 11'b00000000111;
    W_iz[10][18] = 11'b00000000000;
    W_iz[10][19] = 11'b00000000010;
    W_iz[10][20] = 11'b00000000010;
    W_iz[10][21] = 11'b11111111110;
    W_iz[10][22] = 11'b00000000100;
    W_iz[10][23] = 11'b00000000111;
    W_iz[10][24] = 11'b00000000011;
    W_iz[10][25] = 11'b00000000001;
    W_iz[10][26] = 11'b00000000000;
    W_iz[10][27] = 11'b11111111001;
    W_iz[10][28] = 11'b11111111110;
    W_iz[10][29] = 11'b00000001000;
    W_iz[10][30] = 11'b11111111101;
    W_iz[10][31] = 11'b11111111101;
    W_iz[10][32] = 11'b00000000000;
    W_iz[10][33] = 11'b00000000011;
    W_iz[10][34] = 11'b11111111111;
    W_iz[10][35] = 11'b11111111110;
    W_iz[10][36] = 11'b00000000000;
    W_iz[10][37] = 11'b00000000001;
    W_iz[10][38] = 11'b00000000100;
    W_iz[10][39] = 11'b00000000000;
    W_iz[10][40] = 11'b00000000100;
    W_iz[10][41] = 11'b11111111110;
    W_iz[10][42] = 11'b00000000100;
    W_iz[10][43] = 11'b00000000000;
    W_iz[10][44] = 11'b00000000001;
    W_iz[10][45] = 11'b00000000010;
    W_iz[10][46] = 11'b00000000010;
    W_iz[10][47] = 11'b00000000001;
    W_iz[10][48] = 11'b00000000010;
    W_iz[10][49] = 11'b00000000001;
    W_iz[10][50] = 11'b11111111100;
    W_iz[10][51] = 11'b00000000011;
    W_iz[10][52] = 11'b00000000011;
    W_iz[10][53] = 11'b00000000010;
    W_iz[10][54] = 11'b11111111001;
    W_iz[10][55] = 11'b00000000010;
    W_iz[10][56] = 11'b00000000010;
    W_iz[10][57] = 11'b11111111011;
    W_iz[10][58] = 11'b11111111100;
    W_iz[10][59] = 11'b11111111101;
    W_iz[10][60] = 11'b00000000101;
    W_iz[10][61] = 11'b00000000010;
    W_iz[10][62] = 11'b00000000101;
    W_iz[10][63] = 11'b00000001001;
    W_iz[11][0] = 11'b00000000000;
    W_iz[11][1] = 11'b00000001000;
    W_iz[11][2] = 11'b00000000000;
    W_iz[11][3] = 11'b00000000110;
    W_iz[11][4] = 11'b11111111010;
    W_iz[11][5] = 11'b00000000001;
    W_iz[11][6] = 11'b00000000001;
    W_iz[11][7] = 11'b11111111110;
    W_iz[11][8] = 11'b11111111111;
    W_iz[11][9] = 11'b00000000101;
    W_iz[11][10] = 11'b11111111100;
    W_iz[11][11] = 11'b11111111111;
    W_iz[11][12] = 11'b11111111100;
    W_iz[11][13] = 11'b11111111111;
    W_iz[11][14] = 11'b11111111110;
    W_iz[11][15] = 11'b11111111111;
    W_iz[11][16] = 11'b00000000000;
    W_iz[11][17] = 11'b00000000001;
    W_iz[11][18] = 11'b11111111101;
    W_iz[11][19] = 11'b00000000100;
    W_iz[11][20] = 11'b11111111110;
    W_iz[11][21] = 11'b00000000010;
    W_iz[11][22] = 11'b00000000011;
    W_iz[11][23] = 11'b00000000010;
    W_iz[11][24] = 11'b00000000111;
    W_iz[11][25] = 11'b00000000001;
    W_iz[11][26] = 11'b11111111111;
    W_iz[11][27] = 11'b11111111110;
    W_iz[11][28] = 11'b00000000001;
    W_iz[11][29] = 11'b00000000001;
    W_iz[11][30] = 11'b11111111100;
    W_iz[11][31] = 11'b00000001000;
    W_iz[11][32] = 11'b00000000100;
    W_iz[11][33] = 11'b11111111011;
    W_iz[11][34] = 11'b00000000010;
    W_iz[11][35] = 11'b00000000001;
    W_iz[11][36] = 11'b00000000001;
    W_iz[11][37] = 11'b11111111001;
    W_iz[11][38] = 11'b00000000011;
    W_iz[11][39] = 11'b00000000000;
    W_iz[11][40] = 11'b00000000000;
    W_iz[11][41] = 11'b00000000101;
    W_iz[11][42] = 11'b11111111011;
    W_iz[11][43] = 11'b00000000001;
    W_iz[11][44] = 11'b11111111101;
    W_iz[11][45] = 11'b11111111110;
    W_iz[11][46] = 11'b00000000110;
    W_iz[11][47] = 11'b11111111101;
    W_iz[11][48] = 11'b11111111110;
    W_iz[11][49] = 11'b11111111111;
    W_iz[11][50] = 11'b11111111100;
    W_iz[11][51] = 11'b11111111101;
    W_iz[11][52] = 11'b11111111101;
    W_iz[11][53] = 11'b11111111100;
    W_iz[11][54] = 11'b11111111110;
    W_iz[11][55] = 11'b11111111001;
    W_iz[11][56] = 11'b11111111101;
    W_iz[11][57] = 11'b00000000100;
    W_iz[11][58] = 11'b11111111100;
    W_iz[11][59] = 11'b11111111101;
    W_iz[11][60] = 11'b11111111101;
    W_iz[11][61] = 11'b11111111101;
    W_iz[11][62] = 11'b11111111010;
    W_iz[11][63] = 11'b11111111110;
    W_iz[12][0] = 11'b00000000000;
    W_iz[12][1] = 11'b11111111110;
    W_iz[12][2] = 11'b11111111111;
    W_iz[12][3] = 11'b11111111101;
    W_iz[12][4] = 11'b00000000000;
    W_iz[12][5] = 11'b00000000011;
    W_iz[12][6] = 11'b11111111100;
    W_iz[12][7] = 11'b11111111011;
    W_iz[12][8] = 11'b11111111001;
    W_iz[12][9] = 11'b11111111101;
    W_iz[12][10] = 11'b11111111001;
    W_iz[12][11] = 11'b11111111110;
    W_iz[12][12] = 11'b11111111111;
    W_iz[12][13] = 11'b00000000011;
    W_iz[12][14] = 11'b00000000001;
    W_iz[12][15] = 11'b11111111111;
    W_iz[12][16] = 11'b11111111100;
    W_iz[12][17] = 11'b11111111101;
    W_iz[12][18] = 11'b11111111100;
    W_iz[12][19] = 11'b11111111011;
    W_iz[12][20] = 11'b11111111111;
    W_iz[12][21] = 11'b00000000011;
    W_iz[12][22] = 11'b00000001000;
    W_iz[12][23] = 11'b00000000101;
    W_iz[12][24] = 11'b11111111001;
    W_iz[12][25] = 11'b11111111010;
    W_iz[12][26] = 11'b00000000000;
    W_iz[12][27] = 11'b11111111001;
    W_iz[12][28] = 11'b00000000110;
    W_iz[12][29] = 11'b00000000000;
    W_iz[12][30] = 11'b00000000110;
    W_iz[12][31] = 11'b11111111100;
    W_iz[12][32] = 11'b11111111001;
    W_iz[12][33] = 11'b11111111010;
    W_iz[12][34] = 11'b11111111100;
    W_iz[12][35] = 11'b11111111100;
    W_iz[12][36] = 11'b11111111010;
    W_iz[12][37] = 11'b11111111011;
    W_iz[12][38] = 11'b11111111101;
    W_iz[12][39] = 11'b00000000010;
    W_iz[12][40] = 11'b00000000001;
    W_iz[12][41] = 11'b11111111100;
    W_iz[12][42] = 11'b11111111111;
    W_iz[12][43] = 11'b11111111101;
    W_iz[12][44] = 11'b11111111000;
    W_iz[12][45] = 11'b11111111111;
    W_iz[12][46] = 11'b11111111111;
    W_iz[12][47] = 11'b11111111111;
    W_iz[12][48] = 11'b00000000000;
    W_iz[12][49] = 11'b11111111110;
    W_iz[12][50] = 11'b00000000101;
    W_iz[12][51] = 11'b11111111101;
    W_iz[12][52] = 11'b00000000111;
    W_iz[12][53] = 11'b00000000100;
    W_iz[12][54] = 11'b00000001000;
    W_iz[12][55] = 11'b00000000110;
    W_iz[12][56] = 11'b00000000011;
    W_iz[12][57] = 11'b11111111001;
    W_iz[12][58] = 11'b00000000100;
    W_iz[12][59] = 11'b00000001110;
    W_iz[12][60] = 11'b00000001010;
    W_iz[12][61] = 11'b00000001011;
    W_iz[12][62] = 11'b00000001101;
    W_iz[12][63] = 11'b00000001100;
    W_iz[13][0] = 11'b00000000001;
    W_iz[13][1] = 11'b00000000001;
    W_iz[13][2] = 11'b00000000010;
    W_iz[13][3] = 11'b11111111111;
    W_iz[13][4] = 11'b11111111111;
    W_iz[13][5] = 11'b11111111011;
    W_iz[13][6] = 11'b00000000110;
    W_iz[13][7] = 11'b11111111001;
    W_iz[13][8] = 11'b11111111010;
    W_iz[13][9] = 11'b11111111110;
    W_iz[13][10] = 11'b00000000000;
    W_iz[13][11] = 11'b11111111111;
    W_iz[13][12] = 11'b11111111100;
    W_iz[13][13] = 11'b11111111111;
    W_iz[13][14] = 11'b11111111100;
    W_iz[13][15] = 11'b11111111100;
    W_iz[13][16] = 11'b00000000101;
    W_iz[13][17] = 11'b11111111011;
    W_iz[13][18] = 11'b00000000001;
    W_iz[13][19] = 11'b11111111010;
    W_iz[13][20] = 11'b11111111111;
    W_iz[13][21] = 11'b00000000000;
    W_iz[13][22] = 11'b00000000011;
    W_iz[13][23] = 11'b00000000010;
    W_iz[13][24] = 11'b11111111111;
    W_iz[13][25] = 11'b11111111101;
    W_iz[13][26] = 11'b11111111111;
    W_iz[13][27] = 11'b00000000011;
    W_iz[13][28] = 11'b00000000001;
    W_iz[13][29] = 11'b11111111100;
    W_iz[13][30] = 11'b11111111110;
    W_iz[13][31] = 11'b11111111001;
    W_iz[13][32] = 11'b00000000000;
    W_iz[13][33] = 11'b11111111000;
    W_iz[13][34] = 11'b11111111110;
    W_iz[13][35] = 11'b00000000100;
    W_iz[13][36] = 11'b11111111100;
    W_iz[13][37] = 11'b11111111010;
    W_iz[13][38] = 11'b11111110111;
    W_iz[13][39] = 11'b00000000101;
    W_iz[13][40] = 11'b11111111101;
    W_iz[13][41] = 11'b11111111111;
    W_iz[13][42] = 11'b00000000000;
    W_iz[13][43] = 11'b11111111101;
    W_iz[13][44] = 11'b00000000001;
    W_iz[13][45] = 11'b11111111101;
    W_iz[13][46] = 11'b11111111111;
    W_iz[13][47] = 11'b00000000100;
    W_iz[13][48] = 11'b00000000010;
    W_iz[13][49] = 11'b00000000010;
    W_iz[13][50] = 11'b00000000001;
    W_iz[13][51] = 11'b00000000001;
    W_iz[13][52] = 11'b11111111110;
    W_iz[13][53] = 11'b11111111101;
    W_iz[13][54] = 11'b00000000010;
    W_iz[13][55] = 11'b00000000000;
    W_iz[13][56] = 11'b00000000001;
    W_iz[13][57] = 11'b11111111011;
    W_iz[13][58] = 11'b11111111100;
    W_iz[13][59] = 11'b11111111110;
    W_iz[13][60] = 11'b00000000111;
    W_iz[13][61] = 11'b00000000101;
    W_iz[13][62] = 11'b11111111110;
    W_iz[13][63] = 11'b00000000101;
    W_iz[14][0] = 11'b00000000110;
    W_iz[14][1] = 11'b11111111110;
    W_iz[14][2] = 11'b00000001001;
    W_iz[14][3] = 11'b11111111110;
    W_iz[14][4] = 11'b00000000101;
    W_iz[14][5] = 11'b00000000001;
    W_iz[14][6] = 11'b11111111001;
    W_iz[14][7] = 11'b00000001001;
    W_iz[14][8] = 11'b00000001011;
    W_iz[14][9] = 11'b00000000110;
    W_iz[14][10] = 11'b00000001000;
    W_iz[14][11] = 11'b00000000000;
    W_iz[14][12] = 11'b00000000000;
    W_iz[14][13] = 11'b00000000010;
    W_iz[14][14] = 11'b11111111110;
    W_iz[14][15] = 11'b11111111001;
    W_iz[14][16] = 11'b11111111101;
    W_iz[14][17] = 11'b00000000101;
    W_iz[14][18] = 11'b00000000000;
    W_iz[14][19] = 11'b00000000000;
    W_iz[14][20] = 11'b11111111111;
    W_iz[14][21] = 11'b11111111011;
    W_iz[14][22] = 11'b00000001001;
    W_iz[14][23] = 11'b00000000000;
    W_iz[14][24] = 11'b11111111011;
    W_iz[14][25] = 11'b00000000011;
    W_iz[14][26] = 11'b11111111010;
    W_iz[14][27] = 11'b11111111100;
    W_iz[14][28] = 11'b00000000110;
    W_iz[14][29] = 11'b00000000101;
    W_iz[14][30] = 11'b11111111011;
    W_iz[14][31] = 11'b00000000101;
    W_iz[14][32] = 11'b00000000000;
    W_iz[14][33] = 11'b00000000011;
    W_iz[14][34] = 11'b00000000111;
    W_iz[14][35] = 11'b00000001000;
    W_iz[14][36] = 11'b11111111111;
    W_iz[14][37] = 11'b00000000010;
    W_iz[14][38] = 11'b11111111000;
    W_iz[14][39] = 11'b11111111111;
    W_iz[14][40] = 11'b00000000100;
    W_iz[14][41] = 11'b11111111101;
    W_iz[14][42] = 11'b00000001001;
    W_iz[14][43] = 11'b00000000010;
    W_iz[14][44] = 11'b00000000100;
    W_iz[14][45] = 11'b11111111100;
    W_iz[14][46] = 11'b11111111001;
    W_iz[14][47] = 11'b00000001000;
    W_iz[14][48] = 11'b11111111010;
    W_iz[14][49] = 11'b11111111100;
    W_iz[14][50] = 11'b00000000100;
    W_iz[14][51] = 11'b11111111111;
    W_iz[14][52] = 11'b00000000100;
    W_iz[14][53] = 11'b11111110010;
    W_iz[14][54] = 11'b11111111110;
    W_iz[14][55] = 11'b00000000001;
    W_iz[14][56] = 11'b11111111011;
    W_iz[14][57] = 11'b11111111110;
    W_iz[14][58] = 11'b11111111011;
    W_iz[14][59] = 11'b11111111010;
    W_iz[14][60] = 11'b11111111110;
    W_iz[14][61] = 11'b11111110100;
    W_iz[14][62] = 11'b11111110001;
    W_iz[14][63] = 11'b11111110000;
    W_iz[15][0] = 11'b11111110101;
    W_iz[15][1] = 11'b11111110101;
    W_iz[15][2] = 11'b00000000011;
    W_iz[15][3] = 11'b11111111110;
    W_iz[15][4] = 11'b00000000110;
    W_iz[15][5] = 11'b00000001000;
    W_iz[15][6] = 11'b11111111001;
    W_iz[15][7] = 11'b00000000010;
    W_iz[15][8] = 11'b11111111011;
    W_iz[15][9] = 11'b11111110100;
    W_iz[15][10] = 11'b11111111100;
    W_iz[15][11] = 11'b00000000101;
    W_iz[15][12] = 11'b00000000110;
    W_iz[15][13] = 11'b11111111010;
    W_iz[15][14] = 11'b00000000110;
    W_iz[15][15] = 11'b00000000000;
    W_iz[15][16] = 11'b00000000001;
    W_iz[15][17] = 11'b11111111101;
    W_iz[15][18] = 11'b00000000001;
    W_iz[15][19] = 11'b00000000111;
    W_iz[15][20] = 11'b11111111100;
    W_iz[15][21] = 11'b11111111101;
    W_iz[15][22] = 11'b00000001000;
    W_iz[15][23] = 11'b11111111101;
    W_iz[15][24] = 11'b00000000111;
    W_iz[15][25] = 11'b00000000011;
    W_iz[15][26] = 11'b00000000100;
    W_iz[15][27] = 11'b11111111110;
    W_iz[15][28] = 11'b00000000110;
    W_iz[15][29] = 11'b00000001001;
    W_iz[15][30] = 11'b00000000110;
    W_iz[15][31] = 11'b00000000011;
    W_iz[15][32] = 11'b11111111011;
    W_iz[15][33] = 11'b11111111101;
    W_iz[15][34] = 11'b11111110100;
    W_iz[15][35] = 11'b11111111010;
    W_iz[15][36] = 11'b00000001000;
    W_iz[15][37] = 11'b00000000000;
    W_iz[15][38] = 11'b00000000110;
    W_iz[15][39] = 11'b11111110111;
    W_iz[15][40] = 11'b00000000000;
    W_iz[15][41] = 11'b11111111000;
    W_iz[15][42] = 11'b11111110111;
    W_iz[15][43] = 11'b11111110111;
    W_iz[15][44] = 11'b11111111011;
    W_iz[15][45] = 11'b00000000001;
    W_iz[15][46] = 11'b00000010010;
    W_iz[15][47] = 11'b11111111011;
    W_iz[15][48] = 11'b11111111111;
    W_iz[15][49] = 11'b11111111011;
    W_iz[15][50] = 11'b11111111000;
    W_iz[15][51] = 11'b00000001100;
    W_iz[15][52] = 11'b11111110111;
    W_iz[15][53] = 11'b00000000011;
    W_iz[15][54] = 11'b00000001001;
    W_iz[15][55] = 11'b00000000001;
    W_iz[15][56] = 11'b00000010010;
    W_iz[15][57] = 11'b00000000010;
    W_iz[15][58] = 11'b00000010011;
    W_iz[15][59] = 11'b00000000011;
    W_iz[15][60] = 11'b11111111000;
    W_iz[15][61] = 11'b00000001001;
    W_iz[15][62] = 11'b00000001100;
    W_iz[15][63] = 11'b11111111000;

    // Initialize W_in weights
    W_in[0][0] = 11'b11111111100;
    W_in[0][1] = 11'b00000000010;
    W_in[0][2] = 11'b11111111110;
    W_in[0][3] = 11'b00000000100;
    W_in[0][4] = 11'b11111111111;
    W_in[0][5] = 11'b11111111110;
    W_in[0][6] = 11'b11111111001;
    W_in[0][7] = 11'b11111111100;
    W_in[0][8] = 11'b11111111110;
    W_in[0][9] = 11'b00000000101;
    W_in[0][10] = 11'b00000000010;
    W_in[0][11] = 11'b00000000111;
    W_in[0][12] = 11'b11111111110;
    W_in[0][13] = 11'b00000000100;
    W_in[0][14] = 11'b00000000100;
    W_in[0][15] = 11'b00000000010;
    W_in[0][16] = 11'b11111111111;
    W_in[0][17] = 11'b00000000101;
    W_in[0][18] = 11'b00000001000;
    W_in[0][19] = 11'b00000000100;
    W_in[0][20] = 11'b11111111111;
    W_in[0][21] = 11'b00000000001;
    W_in[0][22] = 11'b00000000110;
    W_in[0][23] = 11'b00000000001;
    W_in[0][24] = 11'b00000000000;
    W_in[0][25] = 11'b11111111111;
    W_in[0][26] = 11'b11111111001;
    W_in[0][27] = 11'b00000000010;
    W_in[0][28] = 11'b00000000100;
    W_in[0][29] = 11'b00000000000;
    W_in[0][30] = 11'b00000000101;
    W_in[0][31] = 11'b00000000100;
    W_in[0][32] = 11'b11111111111;
    W_in[0][33] = 11'b11111111011;
    W_in[0][34] = 11'b11111111010;
    W_in[0][35] = 11'b11111111101;
    W_in[0][36] = 11'b11111111101;
    W_in[0][37] = 11'b11111110110;
    W_in[0][38] = 11'b00000000010;
    W_in[0][39] = 11'b11111111111;
    W_in[0][40] = 11'b11111111111;
    W_in[0][41] = 11'b00000000111;
    W_in[0][42] = 11'b11111111011;
    W_in[0][43] = 11'b00000000100;
    W_in[0][44] = 11'b00000000000;
    W_in[0][45] = 11'b11111111100;
    W_in[0][46] = 11'b11111111011;
    W_in[0][47] = 11'b00000000101;
    W_in[0][48] = 11'b00000000010;
    W_in[0][49] = 11'b00000001001;
    W_in[0][50] = 11'b00000000000;
    W_in[0][51] = 11'b00000000010;
    W_in[0][52] = 11'b11111111110;
    W_in[0][53] = 11'b11111111010;
    W_in[0][54] = 11'b11111111001;
    W_in[0][55] = 11'b11111111101;
    W_in[0][56] = 11'b00000000111;
    W_in[0][57] = 11'b11111111110;
    W_in[0][58] = 11'b00000001000;
    W_in[0][59] = 11'b11111111110;
    W_in[0][60] = 11'b11111110111;
    W_in[0][61] = 11'b11111110010;
    W_in[0][62] = 11'b11111110000;
    W_in[0][63] = 11'b00000000011;
    W_in[1][0] = 11'b00000000110;
    W_in[1][1] = 11'b00000000010;
    W_in[1][2] = 11'b00000000001;
    W_in[1][3] = 11'b00000000000;
    W_in[1][4] = 11'b00000000001;
    W_in[1][5] = 11'b00000000101;
    W_in[1][6] = 11'b11111111010;
    W_in[1][7] = 11'b11111111011;
    W_in[1][8] = 11'b00000000000;
    W_in[1][9] = 11'b00000001000;
    W_in[1][10] = 11'b00000000100;
    W_in[1][11] = 11'b11111111000;
    W_in[1][12] = 11'b11111111011;
    W_in[1][13] = 11'b00000000101;
    W_in[1][14] = 11'b11111111110;
    W_in[1][15] = 11'b00000000110;
    W_in[1][16] = 11'b11111111000;
    W_in[1][17] = 11'b00000000100;
    W_in[1][18] = 11'b00000001001;
    W_in[1][19] = 11'b11111111011;
    W_in[1][20] = 11'b11111111011;
    W_in[1][21] = 11'b11111111001;
    W_in[1][22] = 11'b00000000100;
    W_in[1][23] = 11'b00000001010;
    W_in[1][24] = 11'b00000000100;
    W_in[1][25] = 11'b11111111100;
    W_in[1][26] = 11'b11111111101;
    W_in[1][27] = 11'b11111111100;
    W_in[1][28] = 11'b11111111101;
    W_in[1][29] = 11'b11111111010;
    W_in[1][30] = 11'b11111111110;
    W_in[1][31] = 11'b11111111010;
    W_in[1][32] = 11'b00000000101;
    W_in[1][33] = 11'b11111111110;
    W_in[1][34] = 11'b11111111100;
    W_in[1][35] = 11'b00000000101;
    W_in[1][36] = 11'b11111110111;
    W_in[1][37] = 11'b00000000001;
    W_in[1][38] = 11'b00000000000;
    W_in[1][39] = 11'b11111111100;
    W_in[1][40] = 11'b00000000110;
    W_in[1][41] = 11'b00000000011;
    W_in[1][42] = 11'b00000000111;
    W_in[1][43] = 11'b00000000110;
    W_in[1][44] = 11'b00000000000;
    W_in[1][45] = 11'b00000000111;
    W_in[1][46] = 11'b00000000010;
    W_in[1][47] = 11'b11111111110;
    W_in[1][48] = 11'b11111111010;
    W_in[1][49] = 11'b11111111111;
    W_in[1][50] = 11'b11111111101;
    W_in[1][51] = 11'b00000000100;
    W_in[1][52] = 11'b00000000101;
    W_in[1][53] = 11'b00000000011;
    W_in[1][54] = 11'b11111111000;
    W_in[1][55] = 11'b00000001010;
    W_in[1][56] = 11'b00000000101;
    W_in[1][57] = 11'b11111111110;
    W_in[1][58] = 11'b11111111111;
    W_in[1][59] = 11'b00000000111;
    W_in[1][60] = 11'b11111110111;
    W_in[1][61] = 11'b00000000000;
    W_in[1][62] = 11'b11111111101;
    W_in[1][63] = 11'b11111111101;
    W_in[2][0] = 11'b00000000011;
    W_in[2][1] = 11'b00000000100;
    W_in[2][2] = 11'b11111111111;
    W_in[2][3] = 11'b00000000010;
    W_in[2][4] = 11'b00000000110;
    W_in[2][5] = 11'b00000000011;
    W_in[2][6] = 11'b11111110111;
    W_in[2][7] = 11'b00000000011;
    W_in[2][8] = 11'b11111110100;
    W_in[2][9] = 11'b11111111110;
    W_in[2][10] = 11'b00000000000;
    W_in[2][11] = 11'b11111111100;
    W_in[2][12] = 11'b11111111001;
    W_in[2][13] = 11'b00000000011;
    W_in[2][14] = 11'b00000000000;
    W_in[2][15] = 11'b11111110101;
    W_in[2][16] = 11'b00000000100;
    W_in[2][17] = 11'b00000000101;
    W_in[2][18] = 11'b11111110100;
    W_in[2][19] = 11'b11111111000;
    W_in[2][20] = 11'b00000000111;
    W_in[2][21] = 11'b11111111010;
    W_in[2][22] = 11'b00000000011;
    W_in[2][23] = 11'b11111111010;
    W_in[2][24] = 11'b00000000011;
    W_in[2][25] = 11'b11111111011;
    W_in[2][26] = 11'b00000001001;
    W_in[2][27] = 11'b11111111110;
    W_in[2][28] = 11'b00000000110;
    W_in[2][29] = 11'b00000001001;
    W_in[2][30] = 11'b11111111111;
    W_in[2][31] = 11'b00000000000;
    W_in[2][32] = 11'b00000001011;
    W_in[2][33] = 11'b11111111000;
    W_in[2][34] = 11'b11111111000;
    W_in[2][35] = 11'b11111111100;
    W_in[2][36] = 11'b00000001010;
    W_in[2][37] = 11'b00000001000;
    W_in[2][38] = 11'b11111111011;
    W_in[2][39] = 11'b11111110101;
    W_in[2][40] = 11'b00000000100;
    W_in[2][41] = 11'b11111111111;
    W_in[2][42] = 11'b11111111000;
    W_in[2][43] = 11'b00000000001;
    W_in[2][44] = 11'b11111111101;
    W_in[2][45] = 11'b00000000101;
    W_in[2][46] = 11'b11111111110;
    W_in[2][47] = 11'b11111111110;
    W_in[2][48] = 11'b11111111101;
    W_in[2][49] = 11'b00000000000;
    W_in[2][50] = 11'b11111111000;
    W_in[2][51] = 11'b11111111101;
    W_in[2][52] = 11'b11111111000;
    W_in[2][53] = 11'b00000000111;
    W_in[2][54] = 11'b11111111111;
    W_in[2][55] = 11'b11111111100;
    W_in[2][56] = 11'b11111111101;
    W_in[2][57] = 11'b00000000111;
    W_in[2][58] = 11'b00000001000;
    W_in[2][59] = 11'b00000001010;
    W_in[2][60] = 11'b00000001111;
    W_in[2][61] = 11'b00000001010;
    W_in[2][62] = 11'b00000010001;
    W_in[2][63] = 11'b00000001101;
    W_in[3][0] = 11'b11111110101;
    W_in[3][1] = 11'b00000001000;
    W_in[3][2] = 11'b00000000001;
    W_in[3][3] = 11'b00000001001;
    W_in[3][4] = 11'b11111110110;
    W_in[3][5] = 11'b00000000010;
    W_in[3][6] = 11'b11111110111;
    W_in[3][7] = 11'b00000000101;
    W_in[3][8] = 11'b11111110010;
    W_in[3][9] = 11'b11111110101;
    W_in[3][10] = 11'b00000001001;
    W_in[3][11] = 11'b11111110101;
    W_in[3][12] = 11'b11111110101;
    W_in[3][13] = 11'b00000000101;
    W_in[3][14] = 11'b00000000100;
    W_in[3][15] = 11'b00000000100;
    W_in[3][16] = 11'b00000001011;
    W_in[3][17] = 11'b11111111110;
    W_in[3][18] = 11'b00000000000;
    W_in[3][19] = 11'b00000001101;
    W_in[3][20] = 11'b11111111110;
    W_in[3][21] = 11'b11111111000;
    W_in[3][22] = 11'b11111111101;
    W_in[3][23] = 11'b11111111100;
    W_in[3][24] = 11'b11111110110;
    W_in[3][25] = 11'b11111111110;
    W_in[3][26] = 11'b11111111000;
    W_in[3][27] = 11'b11111110110;
    W_in[3][28] = 11'b00000001101;
    W_in[3][29] = 11'b00000000100;
    W_in[3][30] = 11'b00000000001;
    W_in[3][31] = 11'b00000000111;
    W_in[3][32] = 11'b00000000100;
    W_in[3][33] = 11'b11111111110;
    W_in[3][34] = 11'b00000000111;
    W_in[3][35] = 11'b00000000100;
    W_in[3][36] = 11'b11111110111;
    W_in[3][37] = 11'b11111110110;
    W_in[3][38] = 11'b00000000100;
    W_in[3][39] = 11'b00000000000;
    W_in[3][40] = 11'b11111110100;
    W_in[3][41] = 11'b11111110110;
    W_in[3][42] = 11'b00000001000;
    W_in[3][43] = 11'b00000000001;
    W_in[3][44] = 11'b00000000011;
    W_in[3][45] = 11'b00000001100;
    W_in[3][46] = 11'b11111111111;
    W_in[3][47] = 11'b00000001010;
    W_in[3][48] = 11'b00000000001;
    W_in[3][49] = 11'b11111111111;
    W_in[3][50] = 11'b11111111011;
    W_in[3][51] = 11'b00000000110;
    W_in[3][52] = 11'b11111111110;
    W_in[3][53] = 11'b11111110110;
    W_in[3][54] = 11'b00000001100;
    W_in[3][55] = 11'b00000000010;
    W_in[3][56] = 11'b11111111010;
    W_in[3][57] = 11'b00000000110;
    W_in[3][58] = 11'b11111111011;
    W_in[3][59] = 11'b00000001011;
    W_in[3][60] = 11'b00000001011;
    W_in[3][61] = 11'b00000000011;
    W_in[3][62] = 11'b00000000001;
    W_in[3][63] = 11'b00000001001;
    W_in[4][0] = 11'b00000000011;
    W_in[4][1] = 11'b00000000101;
    W_in[4][2] = 11'b00000000100;
    W_in[4][3] = 11'b00000000100;
    W_in[4][4] = 11'b11111111110;
    W_in[4][5] = 11'b11111111011;
    W_in[4][6] = 11'b00000000100;
    W_in[4][7] = 11'b00000000010;
    W_in[4][8] = 11'b11111111001;
    W_in[4][9] = 11'b00000000001;
    W_in[4][10] = 11'b00000001000;
    W_in[4][11] = 11'b00000000000;
    W_in[4][12] = 11'b00000000101;
    W_in[4][13] = 11'b00000000001;
    W_in[4][14] = 11'b00000000001;
    W_in[4][15] = 11'b00000000110;
    W_in[4][16] = 11'b11111111111;
    W_in[4][17] = 11'b00000000111;
    W_in[4][18] = 11'b11111111111;
    W_in[4][19] = 11'b00000000101;
    W_in[4][20] = 11'b11111111111;
    W_in[4][21] = 11'b00000000100;
    W_in[4][22] = 11'b00000000011;
    W_in[4][23] = 11'b00000000011;
    W_in[4][24] = 11'b11111111011;
    W_in[4][25] = 11'b00000000100;
    W_in[4][26] = 11'b00000000100;
    W_in[4][27] = 11'b00000000011;
    W_in[4][28] = 11'b00000000111;
    W_in[4][29] = 11'b11111111001;
    W_in[4][30] = 11'b11111111110;
    W_in[4][31] = 11'b00000000011;
    W_in[4][32] = 11'b00000000010;
    W_in[4][33] = 11'b00000000100;
    W_in[4][34] = 11'b00000000100;
    W_in[4][35] = 11'b00000000001;
    W_in[4][36] = 11'b00000001000;
    W_in[4][37] = 11'b00000000011;
    W_in[4][38] = 11'b11111111110;
    W_in[4][39] = 11'b00000000010;
    W_in[4][40] = 11'b00000000101;
    W_in[4][41] = 11'b11111111010;
    W_in[4][42] = 11'b00000000010;
    W_in[4][43] = 11'b11111111101;
    W_in[4][44] = 11'b00000000000;
    W_in[4][45] = 11'b11111111100;
    W_in[4][46] = 11'b11111111010;
    W_in[4][47] = 11'b00000000111;
    W_in[4][48] = 11'b11111111110;
    W_in[4][49] = 11'b11111111101;
    W_in[4][50] = 11'b11111111111;
    W_in[4][51] = 11'b00000000000;
    W_in[4][52] = 11'b11111111001;
    W_in[4][53] = 11'b11111111101;
    W_in[4][54] = 11'b00000000010;
    W_in[4][55] = 11'b11111111101;
    W_in[4][56] = 11'b00000000101;
    W_in[4][57] = 11'b11111111101;
    W_in[4][58] = 11'b11111111101;
    W_in[4][59] = 11'b00000000100;
    W_in[4][60] = 11'b11111111011;
    W_in[4][61] = 11'b11111111010;
    W_in[4][62] = 11'b11111111010;
    W_in[4][63] = 11'b00000000100;
    W_in[5][0] = 11'b11111111100;
    W_in[5][1] = 11'b11111111101;
    W_in[5][2] = 11'b00000000110;
    W_in[5][3] = 11'b00000000101;
    W_in[5][4] = 11'b00000000001;
    W_in[5][5] = 11'b00000000010;
    W_in[5][6] = 11'b00000000010;
    W_in[5][7] = 11'b00000000001;
    W_in[5][8] = 11'b00000000001;
    W_in[5][9] = 11'b00000000001;
    W_in[5][10] = 11'b11111111111;
    W_in[5][11] = 11'b00000000000;
    W_in[5][12] = 11'b00000000001;
    W_in[5][13] = 11'b00000000100;
    W_in[5][14] = 11'b11111111011;
    W_in[5][15] = 11'b00000000001;
    W_in[5][16] = 11'b00000000000;
    W_in[5][17] = 11'b00000000000;
    W_in[5][18] = 11'b00000000000;
    W_in[5][19] = 11'b11111111101;
    W_in[5][20] = 11'b00000000000;
    W_in[5][21] = 11'b00000000001;
    W_in[5][22] = 11'b11111111110;
    W_in[5][23] = 11'b11111111101;
    W_in[5][24] = 11'b00000000000;
    W_in[5][25] = 11'b00000000110;
    W_in[5][26] = 11'b11111111010;
    W_in[5][27] = 11'b11111111010;
    W_in[5][28] = 11'b00000000111;
    W_in[5][29] = 11'b00000000010;
    W_in[5][30] = 11'b00000000000;
    W_in[5][31] = 11'b00000000000;
    W_in[5][32] = 11'b11111111100;
    W_in[5][33] = 11'b00000000000;
    W_in[5][34] = 11'b11111111111;
    W_in[5][35] = 11'b00000000000;
    W_in[5][36] = 11'b00000000010;
    W_in[5][37] = 11'b00000000001;
    W_in[5][38] = 11'b00000000010;
    W_in[5][39] = 11'b00000000100;
    W_in[5][40] = 11'b00000000010;
    W_in[5][41] = 11'b00000000000;
    W_in[5][42] = 11'b00000000000;
    W_in[5][43] = 11'b00000000010;
    W_in[5][44] = 11'b00000000001;
    W_in[5][45] = 11'b00000000010;
    W_in[5][46] = 11'b00000000000;
    W_in[5][47] = 11'b11111111111;
    W_in[5][48] = 11'b11111111111;
    W_in[5][49] = 11'b11111111001;
    W_in[5][50] = 11'b00000000100;
    W_in[5][51] = 11'b00000000101;
    W_in[5][52] = 11'b11111111110;
    W_in[5][53] = 11'b11111111101;
    W_in[5][54] = 11'b11111111101;
    W_in[5][55] = 11'b11111111101;
    W_in[5][56] = 11'b11111111110;
    W_in[5][57] = 11'b00000000110;
    W_in[5][58] = 11'b00000000100;
    W_in[5][59] = 11'b11111111100;
    W_in[5][60] = 11'b11111111111;
    W_in[5][61] = 11'b11111111110;
    W_in[5][62] = 11'b00000000101;
    W_in[5][63] = 11'b11111111101;
    W_in[6][0] = 11'b11111111101;
    W_in[6][1] = 11'b11111111110;
    W_in[6][2] = 11'b11111111001;
    W_in[6][3] = 11'b11111111100;
    W_in[6][4] = 11'b11111111110;
    W_in[6][5] = 11'b11111111111;
    W_in[6][6] = 11'b00000000001;
    W_in[6][7] = 11'b11111111011;
    W_in[6][8] = 11'b11111111111;
    W_in[6][9] = 11'b11111111111;
    W_in[6][10] = 11'b11111111111;
    W_in[6][11] = 11'b11111111001;
    W_in[6][12] = 11'b11111111111;
    W_in[6][13] = 11'b00000000010;
    W_in[6][14] = 11'b11111111111;
    W_in[6][15] = 11'b00000000011;
    W_in[6][16] = 11'b11111111011;
    W_in[6][17] = 11'b00000000111;
    W_in[6][18] = 11'b00000000000;
    W_in[6][19] = 11'b00000000010;
    W_in[6][20] = 11'b00000000010;
    W_in[6][21] = 11'b11111111110;
    W_in[6][22] = 11'b00000000100;
    W_in[6][23] = 11'b00000000111;
    W_in[6][24] = 11'b00000000011;
    W_in[6][25] = 11'b00000000001;
    W_in[6][26] = 11'b00000000000;
    W_in[6][27] = 11'b11111111001;
    W_in[6][28] = 11'b11111111110;
    W_in[6][29] = 11'b00000001000;
    W_in[6][30] = 11'b11111111101;
    W_in[6][31] = 11'b11111111101;
    W_in[6][32] = 11'b00000000000;
    W_in[6][33] = 11'b00000000011;
    W_in[6][34] = 11'b11111111111;
    W_in[6][35] = 11'b11111111110;
    W_in[6][36] = 11'b00000000000;
    W_in[6][37] = 11'b00000000001;
    W_in[6][38] = 11'b00000000100;
    W_in[6][39] = 11'b00000000000;
    W_in[6][40] = 11'b00000000100;
    W_in[6][41] = 11'b11111111110;
    W_in[6][42] = 11'b00000000100;
    W_in[6][43] = 11'b00000000000;
    W_in[6][44] = 11'b00000000001;
    W_in[6][45] = 11'b00000000010;
    W_in[6][46] = 11'b00000000010;
    W_in[6][47] = 11'b00000000001;
    W_in[6][48] = 11'b00000000010;
    W_in[6][49] = 11'b00000000001;
    W_in[6][50] = 11'b11111111100;
    W_in[6][51] = 11'b00000000011;
    W_in[6][52] = 11'b00000000011;
    W_in[6][53] = 11'b00000000010;
    W_in[6][54] = 11'b11111111001;
    W_in[6][55] = 11'b00000000010;
    W_in[6][56] = 11'b00000000010;
    W_in[6][57] = 11'b11111111011;
    W_in[6][58] = 11'b11111111100;
    W_in[6][59] = 11'b11111111101;
    W_in[6][60] = 11'b00000000101;
    W_in[6][61] = 11'b00000000010;
    W_in[6][62] = 11'b00000000101;
    W_in[6][63] = 11'b00000001001;
    W_in[7][0] = 11'b00000000000;
    W_in[7][1] = 11'b00000001000;
    W_in[7][2] = 11'b00000000000;
    W_in[7][3] = 11'b00000000110;
    W_in[7][4] = 11'b11111111010;
    W_in[7][5] = 11'b00000000001;
    W_in[7][6] = 11'b00000000001;
    W_in[7][7] = 11'b11111111110;
    W_in[7][8] = 11'b11111111111;
    W_in[7][9] = 11'b00000000101;
    W_in[7][10] = 11'b11111111100;
    W_in[7][11] = 11'b11111111111;
    W_in[7][12] = 11'b11111111100;
    W_in[7][13] = 11'b11111111111;
    W_in[7][14] = 11'b11111111110;
    W_in[7][15] = 11'b11111111111;
    W_in[7][16] = 11'b00000000000;
    W_in[7][17] = 11'b00000000001;
    W_in[7][18] = 11'b11111111101;
    W_in[7][19] = 11'b00000000100;
    W_in[7][20] = 11'b11111111110;
    W_in[7][21] = 11'b00000000010;
    W_in[7][22] = 11'b00000000011;
    W_in[7][23] = 11'b00000000010;
    W_in[7][24] = 11'b00000000111;
    W_in[7][25] = 11'b00000000001;
    W_in[7][26] = 11'b11111111111;
    W_in[7][27] = 11'b11111111110;
    W_in[7][28] = 11'b00000000001;
    W_in[7][29] = 11'b00000000001;
    W_in[7][30] = 11'b11111111100;
    W_in[7][31] = 11'b00000001000;
    W_in[7][32] = 11'b00000000100;
    W_in[7][33] = 11'b11111111011;
    W_in[7][34] = 11'b00000000010;
    W_in[7][35] = 11'b00000000001;
    W_in[7][36] = 11'b00000000001;
    W_in[7][37] = 11'b11111111001;
    W_in[7][38] = 11'b00000000011;
    W_in[7][39] = 11'b00000000000;
    W_in[7][40] = 11'b00000000000;
    W_in[7][41] = 11'b00000000101;
    W_in[7][42] = 11'b11111111011;
    W_in[7][43] = 11'b00000000001;
    W_in[7][44] = 11'b11111111101;
    W_in[7][45] = 11'b11111111110;
    W_in[7][46] = 11'b00000000110;
    W_in[7][47] = 11'b11111111101;
    W_in[7][48] = 11'b11111111110;
    W_in[7][49] = 11'b11111111111;
    W_in[7][50] = 11'b11111111100;
    W_in[7][51] = 11'b11111111101;
    W_in[7][52] = 11'b11111111101;
    W_in[7][53] = 11'b11111111100;
    W_in[7][54] = 11'b11111111110;
    W_in[7][55] = 11'b11111111001;
    W_in[7][56] = 11'b11111111101;
    W_in[7][57] = 11'b00000000100;
    W_in[7][58] = 11'b11111111100;
    W_in[7][59] = 11'b11111111101;
    W_in[7][60] = 11'b11111111101;
    W_in[7][61] = 11'b11111111101;
    W_in[7][62] = 11'b11111111010;
    W_in[7][63] = 11'b11111111110;
    W_in[8][0] = 11'b00000000000;
    W_in[8][1] = 11'b11111111110;
    W_in[8][2] = 11'b11111111111;
    W_in[8][3] = 11'b11111111101;
    W_in[8][4] = 11'b00000000000;
    W_in[8][5] = 11'b00000000011;
    W_in[8][6] = 11'b11111111100;
    W_in[8][7] = 11'b11111111011;
    W_in[8][8] = 11'b11111111001;
    W_in[8][9] = 11'b11111111101;
    W_in[8][10] = 11'b11111111001;
    W_in[8][11] = 11'b11111111110;
    W_in[8][12] = 11'b11111111111;
    W_in[8][13] = 11'b00000000011;
    W_in[8][14] = 11'b00000000001;
    W_in[8][15] = 11'b11111111111;
    W_in[8][16] = 11'b11111111100;
    W_in[8][17] = 11'b11111111101;
    W_in[8][18] = 11'b11111111100;
    W_in[8][19] = 11'b11111111011;
    W_in[8][20] = 11'b11111111111;
    W_in[8][21] = 11'b00000000011;
    W_in[8][22] = 11'b00000001000;
    W_in[8][23] = 11'b00000000101;
    W_in[8][24] = 11'b11111111001;
    W_in[8][25] = 11'b11111111010;
    W_in[8][26] = 11'b00000000000;
    W_in[8][27] = 11'b11111111001;
    W_in[8][28] = 11'b00000000110;
    W_in[8][29] = 11'b00000000000;
    W_in[8][30] = 11'b00000000110;
    W_in[8][31] = 11'b11111111100;
    W_in[8][32] = 11'b11111111001;
    W_in[8][33] = 11'b11111111010;
    W_in[8][34] = 11'b11111111100;
    W_in[8][35] = 11'b11111111100;
    W_in[8][36] = 11'b11111111010;
    W_in[8][37] = 11'b11111111011;
    W_in[8][38] = 11'b11111111101;
    W_in[8][39] = 11'b00000000010;
    W_in[8][40] = 11'b00000000001;
    W_in[8][41] = 11'b11111111100;
    W_in[8][42] = 11'b11111111111;
    W_in[8][43] = 11'b11111111101;
    W_in[8][44] = 11'b11111111000;
    W_in[8][45] = 11'b11111111111;
    W_in[8][46] = 11'b11111111111;
    W_in[8][47] = 11'b11111111111;
    W_in[8][48] = 11'b00000000000;
    W_in[8][49] = 11'b11111111110;
    W_in[8][50] = 11'b00000000101;
    W_in[8][51] = 11'b11111111101;
    W_in[8][52] = 11'b00000000111;
    W_in[8][53] = 11'b00000000100;
    W_in[8][54] = 11'b00000001000;
    W_in[8][55] = 11'b00000000110;
    W_in[8][56] = 11'b00000000011;
    W_in[8][57] = 11'b11111111001;
    W_in[8][58] = 11'b00000000100;
    W_in[8][59] = 11'b00000001110;
    W_in[8][60] = 11'b00000001010;
    W_in[8][61] = 11'b00000001011;
    W_in[8][62] = 11'b00000001101;
    W_in[8][63] = 11'b00000001100;
    W_in[9][0] = 11'b00000000001;
    W_in[9][1] = 11'b00000000001;
    W_in[9][2] = 11'b00000000010;
    W_in[9][3] = 11'b11111111111;
    W_in[9][4] = 11'b11111111111;
    W_in[9][5] = 11'b11111111011;
    W_in[9][6] = 11'b00000000110;
    W_in[9][7] = 11'b11111111001;
    W_in[9][8] = 11'b11111111010;
    W_in[9][9] = 11'b11111111110;
    W_in[9][10] = 11'b00000000000;
    W_in[9][11] = 11'b11111111111;
    W_in[9][12] = 11'b11111111100;
    W_in[9][13] = 11'b11111111111;
    W_in[9][14] = 11'b11111111100;
    W_in[9][15] = 11'b11111111100;
    W_in[9][16] = 11'b00000000101;
    W_in[9][17] = 11'b11111111011;
    W_in[9][18] = 11'b00000000001;
    W_in[9][19] = 11'b11111111010;
    W_in[9][20] = 11'b11111111111;
    W_in[9][21] = 11'b00000000000;
    W_in[9][22] = 11'b00000000011;
    W_in[9][23] = 11'b00000000010;
    W_in[9][24] = 11'b11111111111;
    W_in[9][25] = 11'b11111111101;
    W_in[9][26] = 11'b11111111111;
    W_in[9][27] = 11'b00000000011;
    W_in[9][28] = 11'b00000000001;
    W_in[9][29] = 11'b11111111100;
    W_in[9][30] = 11'b11111111110;
    W_in[9][31] = 11'b11111111001;
    W_in[9][32] = 11'b00000000000;
    W_in[9][33] = 11'b11111111000;
    W_in[9][34] = 11'b11111111110;
    W_in[9][35] = 11'b00000000100;
    W_in[9][36] = 11'b11111111100;
    W_in[9][37] = 11'b11111111010;
    W_in[9][38] = 11'b11111110111;
    W_in[9][39] = 11'b00000000101;
    W_in[9][40] = 11'b11111111101;
    W_in[9][41] = 11'b11111111111;
    W_in[9][42] = 11'b00000000000;
    W_in[9][43] = 11'b11111111101;
    W_in[9][44] = 11'b00000000001;
    W_in[9][45] = 11'b11111111101;
    W_in[9][46] = 11'b11111111111;
    W_in[9][47] = 11'b00000000100;
    W_in[9][48] = 11'b00000000010;
    W_in[9][49] = 11'b00000000010;
    W_in[9][50] = 11'b00000000001;
    W_in[9][51] = 11'b00000000001;
    W_in[9][52] = 11'b11111111110;
    W_in[9][53] = 11'b11111111101;
    W_in[9][54] = 11'b00000000010;
    W_in[9][55] = 11'b00000000000;
    W_in[9][56] = 11'b00000000001;
    W_in[9][57] = 11'b11111111011;
    W_in[9][58] = 11'b11111111100;
    W_in[9][59] = 11'b11111111110;
    W_in[9][60] = 11'b00000000111;
    W_in[9][61] = 11'b00000000101;
    W_in[9][62] = 11'b11111111110;
    W_in[9][63] = 11'b00000000101;
    W_in[10][0] = 11'b00000000110;
    W_in[10][1] = 11'b11111111110;
    W_in[10][2] = 11'b00000001001;
    W_in[10][3] = 11'b11111111110;
    W_in[10][4] = 11'b00000000101;
    W_in[10][5] = 11'b00000000001;
    W_in[10][6] = 11'b11111111001;
    W_in[10][7] = 11'b00000001001;
    W_in[10][8] = 11'b00000001011;
    W_in[10][9] = 11'b00000000110;
    W_in[10][10] = 11'b00000001000;
    W_in[10][11] = 11'b00000000000;
    W_in[10][12] = 11'b00000000000;
    W_in[10][13] = 11'b00000000010;
    W_in[10][14] = 11'b11111111110;
    W_in[10][15] = 11'b11111111001;
    W_in[10][16] = 11'b11111111101;
    W_in[10][17] = 11'b00000000101;
    W_in[10][18] = 11'b00000000000;
    W_in[10][19] = 11'b00000000000;
    W_in[10][20] = 11'b11111111111;
    W_in[10][21] = 11'b11111111011;
    W_in[10][22] = 11'b00000001001;
    W_in[10][23] = 11'b00000000000;
    W_in[10][24] = 11'b11111111011;
    W_in[10][25] = 11'b00000000011;
    W_in[10][26] = 11'b11111111010;
    W_in[10][27] = 11'b11111111100;
    W_in[10][28] = 11'b00000000110;
    W_in[10][29] = 11'b00000000101;
    W_in[10][30] = 11'b11111111011;
    W_in[10][31] = 11'b00000000101;
    W_in[10][32] = 11'b00000000000;
    W_in[10][33] = 11'b00000000011;
    W_in[10][34] = 11'b00000000111;
    W_in[10][35] = 11'b00000001000;
    W_in[10][36] = 11'b11111111111;
    W_in[10][37] = 11'b00000000010;
    W_in[10][38] = 11'b11111111000;
    W_in[10][39] = 11'b11111111111;
    W_in[10][40] = 11'b00000000100;
    W_in[10][41] = 11'b11111111101;
    W_in[10][42] = 11'b00000001001;
    W_in[10][43] = 11'b00000000010;
    W_in[10][44] = 11'b00000000100;
    W_in[10][45] = 11'b11111111100;
    W_in[10][46] = 11'b11111111001;
    W_in[10][47] = 11'b00000001000;
    W_in[10][48] = 11'b11111111010;
    W_in[10][49] = 11'b11111111100;
    W_in[10][50] = 11'b00000000100;
    W_in[10][51] = 11'b11111111111;
    W_in[10][52] = 11'b00000000100;
    W_in[10][53] = 11'b11111110010;
    W_in[10][54] = 11'b11111111110;
    W_in[10][55] = 11'b00000000001;
    W_in[10][56] = 11'b11111111011;
    W_in[10][57] = 11'b11111111110;
    W_in[10][58] = 11'b11111111011;
    W_in[10][59] = 11'b11111111010;
    W_in[10][60] = 11'b11111111110;
    W_in[10][61] = 11'b11111110100;
    W_in[10][62] = 11'b11111110001;
    W_in[10][63] = 11'b11111110000;
    W_in[11][0] = 11'b11111110101;
    W_in[11][1] = 11'b11111110101;
    W_in[11][2] = 11'b00000000011;
    W_in[11][3] = 11'b11111111110;
    W_in[11][4] = 11'b00000000110;
    W_in[11][5] = 11'b00000001000;
    W_in[11][6] = 11'b11111111001;
    W_in[11][7] = 11'b00000000010;
    W_in[11][8] = 11'b11111111011;
    W_in[11][9] = 11'b11111110100;
    W_in[11][10] = 11'b11111111100;
    W_in[11][11] = 11'b00000000101;
    W_in[11][12] = 11'b00000000110;
    W_in[11][13] = 11'b11111111010;
    W_in[11][14] = 11'b00000000110;
    W_in[11][15] = 11'b00000000000;
    W_in[11][16] = 11'b00000000001;
    W_in[11][17] = 11'b11111111101;
    W_in[11][18] = 11'b00000000001;
    W_in[11][19] = 11'b00000000111;
    W_in[11][20] = 11'b11111111100;
    W_in[11][21] = 11'b11111111101;
    W_in[11][22] = 11'b00000001000;
    W_in[11][23] = 11'b11111111101;
    W_in[11][24] = 11'b00000000111;
    W_in[11][25] = 11'b00000000011;
    W_in[11][26] = 11'b00000000100;
    W_in[11][27] = 11'b11111111110;
    W_in[11][28] = 11'b00000000110;
    W_in[11][29] = 11'b00000001001;
    W_in[11][30] = 11'b00000000110;
    W_in[11][31] = 11'b00000000011;
    W_in[11][32] = 11'b11111111011;
    W_in[11][33] = 11'b11111111101;
    W_in[11][34] = 11'b11111110100;
    W_in[11][35] = 11'b11111111010;
    W_in[11][36] = 11'b00000001000;
    W_in[11][37] = 11'b00000000000;
    W_in[11][38] = 11'b00000000110;
    W_in[11][39] = 11'b11111110111;
    W_in[11][40] = 11'b00000000000;
    W_in[11][41] = 11'b11111111000;
    W_in[11][42] = 11'b11111110111;
    W_in[11][43] = 11'b11111110111;
    W_in[11][44] = 11'b11111111011;
    W_in[11][45] = 11'b00000000001;
    W_in[11][46] = 11'b00000010010;
    W_in[11][47] = 11'b11111111011;
    W_in[11][48] = 11'b11111111111;
    W_in[11][49] = 11'b11111111011;
    W_in[11][50] = 11'b11111111000;
    W_in[11][51] = 11'b00000001100;
    W_in[11][52] = 11'b11111110111;
    W_in[11][53] = 11'b00000000011;
    W_in[11][54] = 11'b00000001001;
    W_in[11][55] = 11'b00000000001;
    W_in[11][56] = 11'b00000010010;
    W_in[11][57] = 11'b00000000010;
    W_in[11][58] = 11'b00000010011;
    W_in[11][59] = 11'b00000000011;
    W_in[11][60] = 11'b11111111000;
    W_in[11][61] = 11'b00000001001;
    W_in[11][62] = 11'b00000001100;
    W_in[11][63] = 11'b11111111000;
    W_in[12][0] = 11'b11111111100;
    W_in[12][1] = 11'b00000000010;
    W_in[12][2] = 11'b11111111110;
    W_in[12][3] = 11'b00000000100;
    W_in[12][4] = 11'b11111111111;
    W_in[12][5] = 11'b11111111110;
    W_in[12][6] = 11'b11111111001;
    W_in[12][7] = 11'b11111111100;
    W_in[12][8] = 11'b11111111110;
    W_in[12][9] = 11'b00000000101;
    W_in[12][10] = 11'b00000000010;
    W_in[12][11] = 11'b00000000111;
    W_in[12][12] = 11'b11111111110;
    W_in[12][13] = 11'b00000000100;
    W_in[12][14] = 11'b00000000100;
    W_in[12][15] = 11'b00000000010;
    W_in[12][16] = 11'b11111111111;
    W_in[12][17] = 11'b00000000101;
    W_in[12][18] = 11'b00000001000;
    W_in[12][19] = 11'b00000000100;
    W_in[12][20] = 11'b11111111111;
    W_in[12][21] = 11'b00000000001;
    W_in[12][22] = 11'b00000000110;
    W_in[12][23] = 11'b00000000001;
    W_in[12][24] = 11'b00000000000;
    W_in[12][25] = 11'b11111111111;
    W_in[12][26] = 11'b11111111001;
    W_in[12][27] = 11'b00000000010;
    W_in[12][28] = 11'b00000000100;
    W_in[12][29] = 11'b00000000000;
    W_in[12][30] = 11'b00000000101;
    W_in[12][31] = 11'b00000000100;
    W_in[12][32] = 11'b11111111111;
    W_in[12][33] = 11'b11111111011;
    W_in[12][34] = 11'b11111111010;
    W_in[12][35] = 11'b11111111101;
    W_in[12][36] = 11'b11111111101;
    W_in[12][37] = 11'b11111110110;
    W_in[12][38] = 11'b00000000010;
    W_in[12][39] = 11'b11111111111;
    W_in[12][40] = 11'b11111111111;
    W_in[12][41] = 11'b00000000111;
    W_in[12][42] = 11'b11111111011;
    W_in[12][43] = 11'b00000000100;
    W_in[12][44] = 11'b00000000000;
    W_in[12][45] = 11'b11111111100;
    W_in[12][46] = 11'b11111111011;
    W_in[12][47] = 11'b00000000101;
    W_in[12][48] = 11'b00000000010;
    W_in[12][49] = 11'b00000001001;
    W_in[12][50] = 11'b00000000000;
    W_in[12][51] = 11'b00000000010;
    W_in[12][52] = 11'b11111111110;
    W_in[12][53] = 11'b11111111010;
    W_in[12][54] = 11'b11111111001;
    W_in[12][55] = 11'b11111111101;
    W_in[12][56] = 11'b00000000111;
    W_in[12][57] = 11'b11111111110;
    W_in[12][58] = 11'b00000001000;
    W_in[12][59] = 11'b11111111110;
    W_in[12][60] = 11'b11111110111;
    W_in[12][61] = 11'b11111110010;
    W_in[12][62] = 11'b11111110000;
    W_in[12][63] = 11'b00000000011;
    W_in[13][0] = 11'b00000000110;
    W_in[13][1] = 11'b00000000010;
    W_in[13][2] = 11'b00000000001;
    W_in[13][3] = 11'b00000000000;
    W_in[13][4] = 11'b00000000001;
    W_in[13][5] = 11'b00000000101;
    W_in[13][6] = 11'b11111111010;
    W_in[13][7] = 11'b11111111011;
    W_in[13][8] = 11'b00000000000;
    W_in[13][9] = 11'b00000001000;
    W_in[13][10] = 11'b00000000100;
    W_in[13][11] = 11'b11111111000;
    W_in[13][12] = 11'b11111111011;
    W_in[13][13] = 11'b00000000101;
    W_in[13][14] = 11'b11111111110;
    W_in[13][15] = 11'b00000000110;
    W_in[13][16] = 11'b11111111000;
    W_in[13][17] = 11'b00000000100;
    W_in[13][18] = 11'b00000001001;
    W_in[13][19] = 11'b11111111011;
    W_in[13][20] = 11'b11111111011;
    W_in[13][21] = 11'b11111111001;
    W_in[13][22] = 11'b00000000100;
    W_in[13][23] = 11'b00000001010;
    W_in[13][24] = 11'b00000000100;
    W_in[13][25] = 11'b11111111100;
    W_in[13][26] = 11'b11111111101;
    W_in[13][27] = 11'b11111111100;
    W_in[13][28] = 11'b11111111101;
    W_in[13][29] = 11'b11111111010;
    W_in[13][30] = 11'b11111111110;
    W_in[13][31] = 11'b11111111010;
    W_in[13][32] = 11'b00000000101;
    W_in[13][33] = 11'b11111111110;
    W_in[13][34] = 11'b11111111100;
    W_in[13][35] = 11'b00000000101;
    W_in[13][36] = 11'b11111110111;
    W_in[13][37] = 11'b00000000001;
    W_in[13][38] = 11'b00000000000;
    W_in[13][39] = 11'b11111111100;
    W_in[13][40] = 11'b00000000110;
    W_in[13][41] = 11'b00000000011;
    W_in[13][42] = 11'b00000000111;
    W_in[13][43] = 11'b00000000110;
    W_in[13][44] = 11'b00000000000;
    W_in[13][45] = 11'b00000000111;
    W_in[13][46] = 11'b00000000010;
    W_in[13][47] = 11'b11111111110;
    W_in[13][48] = 11'b11111111010;
    W_in[13][49] = 11'b11111111111;
    W_in[13][50] = 11'b11111111101;
    W_in[13][51] = 11'b00000000100;
    W_in[13][52] = 11'b00000000101;
    W_in[13][53] = 11'b00000000011;
    W_in[13][54] = 11'b11111111000;
    W_in[13][55] = 11'b00000001010;
    W_in[13][56] = 11'b00000000101;
    W_in[13][57] = 11'b11111111110;
    W_in[13][58] = 11'b11111111111;
    W_in[13][59] = 11'b00000000111;
    W_in[13][60] = 11'b11111110111;
    W_in[13][61] = 11'b00000000000;
    W_in[13][62] = 11'b11111111101;
    W_in[13][63] = 11'b11111111101;
    W_in[14][0] = 11'b00000000011;
    W_in[14][1] = 11'b00000000100;
    W_in[14][2] = 11'b11111111111;
    W_in[14][3] = 11'b00000000010;
    W_in[14][4] = 11'b00000000110;
    W_in[14][5] = 11'b00000000011;
    W_in[14][6] = 11'b11111110111;
    W_in[14][7] = 11'b00000000011;
    W_in[14][8] = 11'b11111110100;
    W_in[14][9] = 11'b11111111110;
    W_in[14][10] = 11'b00000000000;
    W_in[14][11] = 11'b11111111100;
    W_in[14][12] = 11'b11111111001;
    W_in[14][13] = 11'b00000000011;
    W_in[14][14] = 11'b00000000000;
    W_in[14][15] = 11'b11111110101;
    W_in[14][16] = 11'b00000000100;
    W_in[14][17] = 11'b00000000101;
    W_in[14][18] = 11'b11111110100;
    W_in[14][19] = 11'b11111111000;
    W_in[14][20] = 11'b00000000111;
    W_in[14][21] = 11'b11111111010;
    W_in[14][22] = 11'b00000000011;
    W_in[14][23] = 11'b11111111010;
    W_in[14][24] = 11'b00000000011;
    W_in[14][25] = 11'b11111111011;
    W_in[14][26] = 11'b00000001001;
    W_in[14][27] = 11'b11111111110;
    W_in[14][28] = 11'b00000000110;
    W_in[14][29] = 11'b00000001001;
    W_in[14][30] = 11'b11111111111;
    W_in[14][31] = 11'b00000000000;
    W_in[14][32] = 11'b00000001011;
    W_in[14][33] = 11'b11111111000;
    W_in[14][34] = 11'b11111111000;
    W_in[14][35] = 11'b11111111100;
    W_in[14][36] = 11'b00000001010;
    W_in[14][37] = 11'b00000001000;
    W_in[14][38] = 11'b11111111011;
    W_in[14][39] = 11'b11111110101;
    W_in[14][40] = 11'b00000000100;
    W_in[14][41] = 11'b11111111111;
    W_in[14][42] = 11'b11111111000;
    W_in[14][43] = 11'b00000000001;
    W_in[14][44] = 11'b11111111101;
    W_in[14][45] = 11'b00000000101;
    W_in[14][46] = 11'b11111111110;
    W_in[14][47] = 11'b11111111110;
    W_in[14][48] = 11'b11111111101;
    W_in[14][49] = 11'b00000000000;
    W_in[14][50] = 11'b11111111000;
    W_in[14][51] = 11'b11111111101;
    W_in[14][52] = 11'b11111111000;
    W_in[14][53] = 11'b00000000111;
    W_in[14][54] = 11'b11111111111;
    W_in[14][55] = 11'b11111111100;
    W_in[14][56] = 11'b11111111101;
    W_in[14][57] = 11'b00000000111;
    W_in[14][58] = 11'b00000001000;
    W_in[14][59] = 11'b00000001010;
    W_in[14][60] = 11'b00000001111;
    W_in[14][61] = 11'b00000001010;
    W_in[14][62] = 11'b00000010001;
    W_in[14][63] = 11'b00000001101;
    W_in[15][0] = 11'b11111110101;
    W_in[15][1] = 11'b00000001000;
    W_in[15][2] = 11'b00000000001;
    W_in[15][3] = 11'b00000001001;
    W_in[15][4] = 11'b11111110110;
    W_in[15][5] = 11'b00000000010;
    W_in[15][6] = 11'b11111110111;
    W_in[15][7] = 11'b00000000101;
    W_in[15][8] = 11'b11111110010;
    W_in[15][9] = 11'b11111110101;
    W_in[15][10] = 11'b00000001001;
    W_in[15][11] = 11'b11111110101;
    W_in[15][12] = 11'b11111110101;
    W_in[15][13] = 11'b00000000101;
    W_in[15][14] = 11'b00000000100;
    W_in[15][15] = 11'b00000000100;
    W_in[15][16] = 11'b00000001011;
    W_in[15][17] = 11'b11111111110;
    W_in[15][18] = 11'b00000000000;
    W_in[15][19] = 11'b00000001101;
    W_in[15][20] = 11'b11111111110;
    W_in[15][21] = 11'b11111111000;
    W_in[15][22] = 11'b11111111101;
    W_in[15][23] = 11'b11111111100;
    W_in[15][24] = 11'b11111110110;
    W_in[15][25] = 11'b11111111110;
    W_in[15][26] = 11'b11111111000;
    W_in[15][27] = 11'b11111110110;
    W_in[15][28] = 11'b00000001101;
    W_in[15][29] = 11'b00000000100;
    W_in[15][30] = 11'b00000000001;
    W_in[15][31] = 11'b00000000111;
    W_in[15][32] = 11'b00000000100;
    W_in[15][33] = 11'b11111111110;
    W_in[15][34] = 11'b00000000111;
    W_in[15][35] = 11'b00000000100;
    W_in[15][36] = 11'b11111110111;
    W_in[15][37] = 11'b11111110110;
    W_in[15][38] = 11'b00000000100;
    W_in[15][39] = 11'b00000000000;
    W_in[15][40] = 11'b11111110100;
    W_in[15][41] = 11'b11111110110;
    W_in[15][42] = 11'b00000001000;
    W_in[15][43] = 11'b00000000001;
    W_in[15][44] = 11'b00000000011;
    W_in[15][45] = 11'b00000001100;
    W_in[15][46] = 11'b11111111111;
    W_in[15][47] = 11'b00000001010;
    W_in[15][48] = 11'b00000000001;
    W_in[15][49] = 11'b11111111111;
    W_in[15][50] = 11'b11111111011;
    W_in[15][51] = 11'b00000000110;
    W_in[15][52] = 11'b11111111110;
    W_in[15][53] = 11'b11111110110;
    W_in[15][54] = 11'b00000001100;
    W_in[15][55] = 11'b00000000010;
    W_in[15][56] = 11'b11111111010;
    W_in[15][57] = 11'b00000000110;
    W_in[15][58] = 11'b11111111011;
    W_in[15][59] = 11'b00000001011;
    W_in[15][60] = 11'b00000001011;
    W_in[15][61] = 11'b00000000011;
    W_in[15][62] = 11'b00000000001;
    W_in[15][63] = 11'b00000001001;

    // Initialize W_hr weights
    W_hr[0][0] = 11'b00000000000;
    W_hr[0][1] = 11'b00000000001;
    W_hr[0][2] = 11'b00000000010;
    W_hr[0][3] = 11'b11111111011;
    W_hr[0][4] = 11'b00000001001;
    W_hr[0][5] = 11'b00000001001;
    W_hr[0][6] = 11'b00000001001;
    W_hr[0][7] = 11'b11111110111;
    W_hr[0][8] = 11'b00000001000;
    W_hr[0][9] = 11'b00000001001;
    W_hr[0][10] = 11'b11111111100;
    W_hr[0][11] = 11'b11111111011;
    W_hr[0][12] = 11'b00000000100;
    W_hr[0][13] = 11'b00000000101;
    W_hr[0][14] = 11'b00000001011;
    W_hr[0][15] = 11'b11111111000;
    W_hr[1][0] = 11'b00000000111;
    W_hr[1][1] = 11'b00000000100;
    W_hr[1][2] = 11'b11111111101;
    W_hr[1][3] = 11'b00000000100;
    W_hr[1][4] = 11'b00000001101;
    W_hr[1][5] = 11'b11111110100;
    W_hr[1][6] = 11'b00000000000;
    W_hr[1][7] = 11'b00000001001;
    W_hr[1][8] = 11'b00000000111;
    W_hr[1][9] = 11'b00000000000;
    W_hr[1][10] = 11'b11111110000;
    W_hr[1][11] = 11'b00000001110;
    W_hr[1][12] = 11'b00000001100;
    W_hr[1][13] = 11'b00000000100;
    W_hr[1][14] = 11'b11111110111;
    W_hr[1][15] = 11'b00000010101;
    W_hr[2][0] = 11'b11111111111;
    W_hr[2][1] = 11'b11111111110;
    W_hr[2][2] = 11'b00000000101;
    W_hr[2][3] = 11'b11111111010;
    W_hr[2][4] = 11'b11111111010;
    W_hr[2][5] = 11'b11111111111;
    W_hr[2][6] = 11'b00000010111;
    W_hr[2][7] = 11'b11111110100;
    W_hr[2][8] = 11'b11111111111;
    W_hr[2][9] = 11'b00000001110;
    W_hr[2][10] = 11'b00000010100;
    W_hr[2][11] = 11'b11111110010;
    W_hr[2][12] = 11'b11111111011;
    W_hr[2][13] = 11'b11111110110;
    W_hr[2][14] = 11'b11111111001;
    W_hr[2][15] = 11'b00000001010;
    W_hr[3][0] = 11'b00000000000;
    W_hr[3][1] = 11'b00000000001;
    W_hr[3][2] = 11'b00000000010;
    W_hr[3][3] = 11'b11111111011;
    W_hr[3][4] = 11'b00000001001;
    W_hr[3][5] = 11'b00000001001;
    W_hr[3][6] = 11'b00000001001;
    W_hr[3][7] = 11'b11111110111;
    W_hr[3][8] = 11'b00000001000;
    W_hr[3][9] = 11'b00000001001;
    W_hr[3][10] = 11'b11111111100;
    W_hr[3][11] = 11'b11111111011;
    W_hr[3][12] = 11'b00000000100;
    W_hr[3][13] = 11'b00000000101;
    W_hr[3][14] = 11'b00000001011;
    W_hr[3][15] = 11'b11111111000;
    W_hr[4][0] = 11'b00000000111;
    W_hr[4][1] = 11'b00000000100;
    W_hr[4][2] = 11'b11111111101;
    W_hr[4][3] = 11'b00000000100;
    W_hr[4][4] = 11'b00000001101;
    W_hr[4][5] = 11'b11111110100;
    W_hr[4][6] = 11'b00000000000;
    W_hr[4][7] = 11'b00000001001;
    W_hr[4][8] = 11'b00000000111;
    W_hr[4][9] = 11'b00000000000;
    W_hr[4][10] = 11'b11111110000;
    W_hr[4][11] = 11'b00000001110;
    W_hr[4][12] = 11'b00000001100;
    W_hr[4][13] = 11'b00000000100;
    W_hr[4][14] = 11'b11111110111;
    W_hr[4][15] = 11'b00000010101;
    W_hr[5][0] = 11'b11111111111;
    W_hr[5][1] = 11'b11111111110;
    W_hr[5][2] = 11'b00000000101;
    W_hr[5][3] = 11'b11111111010;
    W_hr[5][4] = 11'b11111111010;
    W_hr[5][5] = 11'b11111111111;
    W_hr[5][6] = 11'b00000010111;
    W_hr[5][7] = 11'b11111110100;
    W_hr[5][8] = 11'b11111111111;
    W_hr[5][9] = 11'b00000001110;
    W_hr[5][10] = 11'b00000010100;
    W_hr[5][11] = 11'b11111110010;
    W_hr[5][12] = 11'b11111111011;
    W_hr[5][13] = 11'b11111110110;
    W_hr[5][14] = 11'b11111111001;
    W_hr[5][15] = 11'b00000001010;
    W_hr[6][0] = 11'b00000000000;
    W_hr[6][1] = 11'b00000000001;
    W_hr[6][2] = 11'b00000000010;
    W_hr[6][3] = 11'b11111111011;
    W_hr[6][4] = 11'b00000001001;
    W_hr[6][5] = 11'b00000001001;
    W_hr[6][6] = 11'b00000001001;
    W_hr[6][7] = 11'b11111110111;
    W_hr[6][8] = 11'b00000001000;
    W_hr[6][9] = 11'b00000001001;
    W_hr[6][10] = 11'b11111111100;
    W_hr[6][11] = 11'b11111111011;
    W_hr[6][12] = 11'b00000000100;
    W_hr[6][13] = 11'b00000000101;
    W_hr[6][14] = 11'b00000001011;
    W_hr[6][15] = 11'b11111111000;
    W_hr[7][0] = 11'b00000000111;
    W_hr[7][1] = 11'b00000000100;
    W_hr[7][2] = 11'b11111111101;
    W_hr[7][3] = 11'b00000000100;
    W_hr[7][4] = 11'b00000001101;
    W_hr[7][5] = 11'b11111110100;
    W_hr[7][6] = 11'b00000000000;
    W_hr[7][7] = 11'b00000001001;
    W_hr[7][8] = 11'b00000000111;
    W_hr[7][9] = 11'b00000000000;
    W_hr[7][10] = 11'b11111110000;
    W_hr[7][11] = 11'b00000001110;
    W_hr[7][12] = 11'b00000001100;
    W_hr[7][13] = 11'b00000000100;
    W_hr[7][14] = 11'b11111110111;
    W_hr[7][15] = 11'b00000010101;
    W_hr[8][0] = 11'b11111111111;
    W_hr[8][1] = 11'b11111111110;
    W_hr[8][2] = 11'b00000000101;
    W_hr[8][3] = 11'b11111111010;
    W_hr[8][4] = 11'b11111111010;
    W_hr[8][5] = 11'b11111111111;
    W_hr[8][6] = 11'b00000010111;
    W_hr[8][7] = 11'b11111110100;
    W_hr[8][8] = 11'b11111111111;
    W_hr[8][9] = 11'b00000001110;
    W_hr[8][10] = 11'b00000010100;
    W_hr[8][11] = 11'b11111110010;
    W_hr[8][12] = 11'b11111111011;
    W_hr[8][13] = 11'b11111110110;
    W_hr[8][14] = 11'b11111111001;
    W_hr[8][15] = 11'b00000001010;
    W_hr[9][0] = 11'b00000000000;
    W_hr[9][1] = 11'b00000000001;
    W_hr[9][2] = 11'b00000000010;
    W_hr[9][3] = 11'b11111111011;
    W_hr[9][4] = 11'b00000001001;
    W_hr[9][5] = 11'b00000001001;
    W_hr[9][6] = 11'b00000001001;
    W_hr[9][7] = 11'b11111110111;
    W_hr[9][8] = 11'b00000001000;
    W_hr[9][9] = 11'b00000001001;
    W_hr[9][10] = 11'b11111111100;
    W_hr[9][11] = 11'b11111111011;
    W_hr[9][12] = 11'b00000000100;
    W_hr[9][13] = 11'b00000000101;
    W_hr[9][14] = 11'b00000001011;
    W_hr[9][15] = 11'b11111111000;
    W_hr[10][0] = 11'b00000000111;
    W_hr[10][1] = 11'b00000000100;
    W_hr[10][2] = 11'b11111111101;
    W_hr[10][3] = 11'b00000000100;
    W_hr[10][4] = 11'b00000001101;
    W_hr[10][5] = 11'b11111110100;
    W_hr[10][6] = 11'b00000000000;
    W_hr[10][7] = 11'b00000001001;
    W_hr[10][8] = 11'b00000000111;
    W_hr[10][9] = 11'b00000000000;
    W_hr[10][10] = 11'b11111110000;
    W_hr[10][11] = 11'b00000001110;
    W_hr[10][12] = 11'b00000001100;
    W_hr[10][13] = 11'b00000000100;
    W_hr[10][14] = 11'b11111110111;
    W_hr[10][15] = 11'b00000010101;
    W_hr[11][0] = 11'b11111111111;
    W_hr[11][1] = 11'b11111111110;
    W_hr[11][2] = 11'b00000000101;
    W_hr[11][3] = 11'b11111111010;
    W_hr[11][4] = 11'b11111111010;
    W_hr[11][5] = 11'b11111111111;
    W_hr[11][6] = 11'b00000010111;
    W_hr[11][7] = 11'b11111110100;
    W_hr[11][8] = 11'b11111111111;
    W_hr[11][9] = 11'b00000001110;
    W_hr[11][10] = 11'b00000010100;
    W_hr[11][11] = 11'b11111110010;
    W_hr[11][12] = 11'b11111111011;
    W_hr[11][13] = 11'b11111110110;
    W_hr[11][14] = 11'b11111111001;
    W_hr[11][15] = 11'b00000001010;
    W_hr[12][0] = 11'b00000000000;
    W_hr[12][1] = 11'b00000000001;
    W_hr[12][2] = 11'b00000000010;
    W_hr[12][3] = 11'b11111111011;
    W_hr[12][4] = 11'b00000001001;
    W_hr[12][5] = 11'b00000001001;
    W_hr[12][6] = 11'b00000001001;
    W_hr[12][7] = 11'b11111110111;
    W_hr[12][8] = 11'b00000001000;
    W_hr[12][9] = 11'b00000001001;
    W_hr[12][10] = 11'b11111111100;
    W_hr[12][11] = 11'b11111111011;
    W_hr[12][12] = 11'b00000000100;
    W_hr[12][13] = 11'b00000000101;
    W_hr[12][14] = 11'b00000001011;
    W_hr[12][15] = 11'b11111111000;
    W_hr[13][0] = 11'b00000000111;
    W_hr[13][1] = 11'b00000000100;
    W_hr[13][2] = 11'b11111111101;
    W_hr[13][3] = 11'b00000000100;
    W_hr[13][4] = 11'b00000001101;
    W_hr[13][5] = 11'b11111110100;
    W_hr[13][6] = 11'b00000000000;
    W_hr[13][7] = 11'b00000001001;
    W_hr[13][8] = 11'b00000000111;
    W_hr[13][9] = 11'b00000000000;
    W_hr[13][10] = 11'b11111110000;
    W_hr[13][11] = 11'b00000001110;
    W_hr[13][12] = 11'b00000001100;
    W_hr[13][13] = 11'b00000000100;
    W_hr[13][14] = 11'b11111110111;
    W_hr[13][15] = 11'b00000010101;
    W_hr[14][0] = 11'b11111111111;
    W_hr[14][1] = 11'b11111111110;
    W_hr[14][2] = 11'b00000000101;
    W_hr[14][3] = 11'b11111111010;
    W_hr[14][4] = 11'b11111111010;
    W_hr[14][5] = 11'b11111111111;
    W_hr[14][6] = 11'b00000010111;
    W_hr[14][7] = 11'b11111110100;
    W_hr[14][8] = 11'b11111111111;
    W_hr[14][9] = 11'b00000001110;
    W_hr[14][10] = 11'b00000010100;
    W_hr[14][11] = 11'b11111110010;
    W_hr[14][12] = 11'b11111111011;
    W_hr[14][13] = 11'b11111110110;
    W_hr[14][14] = 11'b11111111001;
    W_hr[14][15] = 11'b00000001010;
    W_hr[15][0] = 11'b00000000000;
    W_hr[15][1] = 11'b00000000001;
    W_hr[15][2] = 11'b00000000010;
    W_hr[15][3] = 11'b11111111011;
    W_hr[15][4] = 11'b00000001001;
    W_hr[15][5] = 11'b00000001001;
    W_hr[15][6] = 11'b00000001001;
    W_hr[15][7] = 11'b11111110111;
    W_hr[15][8] = 11'b00000001000;
    W_hr[15][9] = 11'b00000001001;
    W_hr[15][10] = 11'b11111111100;
    W_hr[15][11] = 11'b11111111011;
    W_hr[15][12] = 11'b00000000100;
    W_hr[15][13] = 11'b00000000101;
    W_hr[15][14] = 11'b00000001011;
    W_hr[15][15] = 11'b11111111000;

    // Initialize W_hz weights
    W_hz[0][0] = 11'b00000000111;
    W_hz[0][1] = 11'b00000000100;
    W_hz[0][2] = 11'b11111111101;
    W_hz[0][3] = 11'b00000000100;
    W_hz[0][4] = 11'b00000001101;
    W_hz[0][5] = 11'b11111110100;
    W_hz[0][6] = 11'b00000000000;
    W_hz[0][7] = 11'b00000001001;
    W_hz[0][8] = 11'b00000000111;
    W_hz[0][9] = 11'b00000000000;
    W_hz[0][10] = 11'b11111110000;
    W_hz[0][11] = 11'b00000001110;
    W_hz[0][12] = 11'b00000001100;
    W_hz[0][13] = 11'b00000000100;
    W_hz[0][14] = 11'b11111110111;
    W_hz[0][15] = 11'b00000010101;
    W_hz[1][0] = 11'b11111111111;
    W_hz[1][1] = 11'b11111111110;
    W_hz[1][2] = 11'b00000000101;
    W_hz[1][3] = 11'b11111111010;
    W_hz[1][4] = 11'b11111111010;
    W_hz[1][5] = 11'b11111111111;
    W_hz[1][6] = 11'b00000010111;
    W_hz[1][7] = 11'b11111110100;
    W_hz[1][8] = 11'b11111111111;
    W_hz[1][9] = 11'b00000001110;
    W_hz[1][10] = 11'b00000010100;
    W_hz[1][11] = 11'b11111110010;
    W_hz[1][12] = 11'b11111111011;
    W_hz[1][13] = 11'b11111110110;
    W_hz[1][14] = 11'b11111111001;
    W_hz[1][15] = 11'b00000001010;
    W_hz[2][0] = 11'b00000000000;
    W_hz[2][1] = 11'b00000000001;
    W_hz[2][2] = 11'b00000000010;
    W_hz[2][3] = 11'b11111111011;
    W_hz[2][4] = 11'b00000001001;
    W_hz[2][5] = 11'b00000001001;
    W_hz[2][6] = 11'b00000001001;
    W_hz[2][7] = 11'b11111110111;
    W_hz[2][8] = 11'b00000001000;
    W_hz[2][9] = 11'b00000001001;
    W_hz[2][10] = 11'b11111111100;
    W_hz[2][11] = 11'b11111111011;
    W_hz[2][12] = 11'b00000000100;
    W_hz[2][13] = 11'b00000000101;
    W_hz[2][14] = 11'b00000001011;
    W_hz[2][15] = 11'b11111111000;
    W_hz[3][0] = 11'b00000000111;
    W_hz[3][1] = 11'b00000000100;
    W_hz[3][2] = 11'b11111111101;
    W_hz[3][3] = 11'b00000000100;
    W_hz[3][4] = 11'b00000001101;
    W_hz[3][5] = 11'b11111110100;
    W_hz[3][6] = 11'b00000000000;
    W_hz[3][7] = 11'b00000001001;
    W_hz[3][8] = 11'b00000000111;
    W_hz[3][9] = 11'b00000000000;
    W_hz[3][10] = 11'b11111110000;
    W_hz[3][11] = 11'b00000001110;
    W_hz[3][12] = 11'b00000001100;
    W_hz[3][13] = 11'b00000000100;
    W_hz[3][14] = 11'b11111110111;
    W_hz[3][15] = 11'b00000010101;
    W_hz[4][0] = 11'b11111111111;
    W_hz[4][1] = 11'b11111111110;
    W_hz[4][2] = 11'b00000000101;
    W_hz[4][3] = 11'b11111111010;
    W_hz[4][4] = 11'b11111111010;
    W_hz[4][5] = 11'b11111111111;
    W_hz[4][6] = 11'b00000010111;
    W_hz[4][7] = 11'b11111110100;
    W_hz[4][8] = 11'b11111111111;
    W_hz[4][9] = 11'b00000001110;
    W_hz[4][10] = 11'b00000010100;
    W_hz[4][11] = 11'b11111110010;
    W_hz[4][12] = 11'b11111111011;
    W_hz[4][13] = 11'b11111110110;
    W_hz[4][14] = 11'b11111111001;
    W_hz[4][15] = 11'b00000001010;
    W_hz[5][0] = 11'b00000000000;
    W_hz[5][1] = 11'b00000000001;
    W_hz[5][2] = 11'b00000000010;
    W_hz[5][3] = 11'b11111111011;
    W_hz[5][4] = 11'b00000001001;
    W_hz[5][5] = 11'b00000001001;
    W_hz[5][6] = 11'b00000001001;
    W_hz[5][7] = 11'b11111110111;
    W_hz[5][8] = 11'b00000001000;
    W_hz[5][9] = 11'b00000001001;
    W_hz[5][10] = 11'b11111111100;
    W_hz[5][11] = 11'b11111111011;
    W_hz[5][12] = 11'b00000000100;
    W_hz[5][13] = 11'b00000000101;
    W_hz[5][14] = 11'b00000001011;
    W_hz[5][15] = 11'b11111111000;
    W_hz[6][0] = 11'b00000000111;
    W_hz[6][1] = 11'b00000000100;
    W_hz[6][2] = 11'b11111111101;
    W_hz[6][3] = 11'b00000000100;
    W_hz[6][4] = 11'b00000001101;
    W_hz[6][5] = 11'b11111110100;
    W_hz[6][6] = 11'b00000000000;
    W_hz[6][7] = 11'b00000001001;
    W_hz[6][8] = 11'b00000000111;
    W_hz[6][9] = 11'b00000000000;
    W_hz[6][10] = 11'b11111110000;
    W_hz[6][11] = 11'b00000001110;
    W_hz[6][12] = 11'b00000001100;
    W_hz[6][13] = 11'b00000000100;
    W_hz[6][14] = 11'b11111110111;
    W_hz[6][15] = 11'b00000010101;
    W_hz[7][0] = 11'b11111111111;
    W_hz[7][1] = 11'b11111111110;
    W_hz[7][2] = 11'b00000000101;
    W_hz[7][3] = 11'b11111111010;
    W_hz[7][4] = 11'b11111111010;
    W_hz[7][5] = 11'b11111111111;
    W_hz[7][6] = 11'b00000010111;
    W_hz[7][7] = 11'b11111110100;
    W_hz[7][8] = 11'b11111111111;
    W_hz[7][9] = 11'b00000001110;
    W_hz[7][10] = 11'b00000010100;
    W_hz[7][11] = 11'b11111110010;
    W_hz[7][12] = 11'b11111111011;
    W_hz[7][13] = 11'b11111110110;
    W_hz[7][14] = 11'b11111111001;
    W_hz[7][15] = 11'b00000001010;
    W_hz[8][0] = 11'b00000000000;
    W_hz[8][1] = 11'b00000000001;
    W_hz[8][2] = 11'b00000000010;
    W_hz[8][3] = 11'b11111111011;
    W_hz[8][4] = 11'b00000001001;
    W_hz[8][5] = 11'b00000001001;
    W_hz[8][6] = 11'b00000001001;
    W_hz[8][7] = 11'b11111110111;
    W_hz[8][8] = 11'b00000001000;
    W_hz[8][9] = 11'b00000001001;
    W_hz[8][10] = 11'b11111111100;
    W_hz[8][11] = 11'b11111111011;
    W_hz[8][12] = 11'b00000000100;
    W_hz[8][13] = 11'b00000000101;
    W_hz[8][14] = 11'b00000001011;
    W_hz[8][15] = 11'b11111111000;
    W_hz[9][0] = 11'b00000000111;
    W_hz[9][1] = 11'b00000000100;
    W_hz[9][2] = 11'b11111111101;
    W_hz[9][3] = 11'b00000000100;
    W_hz[9][4] = 11'b00000001101;
    W_hz[9][5] = 11'b11111110100;
    W_hz[9][6] = 11'b00000000000;
    W_hz[9][7] = 11'b00000001001;
    W_hz[9][8] = 11'b00000000111;
    W_hz[9][9] = 11'b00000000000;
    W_hz[9][10] = 11'b11111110000;
    W_hz[9][11] = 11'b00000001110;
    W_hz[9][12] = 11'b00000001100;
    W_hz[9][13] = 11'b00000000100;
    W_hz[9][14] = 11'b11111110111;
    W_hz[9][15] = 11'b00000010101;
    W_hz[10][0] = 11'b11111111111;
    W_hz[10][1] = 11'b11111111110;
    W_hz[10][2] = 11'b00000000101;
    W_hz[10][3] = 11'b11111111010;
    W_hz[10][4] = 11'b11111111010;
    W_hz[10][5] = 11'b11111111111;
    W_hz[10][6] = 11'b00000010111;
    W_hz[10][7] = 11'b11111110100;
    W_hz[10][8] = 11'b11111111111;
    W_hz[10][9] = 11'b00000001110;
    W_hz[10][10] = 11'b00000010100;
    W_hz[10][11] = 11'b11111110010;
    W_hz[10][12] = 11'b11111111011;
    W_hz[10][13] = 11'b11111110110;
    W_hz[10][14] = 11'b11111111001;
    W_hz[10][15] = 11'b00000001010;
    W_hz[11][0] = 11'b00000000000;
    W_hz[11][1] = 11'b00000000001;
    W_hz[11][2] = 11'b00000000010;
    W_hz[11][3] = 11'b11111111011;
    W_hz[11][4] = 11'b00000001001;
    W_hz[11][5] = 11'b00000001001;
    W_hz[11][6] = 11'b00000001001;
    W_hz[11][7] = 11'b11111110111;
    W_hz[11][8] = 11'b00000001000;
    W_hz[11][9] = 11'b00000001001;
    W_hz[11][10] = 11'b11111111100;
    W_hz[11][11] = 11'b11111111011;
    W_hz[11][12] = 11'b00000000100;
    W_hz[11][13] = 11'b00000000101;
    W_hz[11][14] = 11'b00000001011;
    W_hz[11][15] = 11'b11111111000;
    W_hz[12][0] = 11'b00000000111;
    W_hz[12][1] = 11'b00000000100;
    W_hz[12][2] = 11'b11111111101;
    W_hz[12][3] = 11'b00000000100;
    W_hz[12][4] = 11'b00000001101;
    W_hz[12][5] = 11'b11111110100;
    W_hz[12][6] = 11'b00000000000;
    W_hz[12][7] = 11'b00000001001;
    W_hz[12][8] = 11'b00000000111;
    W_hz[12][9] = 11'b00000000000;
    W_hz[12][10] = 11'b11111110000;
    W_hz[12][11] = 11'b00000001110;
    W_hz[12][12] = 11'b00000001100;
    W_hz[12][13] = 11'b00000000100;
    W_hz[12][14] = 11'b11111110111;
    W_hz[12][15] = 11'b00000010101;
    W_hz[13][0] = 11'b11111111111;
    W_hz[13][1] = 11'b11111111110;
    W_hz[13][2] = 11'b00000000101;
    W_hz[13][3] = 11'b11111111010;
    W_hz[13][4] = 11'b11111111010;
    W_hz[13][5] = 11'b11111111111;
    W_hz[13][6] = 11'b00000010111;
    W_hz[13][7] = 11'b11111110100;
    W_hz[13][8] = 11'b11111111111;
    W_hz[13][9] = 11'b00000001110;
    W_hz[13][10] = 11'b00000010100;
    W_hz[13][11] = 11'b11111110010;
    W_hz[13][12] = 11'b11111111011;
    W_hz[13][13] = 11'b11111110110;
    W_hz[13][14] = 11'b11111111001;
    W_hz[13][15] = 11'b00000001010;
    W_hz[14][0] = 11'b00000000000;
    W_hz[14][1] = 11'b00000000001;
    W_hz[14][2] = 11'b00000000010;
    W_hz[14][3] = 11'b11111111011;
    W_hz[14][4] = 11'b00000001001;
    W_hz[14][5] = 11'b00000001001;
    W_hz[14][6] = 11'b00000001001;
    W_hz[14][7] = 11'b11111110111;
    W_hz[14][8] = 11'b00000001000;
    W_hz[14][9] = 11'b00000001001;
    W_hz[14][10] = 11'b11111111100;
    W_hz[14][11] = 11'b11111111011;
    W_hz[14][12] = 11'b00000000100;
    W_hz[14][13] = 11'b00000000101;
    W_hz[14][14] = 11'b00000001011;
    W_hz[14][15] = 11'b11111111000;
    W_hz[15][0] = 11'b00000000111;
    W_hz[15][1] = 11'b00000000100;
    W_hz[15][2] = 11'b11111111101;
    W_hz[15][3] = 11'b00000000100;
    W_hz[15][4] = 11'b00000001101;
    W_hz[15][5] = 11'b11111110100;
    W_hz[15][6] = 11'b00000000000;
    W_hz[15][7] = 11'b00000001001;
    W_hz[15][8] = 11'b00000000111;
    W_hz[15][9] = 11'b00000000000;
    W_hz[15][10] = 11'b11111110000;
    W_hz[15][11] = 11'b00000001110;
    W_hz[15][12] = 11'b00000001100;
    W_hz[15][13] = 11'b00000000100;
    W_hz[15][14] = 11'b11111110111;
    W_hz[15][15] = 11'b00000010101;

    // Initialize W_hn weights
    W_hn[0][0] = 11'b11111111111;
    W_hn[0][1] = 11'b11111111110;
    W_hn[0][2] = 11'b00000000101;
    W_hn[0][3] = 11'b11111111010;
    W_hn[0][4] = 11'b11111111010;
    W_hn[0][5] = 11'b11111111111;
    W_hn[0][6] = 11'b00000010111;
    W_hn[0][7] = 11'b11111110100;
    W_hn[0][8] = 11'b11111111111;
    W_hn[0][9] = 11'b00000001110;
    W_hn[0][10] = 11'b00000010100;
    W_hn[0][11] = 11'b11111110010;
    W_hn[0][12] = 11'b11111111011;
    W_hn[0][13] = 11'b11111110110;
    W_hn[0][14] = 11'b11111111001;
    W_hn[0][15] = 11'b00000001010;
    W_hn[1][0] = 11'b00000000000;
    W_hn[1][1] = 11'b00000000001;
    W_hn[1][2] = 11'b00000000010;
    W_hn[1][3] = 11'b11111111011;
    W_hn[1][4] = 11'b00000001001;
    W_hn[1][5] = 11'b00000001001;
    W_hn[1][6] = 11'b00000001001;
    W_hn[1][7] = 11'b11111110111;
    W_hn[1][8] = 11'b00000001000;
    W_hn[1][9] = 11'b00000001001;
    W_hn[1][10] = 11'b11111111100;
    W_hn[1][11] = 11'b11111111011;
    W_hn[1][12] = 11'b00000000100;
    W_hn[1][13] = 11'b00000000101;
    W_hn[1][14] = 11'b00000001011;
    W_hn[1][15] = 11'b11111111000;
    W_hn[2][0] = 11'b00000000111;
    W_hn[2][1] = 11'b00000000100;
    W_hn[2][2] = 11'b11111111101;
    W_hn[2][3] = 11'b00000000100;
    W_hn[2][4] = 11'b00000001101;
    W_hn[2][5] = 11'b11111110100;
    W_hn[2][6] = 11'b00000000000;
    W_hn[2][7] = 11'b00000001001;
    W_hn[2][8] = 11'b00000000111;
    W_hn[2][9] = 11'b00000000000;
    W_hn[2][10] = 11'b11111110000;
    W_hn[2][11] = 11'b00000001110;
    W_hn[2][12] = 11'b00000001100;
    W_hn[2][13] = 11'b00000000100;
    W_hn[2][14] = 11'b11111110111;
    W_hn[2][15] = 11'b00000010101;
    W_hn[3][0] = 11'b11111111111;
    W_hn[3][1] = 11'b11111111110;
    W_hn[3][2] = 11'b00000000101;
    W_hn[3][3] = 11'b11111111010;
    W_hn[3][4] = 11'b11111111010;
    W_hn[3][5] = 11'b11111111111;
    W_hn[3][6] = 11'b00000010111;
    W_hn[3][7] = 11'b11111110100;
    W_hn[3][8] = 11'b11111111111;
    W_hn[3][9] = 11'b00000001110;
    W_hn[3][10] = 11'b00000010100;
    W_hn[3][11] = 11'b11111110010;
    W_hn[3][12] = 11'b11111111011;
    W_hn[3][13] = 11'b11111110110;
    W_hn[3][14] = 11'b11111111001;
    W_hn[3][15] = 11'b00000001010;
    W_hn[4][0] = 11'b00000000000;
    W_hn[4][1] = 11'b00000000001;
    W_hn[4][2] = 11'b00000000010;
    W_hn[4][3] = 11'b11111111011;
    W_hn[4][4] = 11'b00000001001;
    W_hn[4][5] = 11'b00000001001;
    W_hn[4][6] = 11'b00000001001;
    W_hn[4][7] = 11'b11111110111;
    W_hn[4][8] = 11'b00000001000;
    W_hn[4][9] = 11'b00000001001;
    W_hn[4][10] = 11'b11111111100;
    W_hn[4][11] = 11'b11111111011;
    W_hn[4][12] = 11'b00000000100;
    W_hn[4][13] = 11'b00000000101;
    W_hn[4][14] = 11'b00000001011;
    W_hn[4][15] = 11'b11111111000;
    W_hn[5][0] = 11'b00000000111;
    W_hn[5][1] = 11'b00000000100;
    W_hn[5][2] = 11'b11111111101;
    W_hn[5][3] = 11'b00000000100;
    W_hn[5][4] = 11'b00000001101;
    W_hn[5][5] = 11'b11111110100;
    W_hn[5][6] = 11'b00000000000;
    W_hn[5][7] = 11'b00000001001;
    W_hn[5][8] = 11'b00000000111;
    W_hn[5][9] = 11'b00000000000;
    W_hn[5][10] = 11'b11111110000;
    W_hn[5][11] = 11'b00000001110;
    W_hn[5][12] = 11'b00000001100;
    W_hn[5][13] = 11'b00000000100;
    W_hn[5][14] = 11'b11111110111;
    W_hn[5][15] = 11'b00000010101;
    W_hn[6][0] = 11'b11111111111;
    W_hn[6][1] = 11'b11111111110;
    W_hn[6][2] = 11'b00000000101;
    W_hn[6][3] = 11'b11111111010;
    W_hn[6][4] = 11'b11111111010;
    W_hn[6][5] = 11'b11111111111;
    W_hn[6][6] = 11'b00000010111;
    W_hn[6][7] = 11'b11111110100;
    W_hn[6][8] = 11'b11111111111;
    W_hn[6][9] = 11'b00000001110;
    W_hn[6][10] = 11'b00000010100;
    W_hn[6][11] = 11'b11111110010;
    W_hn[6][12] = 11'b11111111011;
    W_hn[6][13] = 11'b11111110110;
    W_hn[6][14] = 11'b11111111001;
    W_hn[6][15] = 11'b00000001010;
    W_hn[7][0] = 11'b00000000000;
    W_hn[7][1] = 11'b00000000001;
    W_hn[7][2] = 11'b00000000010;
    W_hn[7][3] = 11'b11111111011;
    W_hn[7][4] = 11'b00000001001;
    W_hn[7][5] = 11'b00000001001;
    W_hn[7][6] = 11'b00000001001;
    W_hn[7][7] = 11'b11111110111;
    W_hn[7][8] = 11'b00000001000;
    W_hn[7][9] = 11'b00000001001;
    W_hn[7][10] = 11'b11111111100;
    W_hn[7][11] = 11'b11111111011;
    W_hn[7][12] = 11'b00000000100;
    W_hn[7][13] = 11'b00000000101;
    W_hn[7][14] = 11'b00000001011;
    W_hn[7][15] = 11'b11111111000;
    W_hn[8][0] = 11'b00000000111;
    W_hn[8][1] = 11'b00000000100;
    W_hn[8][2] = 11'b11111111101;
    W_hn[8][3] = 11'b00000000100;
    W_hn[8][4] = 11'b00000001101;
    W_hn[8][5] = 11'b11111110100;
    W_hn[8][6] = 11'b00000000000;
    W_hn[8][7] = 11'b00000001001;
    W_hn[8][8] = 11'b00000000111;
    W_hn[8][9] = 11'b00000000000;
    W_hn[8][10] = 11'b11111110000;
    W_hn[8][11] = 11'b00000001110;
    W_hn[8][12] = 11'b00000001100;
    W_hn[8][13] = 11'b00000000100;
    W_hn[8][14] = 11'b11111110111;
    W_hn[8][15] = 11'b00000010101;
    W_hn[9][0] = 11'b11111111111;
    W_hn[9][1] = 11'b11111111110;
    W_hn[9][2] = 11'b00000000101;
    W_hn[9][3] = 11'b11111111010;
    W_hn[9][4] = 11'b11111111010;
    W_hn[9][5] = 11'b11111111111;
    W_hn[9][6] = 11'b00000010111;
    W_hn[9][7] = 11'b11111110100;
    W_hn[9][8] = 11'b11111111111;
    W_hn[9][9] = 11'b00000001110;
    W_hn[9][10] = 11'b00000010100;
    W_hn[9][11] = 11'b11111110010;
    W_hn[9][12] = 11'b11111111011;
    W_hn[9][13] = 11'b11111110110;
    W_hn[9][14] = 11'b11111111001;
    W_hn[9][15] = 11'b00000001010;
    W_hn[10][0] = 11'b00000000000;
    W_hn[10][1] = 11'b00000000001;
    W_hn[10][2] = 11'b00000000010;
    W_hn[10][3] = 11'b11111111011;
    W_hn[10][4] = 11'b00000001001;
    W_hn[10][5] = 11'b00000001001;
    W_hn[10][6] = 11'b00000001001;
    W_hn[10][7] = 11'b11111110111;
    W_hn[10][8] = 11'b00000001000;
    W_hn[10][9] = 11'b00000001001;
    W_hn[10][10] = 11'b11111111100;
    W_hn[10][11] = 11'b11111111011;
    W_hn[10][12] = 11'b00000000100;
    W_hn[10][13] = 11'b00000000101;
    W_hn[10][14] = 11'b00000001011;
    W_hn[10][15] = 11'b11111111000;
    W_hn[11][0] = 11'b00000000111;
    W_hn[11][1] = 11'b00000000100;
    W_hn[11][2] = 11'b11111111101;
    W_hn[11][3] = 11'b00000000100;
    W_hn[11][4] = 11'b00000001101;
    W_hn[11][5] = 11'b11111110100;
    W_hn[11][6] = 11'b00000000000;
    W_hn[11][7] = 11'b00000001001;
    W_hn[11][8] = 11'b00000000111;
    W_hn[11][9] = 11'b00000000000;
    W_hn[11][10] = 11'b11111110000;
    W_hn[11][11] = 11'b00000001110;
    W_hn[11][12] = 11'b00000001100;
    W_hn[11][13] = 11'b00000000100;
    W_hn[11][14] = 11'b11111110111;
    W_hn[11][15] = 11'b00000010101;
    W_hn[12][0] = 11'b11111111111;
    W_hn[12][1] = 11'b11111111110;
    W_hn[12][2] = 11'b00000000101;
    W_hn[12][3] = 11'b11111111010;
    W_hn[12][4] = 11'b11111111010;
    W_hn[12][5] = 11'b11111111111;
    W_hn[12][6] = 11'b00000010111;
    W_hn[12][7] = 11'b11111110100;
    W_hn[12][8] = 11'b11111111111;
    W_hn[12][9] = 11'b00000001110;
    W_hn[12][10] = 11'b00000010100;
    W_hn[12][11] = 11'b11111110010;
    W_hn[12][12] = 11'b11111111011;
    W_hn[12][13] = 11'b11111110110;
    W_hn[12][14] = 11'b11111111001;
    W_hn[12][15] = 11'b00000001010;
    W_hn[13][0] = 11'b00000000000;
    W_hn[13][1] = 11'b00000000001;
    W_hn[13][2] = 11'b00000000010;
    W_hn[13][3] = 11'b11111111011;
    W_hn[13][4] = 11'b00000001001;
    W_hn[13][5] = 11'b00000001001;
    W_hn[13][6] = 11'b00000001001;
    W_hn[13][7] = 11'b11111110111;
    W_hn[13][8] = 11'b00000001000;
    W_hn[13][9] = 11'b00000001001;
    W_hn[13][10] = 11'b11111111100;
    W_hn[13][11] = 11'b11111111011;
    W_hn[13][12] = 11'b00000000100;
    W_hn[13][13] = 11'b00000000101;
    W_hn[13][14] = 11'b00000001011;
    W_hn[13][15] = 11'b11111111000;
    W_hn[14][0] = 11'b00000000111;
    W_hn[14][1] = 11'b00000000100;
    W_hn[14][2] = 11'b11111111101;
    W_hn[14][3] = 11'b00000000100;
    W_hn[14][4] = 11'b00000001101;
    W_hn[14][5] = 11'b11111110100;
    W_hn[14][6] = 11'b00000000000;
    W_hn[14][7] = 11'b00000001001;
    W_hn[14][8] = 11'b00000000111;
    W_hn[14][9] = 11'b00000000000;
    W_hn[14][10] = 11'b11111110000;
    W_hn[14][11] = 11'b00000001110;
    W_hn[14][12] = 11'b00000001100;
    W_hn[14][13] = 11'b00000000100;
    W_hn[14][14] = 11'b11111110111;
    W_hn[14][15] = 11'b00000010101;
    W_hn[15][0] = 11'b11111111111;
    W_hn[15][1] = 11'b11111111110;
    W_hn[15][2] = 11'b00000000101;
    W_hn[15][3] = 11'b11111111010;
    W_hn[15][4] = 11'b11111111010;
    W_hn[15][5] = 11'b11111111111;
    W_hn[15][6] = 11'b00000010111;
    W_hn[15][7] = 11'b11111110100;
    W_hn[15][8] = 11'b11111111111;
    W_hn[15][9] = 11'b00000001110;
    W_hn[15][10] = 11'b00000010100;
    W_hn[15][11] = 11'b11111110010;
    W_hn[15][12] = 11'b11111111011;
    W_hn[15][13] = 11'b11111110110;
    W_hn[15][14] = 11'b11111111001;
    W_hn[15][15] = 11'b00000001010;

    // Initialize biases

    // Initialize b_ir biases
    b_ir[0] = 11'b00000000001;
    b_ir[1] = 11'b00000001000;
    b_ir[2] = 11'b00000001111;
    b_ir[3] = 11'b00000000101;
    b_ir[4] = 11'b00000000110;
    b_ir[5] = 11'b00000000100;
    b_ir[6] = 11'b00000010000;
    b_ir[7] = 11'b00000000000;
    b_ir[8] = 11'b00000001011;
    b_ir[9] = 11'b00000000010;
    b_ir[10] = 11'b00000001110;
    b_ir[11] = 11'b00000000010;
    b_ir[12] = 11'b00000000010;
    b_ir[13] = 11'b00000001010;
    b_ir[14] = 11'b00000000111;
    b_ir[15] = 11'b00000001101;

    // Initialize b_iz biases
    b_iz[0] = 11'b00000000111;
    b_iz[1] = 11'b00000001001;
    b_iz[2] = 11'b00000000101;
    b_iz[3] = 11'b00000011010;
    b_iz[4] = 11'b00000000011;
    b_iz[5] = 11'b00000010011;
    b_iz[6] = 11'b00000000111;
    b_iz[7] = 11'b11111110001;
    b_iz[8] = 11'b00000000001;
    b_iz[9] = 11'b00000001000;
    b_iz[10] = 11'b00000001111;
    b_iz[11] = 11'b00000000101;
    b_iz[12] = 11'b00000000110;
    b_iz[13] = 11'b00000000100;
    b_iz[14] = 11'b00000010000;
    b_iz[15] = 11'b00000000000;

    // Initialize b_in biases
    b_in[0] = 11'b00000001011;
    b_in[1] = 11'b00000000010;
    b_in[2] = 11'b00000001110;
    b_in[3] = 11'b00000000010;
    b_in[4] = 11'b00000000010;
    b_in[5] = 11'b00000001010;
    b_in[6] = 11'b00000000111;
    b_in[7] = 11'b00000001101;
    b_in[8] = 11'b00000000111;
    b_in[9] = 11'b00000001001;
    b_in[10] = 11'b00000000101;
    b_in[11] = 11'b00000011010;
    b_in[12] = 11'b00000000011;
    b_in[13] = 11'b00000010011;
    b_in[14] = 11'b00000000111;
    b_in[15] = 11'b11111110001;

    // Initialize b_hr biases
    b_hr[0] = 11'b00000000001;
    b_hr[1] = 11'b00000001000;
    b_hr[2] = 11'b00000001111;
    b_hr[3] = 11'b00000000101;
    b_hr[4] = 11'b00000000110;
    b_hr[5] = 11'b00000000100;
    b_hr[6] = 11'b00000010000;
    b_hr[7] = 11'b00000000000;
    b_hr[8] = 11'b00000001011;
    b_hr[9] = 11'b00000000010;
    b_hr[10] = 11'b00000001110;
    b_hr[11] = 11'b00000000010;
    b_hr[12] = 11'b00000000010;
    b_hr[13] = 11'b00000001010;
    b_hr[14] = 11'b00000000111;
    b_hr[15] = 11'b00000001101;

    // Initialize b_hz biases
    b_hz[0] = 11'b00000000111;
    b_hz[1] = 11'b00000001001;
    b_hz[2] = 11'b00000000101;
    b_hz[3] = 11'b00000011010;
    b_hz[4] = 11'b00000000011;
    b_hz[5] = 11'b00000010011;
    b_hz[6] = 11'b00000000111;
    b_hz[7] = 11'b11111110001;
    b_hz[8] = 11'b00000000001;
    b_hz[9] = 11'b00000001000;
    b_hz[10] = 11'b00000001111;
    b_hz[11] = 11'b00000000101;
    b_hz[12] = 11'b00000000110;
    b_hz[13] = 11'b00000000100;
    b_hz[14] = 11'b00000010000;
    b_hz[15] = 11'b00000000000;

    // Initialize b_hn biases
    b_hn[0] = 11'b00000001011;
    b_hn[1] = 11'b00000000010;
    b_hn[2] = 11'b00000001110;
    b_hn[3] = 11'b00000000010;
    b_hn[4] = 11'b00000000010;
    b_hn[5] = 11'b00000001010;
    b_hn[6] = 11'b00000000111;
    b_hn[7] = 11'b00000001101;
    b_hn[8] = 11'b00000000111;
    b_hn[9] = 11'b00000001001;
    b_hn[10] = 11'b00000000101;
    b_hn[11] = 11'b00000011010;
    b_hn[12] = 11'b00000000011;
    b_hn[13] = 11'b00000010011;
    b_hn[14] = 11'b00000000111;
    b_hn[15] = 11'b11111110001;

    // Reset sequence
    rst_n = 0;
    start = 0;
    test_start_cycle = 0;
    test_cycles = 0;
    total_cycles = 0;
    test_timeout = 0;
    repeat(10) @(posedge clk);
    rst_n = 1;
    repeat(5) @(posedge clk);

    // Test Vector 1
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000100100;
        x_t[1] = 11'b00000110111;
        x_t[2] = 11'b00001000001;
        x_t[3] = 11'b00001001001;
        x_t[4] = 11'b00000111011;
        x_t[5] = 11'b00000110110;
        x_t[6] = 11'b00000100111;
        x_t[7] = 11'b00000100101;
        x_t[8] = 11'b00000111100;
        x_t[9] = 11'b00001001000;
        x_t[10] = 11'b00001001011;
        x_t[11] = 11'b00001001001;
        x_t[12] = 11'b00001000111;
        x_t[13] = 11'b00000101101;
        x_t[14] = 11'b00000111011;
        x_t[15] = 11'b00001000110;
        x_t[16] = 11'b00001001010;
        x_t[17] = 11'b00001001101;
        x_t[18] = 11'b00001001111;
        x_t[19] = 11'b00001001110;
        x_t[20] = 11'b00000110111;
        x_t[21] = 11'b00000010001;
        x_t[22] = 11'b00000010100;
        x_t[23] = 11'b00000010111;
        x_t[24] = 11'b00000001100;
        x_t[25] = 11'b00000001110;
        x_t[26] = 11'b00000101001;
        x_t[27] = 11'b00000011100;
        x_t[28] = 11'b00000011110;
        x_t[29] = 11'b00000001100;
        x_t[30] = 11'b00000011000;
        x_t[31] = 11'b00000110010;
        x_t[32] = 11'b00000111110;
        x_t[33] = 11'b00000111110;
        x_t[34] = 11'b00000111000;
        x_t[35] = 11'b00000101111;
        x_t[36] = 11'b00000101000;
        x_t[37] = 11'b00000010100;
        x_t[38] = 11'b00000010111;
        x_t[39] = 11'b00000100100;
        x_t[40] = 11'b00000101010;
        x_t[41] = 11'b00000110100;
        x_t[42] = 11'b00000100000;
        x_t[43] = 11'b00000011011;
        x_t[44] = 11'b00000110001;
        x_t[45] = 11'b00000010111;
        x_t[46] = 11'b00000111011;
        x_t[47] = 11'b00001000011;
        x_t[48] = 11'b00000111111;
        x_t[49] = 11'b00001000110;
        x_t[50] = 11'b00001010001;
        x_t[51] = 11'b00001010101;
        x_t[52] = 11'b00001010001;
        x_t[53] = 11'b00001000110;
        x_t[54] = 11'b00000110111;
        x_t[55] = 11'b00000110111;
        x_t[56] = 11'b00001000011;
        x_t[57] = 11'b00001000110;
        x_t[58] = 11'b00001001001;
        x_t[59] = 11'b00000101111;
        x_t[60] = 11'b00000110000;
        x_t[61] = 11'b00000110011;
        x_t[62] = 11'b00000100101;
        x_t[63] = 11'b00000110000;
        
        h_t_prev[0] = 11'b00000100100;
        h_t_prev[1] = 11'b00000110111;
        h_t_prev[2] = 11'b00001000001;
        h_t_prev[3] = 11'b00001001001;
        h_t_prev[4] = 11'b00000111011;
        h_t_prev[5] = 11'b00000110110;
        h_t_prev[6] = 11'b00000100111;
        h_t_prev[7] = 11'b00000100101;
        h_t_prev[8] = 11'b00000111100;
        h_t_prev[9] = 11'b00001001000;
        h_t_prev[10] = 11'b00001001011;
        h_t_prev[11] = 11'b00001001001;
        h_t_prev[12] = 11'b00001000111;
        h_t_prev[13] = 11'b00000101101;
        h_t_prev[14] = 11'b00000111011;
        h_t_prev[15] = 11'b00001000110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 1 timeout!");
                $fdisplay(fd_cycles, "Test Vector   1: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   1: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 1");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 2
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000101110;
        x_t[1] = 11'b00001001001;
        x_t[2] = 11'b00001010010;
        x_t[3] = 11'b00001010101;
        x_t[4] = 11'b00001001111;
        x_t[5] = 11'b00001001100;
        x_t[6] = 11'b00000111111;
        x_t[7] = 11'b00000110111;
        x_t[8] = 11'b00001010001;
        x_t[9] = 11'b00001011010;
        x_t[10] = 11'b00001011011;
        x_t[11] = 11'b00001011111;
        x_t[12] = 11'b00001011010;
        x_t[13] = 11'b00001000000;
        x_t[14] = 11'b00001001101;
        x_t[15] = 11'b00001010111;
        x_t[16] = 11'b00001011000;
        x_t[17] = 11'b00001011101;
        x_t[18] = 11'b00001011110;
        x_t[19] = 11'b00001011101;
        x_t[20] = 11'b00001000011;
        x_t[21] = 11'b00000010011;
        x_t[22] = 11'b00000010100;
        x_t[23] = 11'b00000010110;
        x_t[24] = 11'b00000011000;
        x_t[25] = 11'b00000011010;
        x_t[26] = 11'b00000101101;
        x_t[27] = 11'b00000100001;
        x_t[28] = 11'b00000011010;
        x_t[29] = 11'b00000100011;
        x_t[30] = 11'b00000101010;
        x_t[31] = 11'b00000111000;
        x_t[32] = 11'b00001000010;
        x_t[33] = 11'b00001000000;
        x_t[34] = 11'b00000111010;
        x_t[35] = 11'b00000110101;
        x_t[36] = 11'b00000101001;
        x_t[37] = 11'b00000011001;
        x_t[38] = 11'b00000110101;
        x_t[39] = 11'b00000010110;
        x_t[40] = 11'b00001000010;
        x_t[41] = 11'b11111111101;
        x_t[42] = 11'b00000111010;
        x_t[43] = 11'b00000100101;
        x_t[44] = 11'b00001001000;
        x_t[45] = 11'b00000000101;
        x_t[46] = 11'b00001001001;
        x_t[47] = 11'b00001001001;
        x_t[48] = 11'b00001000000;
        x_t[49] = 11'b00001000001;
        x_t[50] = 11'b00001001110;
        x_t[51] = 11'b00001010010;
        x_t[52] = 11'b00001001001;
        x_t[53] = 11'b00000111100;
        x_t[54] = 11'b00000101010;
        x_t[55] = 11'b00000110101;
        x_t[56] = 11'b00000111110;
        x_t[57] = 11'b00000111110;
        x_t[58] = 11'b00001000010;
        x_t[59] = 11'b00000101001;
        x_t[60] = 11'b00000101110;
        x_t[61] = 11'b00000110100;
        x_t[62] = 11'b00000100110;
        x_t[63] = 11'b00000101101;
        
        h_t_prev[0] = 11'b00000101110;
        h_t_prev[1] = 11'b00001001001;
        h_t_prev[2] = 11'b00001010010;
        h_t_prev[3] = 11'b00001010101;
        h_t_prev[4] = 11'b00001001111;
        h_t_prev[5] = 11'b00001001100;
        h_t_prev[6] = 11'b00000111111;
        h_t_prev[7] = 11'b00000110111;
        h_t_prev[8] = 11'b00001010001;
        h_t_prev[9] = 11'b00001011010;
        h_t_prev[10] = 11'b00001011011;
        h_t_prev[11] = 11'b00001011111;
        h_t_prev[12] = 11'b00001011010;
        h_t_prev[13] = 11'b00001000000;
        h_t_prev[14] = 11'b00001001101;
        h_t_prev[15] = 11'b00001010111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 2 timeout!");
                $fdisplay(fd_cycles, "Test Vector   2: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   2: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 2");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 3
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000111111;
        x_t[1] = 11'b00001000011;
        x_t[2] = 11'b00001000001;
        x_t[3] = 11'b00001000000;
        x_t[4] = 11'b00000110111;
        x_t[5] = 11'b00000101101;
        x_t[6] = 11'b00000011110;
        x_t[7] = 11'b00000110010;
        x_t[8] = 11'b00001000010;
        x_t[9] = 11'b00001000001;
        x_t[10] = 11'b00001000000;
        x_t[11] = 11'b00001000011;
        x_t[12] = 11'b00000110100;
        x_t[13] = 11'b00000001110;
        x_t[14] = 11'b00001000001;
        x_t[15] = 11'b00001000010;
        x_t[16] = 11'b00001000001;
        x_t[17] = 11'b00001000011;
        x_t[18] = 11'b00001000001;
        x_t[19] = 11'b00000111100;
        x_t[20] = 11'b00000011101;
        x_t[21] = 11'b00000100001;
        x_t[22] = 11'b00000011010;
        x_t[23] = 11'b00000010111;
        x_t[24] = 11'b00000101100;
        x_t[25] = 11'b00000101101;
        x_t[26] = 11'b00000100100;
        x_t[27] = 11'b00000011100;
        x_t[28] = 11'b00000011000;
        x_t[29] = 11'b00000111011;
        x_t[30] = 11'b00000101011;
        x_t[31] = 11'b00000101001;
        x_t[32] = 11'b00000110011;
        x_t[33] = 11'b00000101110;
        x_t[34] = 11'b00000100111;
        x_t[35] = 11'b00000100010;
        x_t[36] = 11'b00000011001;
        x_t[37] = 11'b00000010010;
        x_t[38] = 11'b00000110100;
        x_t[39] = 11'b00000000010;
        x_t[40] = 11'b00000111000;
        x_t[41] = 11'b00000000001;
        x_t[42] = 11'b00000110110;
        x_t[43] = 11'b00000100010;
        x_t[44] = 11'b00000111100;
        x_t[45] = 11'b00000000100;
        x_t[46] = 11'b00000111010;
        x_t[47] = 11'b00000110111;
        x_t[48] = 11'b00000101011;
        x_t[49] = 11'b00000101100;
        x_t[50] = 11'b00000111000;
        x_t[51] = 11'b00000111011;
        x_t[52] = 11'b00000110011;
        x_t[53] = 11'b00000101011;
        x_t[54] = 11'b00000100010;
        x_t[55] = 11'b00000100101;
        x_t[56] = 11'b00000110000;
        x_t[57] = 11'b00000101110;
        x_t[58] = 11'b00000110101;
        x_t[59] = 11'b00000100101;
        x_t[60] = 11'b00000100110;
        x_t[61] = 11'b00000101110;
        x_t[62] = 11'b00000100010;
        x_t[63] = 11'b00000101110;
        
        h_t_prev[0] = 11'b00000111111;
        h_t_prev[1] = 11'b00001000011;
        h_t_prev[2] = 11'b00001000001;
        h_t_prev[3] = 11'b00001000000;
        h_t_prev[4] = 11'b00000110111;
        h_t_prev[5] = 11'b00000101101;
        h_t_prev[6] = 11'b00000011110;
        h_t_prev[7] = 11'b00000110010;
        h_t_prev[8] = 11'b00001000010;
        h_t_prev[9] = 11'b00001000001;
        h_t_prev[10] = 11'b00001000000;
        h_t_prev[11] = 11'b00001000011;
        h_t_prev[12] = 11'b00000110100;
        h_t_prev[13] = 11'b00000001110;
        h_t_prev[14] = 11'b00001000001;
        h_t_prev[15] = 11'b00001000010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 3 timeout!");
                $fdisplay(fd_cycles, "Test Vector   3: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   3: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 3");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 4
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000101101;
        x_t[1] = 11'b00000101111;
        x_t[2] = 11'b00000110100;
        x_t[3] = 11'b00000111010;
        x_t[4] = 11'b00000110001;
        x_t[5] = 11'b00000100100;
        x_t[6] = 11'b00000011100;
        x_t[7] = 11'b00000011111;
        x_t[8] = 11'b00000110001;
        x_t[9] = 11'b00000110101;
        x_t[10] = 11'b00000111000;
        x_t[11] = 11'b00000111100;
        x_t[12] = 11'b00000101011;
        x_t[13] = 11'b00000010001;
        x_t[14] = 11'b00000101110;
        x_t[15] = 11'b00000110110;
        x_t[16] = 11'b00000110101;
        x_t[17] = 11'b00000110110;
        x_t[18] = 11'b00000110111;
        x_t[19] = 11'b00000110010;
        x_t[20] = 11'b00000011100;
        x_t[21] = 11'b00000011011;
        x_t[22] = 11'b00000011001;
        x_t[23] = 11'b00000011111;
        x_t[24] = 11'b00000100000;
        x_t[25] = 11'b00000100010;
        x_t[26] = 11'b00000100110;
        x_t[27] = 11'b00000100010;
        x_t[28] = 11'b00000100100;
        x_t[29] = 11'b00000100001;
        x_t[30] = 11'b00000011111;
        x_t[31] = 11'b00000101000;
        x_t[32] = 11'b00000110001;
        x_t[33] = 11'b00000110000;
        x_t[34] = 11'b00000101100;
        x_t[35] = 11'b00000100101;
        x_t[36] = 11'b00000100011;
        x_t[37] = 11'b00000011011;
        x_t[38] = 11'b00000011100;
        x_t[39] = 11'b00000011100;
        x_t[40] = 11'b00000110001;
        x_t[41] = 11'b00000101101;
        x_t[42] = 11'b00000100001;
        x_t[43] = 11'b00000001101;
        x_t[44] = 11'b00000100010;
        x_t[45] = 11'b00000001111;
        x_t[46] = 11'b00000100011;
        x_t[47] = 11'b00000101001;
        x_t[48] = 11'b00000100011;
        x_t[49] = 11'b00000100100;
        x_t[50] = 11'b00000101100;
        x_t[51] = 11'b00000101110;
        x_t[52] = 11'b00000100111;
        x_t[53] = 11'b00000100100;
        x_t[54] = 11'b00000011111;
        x_t[55] = 11'b00000011101;
        x_t[56] = 11'b00000100111;
        x_t[57] = 11'b00000100111;
        x_t[58] = 11'b00000101100;
        x_t[59] = 11'b00000100001;
        x_t[60] = 11'b00000011101;
        x_t[61] = 11'b00000100111;
        x_t[62] = 11'b00000011010;
        x_t[63] = 11'b00000101110;
        
        h_t_prev[0] = 11'b00000101101;
        h_t_prev[1] = 11'b00000101111;
        h_t_prev[2] = 11'b00000110100;
        h_t_prev[3] = 11'b00000111010;
        h_t_prev[4] = 11'b00000110001;
        h_t_prev[5] = 11'b00000100100;
        h_t_prev[6] = 11'b00000011100;
        h_t_prev[7] = 11'b00000011111;
        h_t_prev[8] = 11'b00000110001;
        h_t_prev[9] = 11'b00000110101;
        h_t_prev[10] = 11'b00000111000;
        h_t_prev[11] = 11'b00000111100;
        h_t_prev[12] = 11'b00000101011;
        h_t_prev[13] = 11'b00000010001;
        h_t_prev[14] = 11'b00000101110;
        h_t_prev[15] = 11'b00000110110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 4 timeout!");
                $fdisplay(fd_cycles, "Test Vector   4: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   4: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 4");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 5
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000011100;
        x_t[1] = 11'b00000100110;
        x_t[2] = 11'b00000101001;
        x_t[3] = 11'b00000110001;
        x_t[4] = 11'b00000101100;
        x_t[5] = 11'b00000100000;
        x_t[6] = 11'b00000011101;
        x_t[7] = 11'b00000010100;
        x_t[8] = 11'b00000100001;
        x_t[9] = 11'b00000100111;
        x_t[10] = 11'b00000101010;
        x_t[11] = 11'b00000110000;
        x_t[12] = 11'b00000100001;
        x_t[13] = 11'b00000010000;
        x_t[14] = 11'b00000100010;
        x_t[15] = 11'b00000101000;
        x_t[16] = 11'b00000101000;
        x_t[17] = 11'b00000101000;
        x_t[18] = 11'b00000100111;
        x_t[19] = 11'b00000100010;
        x_t[20] = 11'b00000010010;
        x_t[21] = 11'b00000011111;
        x_t[22] = 11'b00000010101;
        x_t[23] = 11'b00000011011;
        x_t[24] = 11'b00000010110;
        x_t[25] = 11'b00000010111;
        x_t[26] = 11'b00000100000;
        x_t[27] = 11'b00000011101;
        x_t[28] = 11'b00000011111;
        x_t[29] = 11'b00000001110;
        x_t[30] = 11'b00000011001;
        x_t[31] = 11'b00000100001;
        x_t[32] = 11'b00000101000;
        x_t[33] = 11'b00000100110;
        x_t[34] = 11'b00000100101;
        x_t[35] = 11'b00000011011;
        x_t[36] = 11'b00000011010;
        x_t[37] = 11'b00000010100;
        x_t[38] = 11'b00000001100;
        x_t[39] = 11'b00000001110;
        x_t[40] = 11'b00000000110;
        x_t[41] = 11'b00000001100;
        x_t[42] = 11'b00000000100;
        x_t[43] = 11'b11111111011;
        x_t[44] = 11'b00000010001;
        x_t[45] = 11'b00000000100;
        x_t[46] = 11'b00000011101;
        x_t[47] = 11'b00000100100;
        x_t[48] = 11'b00000011101;
        x_t[49] = 11'b00000011111;
        x_t[50] = 11'b00000100101;
        x_t[51] = 11'b00000100101;
        x_t[52] = 11'b00000011101;
        x_t[53] = 11'b00000011010;
        x_t[54] = 11'b00000010011;
        x_t[55] = 11'b00000011010;
        x_t[56] = 11'b00000100100;
        x_t[57] = 11'b00000100011;
        x_t[58] = 11'b00000100101;
        x_t[59] = 11'b00000011010;
        x_t[60] = 11'b00000011000;
        x_t[61] = 11'b00000100001;
        x_t[62] = 11'b00000010010;
        x_t[63] = 11'b00000101010;
        
        h_t_prev[0] = 11'b00000011100;
        h_t_prev[1] = 11'b00000100110;
        h_t_prev[2] = 11'b00000101001;
        h_t_prev[3] = 11'b00000110001;
        h_t_prev[4] = 11'b00000101100;
        h_t_prev[5] = 11'b00000100000;
        h_t_prev[6] = 11'b00000011101;
        h_t_prev[7] = 11'b00000010100;
        h_t_prev[8] = 11'b00000100001;
        h_t_prev[9] = 11'b00000100111;
        h_t_prev[10] = 11'b00000101010;
        h_t_prev[11] = 11'b00000110000;
        h_t_prev[12] = 11'b00000100001;
        h_t_prev[13] = 11'b00000010000;
        h_t_prev[14] = 11'b00000100010;
        h_t_prev[15] = 11'b00000101000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 5 timeout!");
                $fdisplay(fd_cycles, "Test Vector   5: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   5: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 5");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 6
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000010011;
        x_t[1] = 11'b00000011111;
        x_t[2] = 11'b00000100100;
        x_t[3] = 11'b00000101100;
        x_t[4] = 11'b00000100101;
        x_t[5] = 11'b00000010111;
        x_t[6] = 11'b00000010101;
        x_t[7] = 11'b00000001011;
        x_t[8] = 11'b00000011101;
        x_t[9] = 11'b00000100101;
        x_t[10] = 11'b00000101000;
        x_t[11] = 11'b00000101111;
        x_t[12] = 11'b00000011110;
        x_t[13] = 11'b00000001101;
        x_t[14] = 11'b00000100000;
        x_t[15] = 11'b00000100111;
        x_t[16] = 11'b00000100111;
        x_t[17] = 11'b00000101001;
        x_t[18] = 11'b00000100111;
        x_t[19] = 11'b00000100100;
        x_t[20] = 11'b00000010101;
        x_t[21] = 11'b00000010011;
        x_t[22] = 11'b00000010000;
        x_t[23] = 11'b00000010010;
        x_t[24] = 11'b00000010010;
        x_t[25] = 11'b00000010011;
        x_t[26] = 11'b00000011010;
        x_t[27] = 11'b00000010011;
        x_t[28] = 11'b00000010011;
        x_t[29] = 11'b00000001100;
        x_t[30] = 11'b00000011101;
        x_t[31] = 11'b00000011110;
        x_t[32] = 11'b00000101000;
        x_t[33] = 11'b00000100101;
        x_t[34] = 11'b00000100001;
        x_t[35] = 11'b00000011010;
        x_t[36] = 11'b00000010100;
        x_t[37] = 11'b00000001101;
        x_t[38] = 11'b00000001011;
        x_t[39] = 11'b00000001001;
        x_t[40] = 11'b00000010001;
        x_t[41] = 11'b00000000101;
        x_t[42] = 11'b00000010101;
        x_t[43] = 11'b00000011011;
        x_t[44] = 11'b00000011010;
        x_t[45] = 11'b00000001010;
        x_t[46] = 11'b00000011001;
        x_t[47] = 11'b00000011101;
        x_t[48] = 11'b00000010101;
        x_t[49] = 11'b00000011100;
        x_t[50] = 11'b00000100101;
        x_t[51] = 11'b00000101001;
        x_t[52] = 11'b00000100100;
        x_t[53] = 11'b00000100101;
        x_t[54] = 11'b00000011011;
        x_t[55] = 11'b00000010001;
        x_t[56] = 11'b00000011100;
        x_t[57] = 11'b00000011111;
        x_t[58] = 11'b00000100111;
        x_t[59] = 11'b00000011001;
        x_t[60] = 11'b00000010100;
        x_t[61] = 11'b00000011011;
        x_t[62] = 11'b00000001011;
        x_t[63] = 11'b00000100011;
        
        h_t_prev[0] = 11'b00000010011;
        h_t_prev[1] = 11'b00000011111;
        h_t_prev[2] = 11'b00000100100;
        h_t_prev[3] = 11'b00000101100;
        h_t_prev[4] = 11'b00000100101;
        h_t_prev[5] = 11'b00000010111;
        h_t_prev[6] = 11'b00000010101;
        h_t_prev[7] = 11'b00000001011;
        h_t_prev[8] = 11'b00000011101;
        h_t_prev[9] = 11'b00000100101;
        h_t_prev[10] = 11'b00000101000;
        h_t_prev[11] = 11'b00000101111;
        h_t_prev[12] = 11'b00000011110;
        h_t_prev[13] = 11'b00000001101;
        h_t_prev[14] = 11'b00000100000;
        h_t_prev[15] = 11'b00000100111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 6 timeout!");
                $fdisplay(fd_cycles, "Test Vector   6: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   6: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 6");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 7
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000011001;
        x_t[1] = 11'b00000100101;
        x_t[2] = 11'b00000101100;
        x_t[3] = 11'b00000110101;
        x_t[4] = 11'b00000101111;
        x_t[5] = 11'b00000100010;
        x_t[6] = 11'b00000011100;
        x_t[7] = 11'b00000000110;
        x_t[8] = 11'b00000100000;
        x_t[9] = 11'b00000101011;
        x_t[10] = 11'b00000110001;
        x_t[11] = 11'b00000111010;
        x_t[12] = 11'b00000101111;
        x_t[13] = 11'b00000011100;
        x_t[14] = 11'b00000010011;
        x_t[15] = 11'b00000100101;
        x_t[16] = 11'b00000101000;
        x_t[17] = 11'b00000101010;
        x_t[18] = 11'b00000101110;
        x_t[19] = 11'b00000110010;
        x_t[20] = 11'b00000101001;
        x_t[21] = 11'b00000010001;
        x_t[22] = 11'b00000001111;
        x_t[23] = 11'b00000001111;
        x_t[24] = 11'b00000010110;
        x_t[25] = 11'b00000010111;
        x_t[26] = 11'b00000011101;
        x_t[27] = 11'b00000010110;
        x_t[28] = 11'b00000010010;
        x_t[29] = 11'b00000010001;
        x_t[30] = 11'b00000100100;
        x_t[31] = 11'b00000100011;
        x_t[32] = 11'b00000101010;
        x_t[33] = 11'b00000101010;
        x_t[34] = 11'b00000100110;
        x_t[35] = 11'b00000100000;
        x_t[36] = 11'b00000011101;
        x_t[37] = 11'b00000010100;
        x_t[38] = 11'b00000010011;
        x_t[39] = 11'b00000010011;
        x_t[40] = 11'b00000100000;
        x_t[41] = 11'b00000010011;
        x_t[42] = 11'b00000010101;
        x_t[43] = 11'b00001001010;
        x_t[44] = 11'b00000011001;
        x_t[45] = 11'b00000100001;
        x_t[46] = 11'b00000010011;
        x_t[47] = 11'b00000010101;
        x_t[48] = 11'b00000001101;
        x_t[49] = 11'b00000010100;
        x_t[50] = 11'b00000100011;
        x_t[51] = 11'b00000101101;
        x_t[52] = 11'b00000101111;
        x_t[53] = 11'b00000110011;
        x_t[54] = 11'b00000101111;
        x_t[55] = 11'b00000001001;
        x_t[56] = 11'b00000010101;
        x_t[57] = 11'b00000011011;
        x_t[58] = 11'b00000101101;
        x_t[59] = 11'b00000100000;
        x_t[60] = 11'b00000001110;
        x_t[61] = 11'b00000010100;
        x_t[62] = 11'b00000000111;
        x_t[63] = 11'b00000011000;
        
        h_t_prev[0] = 11'b00000011001;
        h_t_prev[1] = 11'b00000100101;
        h_t_prev[2] = 11'b00000101100;
        h_t_prev[3] = 11'b00000110101;
        h_t_prev[4] = 11'b00000101111;
        h_t_prev[5] = 11'b00000100010;
        h_t_prev[6] = 11'b00000011100;
        h_t_prev[7] = 11'b00000000110;
        h_t_prev[8] = 11'b00000100000;
        h_t_prev[9] = 11'b00000101011;
        h_t_prev[10] = 11'b00000110001;
        h_t_prev[11] = 11'b00000111010;
        h_t_prev[12] = 11'b00000101111;
        h_t_prev[13] = 11'b00000011100;
        h_t_prev[14] = 11'b00000010011;
        h_t_prev[15] = 11'b00000100101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 7 timeout!");
                $fdisplay(fd_cycles, "Test Vector   7: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   7: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 7");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 8
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000011001;
        x_t[1] = 11'b00000100011;
        x_t[2] = 11'b00000101001;
        x_t[3] = 11'b00000110101;
        x_t[4] = 11'b00000110001;
        x_t[5] = 11'b00000100111;
        x_t[6] = 11'b00000100110;
        x_t[7] = 11'b00000001001;
        x_t[8] = 11'b00000011100;
        x_t[9] = 11'b00000100101;
        x_t[10] = 11'b00000101110;
        x_t[11] = 11'b00000111010;
        x_t[12] = 11'b00000110011;
        x_t[13] = 11'b00000100111;
        x_t[14] = 11'b00000010011;
        x_t[15] = 11'b00000100000;
        x_t[16] = 11'b00000100010;
        x_t[17] = 11'b00000100110;
        x_t[18] = 11'b00000101110;
        x_t[19] = 11'b00000110100;
        x_t[20] = 11'b00000110000;
        x_t[21] = 11'b00000010110;
        x_t[22] = 11'b00000010010;
        x_t[23] = 11'b00000010101;
        x_t[24] = 11'b00000010110;
        x_t[25] = 11'b00000011000;
        x_t[26] = 11'b00000100001;
        x_t[27] = 11'b00000011011;
        x_t[28] = 11'b00000011000;
        x_t[29] = 11'b00000010001;
        x_t[30] = 11'b00000100001;
        x_t[31] = 11'b00000100110;
        x_t[32] = 11'b00000101011;
        x_t[33] = 11'b00000101001;
        x_t[34] = 11'b00000100111;
        x_t[35] = 11'b00000100001;
        x_t[36] = 11'b00000100011;
        x_t[37] = 11'b00000011100;
        x_t[38] = 11'b00000001101;
        x_t[39] = 11'b00000011000;
        x_t[40] = 11'b00000011000;
        x_t[41] = 11'b00000011001;
        x_t[42] = 11'b00000001110;
        x_t[43] = 11'b00000101010;
        x_t[44] = 11'b00000001110;
        x_t[45] = 11'b00000100100;
        x_t[46] = 11'b00000001101;
        x_t[47] = 11'b00000010010;
        x_t[48] = 11'b00000001011;
        x_t[49] = 11'b00000010011;
        x_t[50] = 11'b00000100001;
        x_t[51] = 11'b00000101100;
        x_t[52] = 11'b00000101011;
        x_t[53] = 11'b00000110001;
        x_t[54] = 11'b00000101010;
        x_t[55] = 11'b00000001001;
        x_t[56] = 11'b00000010100;
        x_t[57] = 11'b00000011010;
        x_t[58] = 11'b00000101000;
        x_t[59] = 11'b00000010111;
        x_t[60] = 11'b00000001001;
        x_t[61] = 11'b00000001110;
        x_t[62] = 11'b00000000011;
        x_t[63] = 11'b00000001100;
        
        h_t_prev[0] = 11'b00000011001;
        h_t_prev[1] = 11'b00000100011;
        h_t_prev[2] = 11'b00000101001;
        h_t_prev[3] = 11'b00000110101;
        h_t_prev[4] = 11'b00000110001;
        h_t_prev[5] = 11'b00000100111;
        h_t_prev[6] = 11'b00000100110;
        h_t_prev[7] = 11'b00000001001;
        h_t_prev[8] = 11'b00000011100;
        h_t_prev[9] = 11'b00000100101;
        h_t_prev[10] = 11'b00000101110;
        h_t_prev[11] = 11'b00000111010;
        h_t_prev[12] = 11'b00000110011;
        h_t_prev[13] = 11'b00000100111;
        h_t_prev[14] = 11'b00000010011;
        h_t_prev[15] = 11'b00000100000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 8 timeout!");
                $fdisplay(fd_cycles, "Test Vector   8: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   8: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 8");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 9
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000010111;
        x_t[1] = 11'b00000011110;
        x_t[2] = 11'b00000100110;
        x_t[3] = 11'b00000101111;
        x_t[4] = 11'b00000101011;
        x_t[5] = 11'b00000100100;
        x_t[6] = 11'b00000100110;
        x_t[7] = 11'b00000000110;
        x_t[8] = 11'b00000010101;
        x_t[9] = 11'b00000011101;
        x_t[10] = 11'b00000100101;
        x_t[11] = 11'b00000110100;
        x_t[12] = 11'b00000101100;
        x_t[13] = 11'b00000101001;
        x_t[14] = 11'b00000001110;
        x_t[15] = 11'b00000011000;
        x_t[16] = 11'b00000011011;
        x_t[17] = 11'b00000100001;
        x_t[18] = 11'b00000100111;
        x_t[19] = 11'b00000101100;
        x_t[20] = 11'b00000101000;
        x_t[21] = 11'b00000011011;
        x_t[22] = 11'b00000010011;
        x_t[23] = 11'b00000010110;
        x_t[24] = 11'b00000011001;
        x_t[25] = 11'b00000011011;
        x_t[26] = 11'b00000100001;
        x_t[27] = 11'b00000011010;
        x_t[28] = 11'b00000010010;
        x_t[29] = 11'b00000010011;
        x_t[30] = 11'b00000100001;
        x_t[31] = 11'b00000100010;
        x_t[32] = 11'b00000101001;
        x_t[33] = 11'b00000100110;
        x_t[34] = 11'b00000100011;
        x_t[35] = 11'b00000011111;
        x_t[36] = 11'b00000011001;
        x_t[37] = 11'b00000010111;
        x_t[38] = 11'b00000010000;
        x_t[39] = 11'b00000001110;
        x_t[40] = 11'b00000010111;
        x_t[41] = 11'b00000001101;
        x_t[42] = 11'b00000001110;
        x_t[43] = 11'b00000100101;
        x_t[44] = 11'b00000000011;
        x_t[45] = 11'b00000010000;
        x_t[46] = 11'b00000010010;
        x_t[47] = 11'b00000010110;
        x_t[48] = 11'b00000001100;
        x_t[49] = 11'b00000010101;
        x_t[50] = 11'b00000011110;
        x_t[51] = 11'b00000100110;
        x_t[52] = 11'b00000100010;
        x_t[53] = 11'b00000100011;
        x_t[54] = 11'b00000011111;
        x_t[55] = 11'b00000010101;
        x_t[56] = 11'b00000011101;
        x_t[57] = 11'b00000011110;
        x_t[58] = 11'b00000100011;
        x_t[59] = 11'b00000010010;
        x_t[60] = 11'b00000001101;
        x_t[61] = 11'b00000001110;
        x_t[62] = 11'b00000000001;
        x_t[63] = 11'b00000001011;
        
        h_t_prev[0] = 11'b00000010111;
        h_t_prev[1] = 11'b00000011110;
        h_t_prev[2] = 11'b00000100110;
        h_t_prev[3] = 11'b00000101111;
        h_t_prev[4] = 11'b00000101011;
        h_t_prev[5] = 11'b00000100100;
        h_t_prev[6] = 11'b00000100110;
        h_t_prev[7] = 11'b00000000110;
        h_t_prev[8] = 11'b00000010101;
        h_t_prev[9] = 11'b00000011101;
        h_t_prev[10] = 11'b00000100101;
        h_t_prev[11] = 11'b00000110100;
        h_t_prev[12] = 11'b00000101100;
        h_t_prev[13] = 11'b00000101001;
        h_t_prev[14] = 11'b00000001110;
        h_t_prev[15] = 11'b00000011000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 9 timeout!");
                $fdisplay(fd_cycles, "Test Vector   9: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   9: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 9");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 10
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000010001;
        x_t[1] = 11'b00000010011;
        x_t[2] = 11'b00000011010;
        x_t[3] = 11'b00000100010;
        x_t[4] = 11'b00000011111;
        x_t[5] = 11'b00000010011;
        x_t[6] = 11'b00000001110;
        x_t[7] = 11'b00000001000;
        x_t[8] = 11'b00000010000;
        x_t[9] = 11'b00000010100;
        x_t[10] = 11'b00000011010;
        x_t[11] = 11'b00000100101;
        x_t[12] = 11'b00000011010;
        x_t[13] = 11'b00000001001;
        x_t[14] = 11'b00000010011;
        x_t[15] = 11'b00000011010;
        x_t[16] = 11'b00000011001;
        x_t[17] = 11'b00000011010;
        x_t[18] = 11'b00000011011;
        x_t[19] = 11'b00000011100;
        x_t[20] = 11'b00000010011;
        x_t[21] = 11'b00000010100;
        x_t[22] = 11'b00000001100;
        x_t[23] = 11'b00000001111;
        x_t[24] = 11'b00000001101;
        x_t[25] = 11'b00000001111;
        x_t[26] = 11'b00000010011;
        x_t[27] = 11'b00000001101;
        x_t[28] = 11'b00000010001;
        x_t[29] = 11'b00000000111;
        x_t[30] = 11'b00000010011;
        x_t[31] = 11'b00000001111;
        x_t[32] = 11'b00000010110;
        x_t[33] = 11'b00000010011;
        x_t[34] = 11'b00000010000;
        x_t[35] = 11'b00000001001;
        x_t[36] = 11'b00000000010;
        x_t[37] = 11'b00000001001;
        x_t[38] = 11'b00000000111;
        x_t[39] = 11'b11111111010;
        x_t[40] = 11'b00000001001;
        x_t[41] = 11'b11111111101;
        x_t[42] = 11'b00000001100;
        x_t[43] = 11'b00000100011;
        x_t[44] = 11'b00000011000;
        x_t[45] = 11'b00000010011;
        x_t[46] = 11'b00000101010;
        x_t[47] = 11'b00000100010;
        x_t[48] = 11'b00000010011;
        x_t[49] = 11'b00000011011;
        x_t[50] = 11'b00000011101;
        x_t[51] = 11'b00000011111;
        x_t[52] = 11'b00000011001;
        x_t[53] = 11'b00000011100;
        x_t[54] = 11'b00000011100;
        x_t[55] = 11'b00000100011;
        x_t[56] = 11'b00000101010;
        x_t[57] = 11'b00000100010;
        x_t[58] = 11'b00000100001;
        x_t[59] = 11'b00000010101;
        x_t[60] = 11'b00000011000;
        x_t[61] = 11'b00000011001;
        x_t[62] = 11'b00000000110;
        x_t[63] = 11'b00000011001;
        
        h_t_prev[0] = 11'b00000010001;
        h_t_prev[1] = 11'b00000010011;
        h_t_prev[2] = 11'b00000011010;
        h_t_prev[3] = 11'b00000100010;
        h_t_prev[4] = 11'b00000011111;
        h_t_prev[5] = 11'b00000010011;
        h_t_prev[6] = 11'b00000001110;
        h_t_prev[7] = 11'b00000001000;
        h_t_prev[8] = 11'b00000010000;
        h_t_prev[9] = 11'b00000010100;
        h_t_prev[10] = 11'b00000011010;
        h_t_prev[11] = 11'b00000100101;
        h_t_prev[12] = 11'b00000011010;
        h_t_prev[13] = 11'b00000001001;
        h_t_prev[14] = 11'b00000010011;
        h_t_prev[15] = 11'b00000011010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 10 timeout!");
                $fdisplay(fd_cycles, "Test Vector  10: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  10: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 10");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 11
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000000110;
        x_t[1] = 11'b00000000111;
        x_t[2] = 11'b00000001011;
        x_t[3] = 11'b00000010001;
        x_t[4] = 11'b00000001101;
        x_t[5] = 11'b00000000000;
        x_t[6] = 11'b11111111100;
        x_t[7] = 11'b11111111111;
        x_t[8] = 11'b00000001100;
        x_t[9] = 11'b00000001111;
        x_t[10] = 11'b00000010001;
        x_t[11] = 11'b00000010010;
        x_t[12] = 11'b00000001011;
        x_t[13] = 11'b11111111100;
        x_t[14] = 11'b00000011000;
        x_t[15] = 11'b00000011100;
        x_t[16] = 11'b00000011000;
        x_t[17] = 11'b00000010111;
        x_t[18] = 11'b00000010001;
        x_t[19] = 11'b00000010001;
        x_t[20] = 11'b00000001011;
        x_t[21] = 11'b00000000111;
        x_t[22] = 11'b00000000010;
        x_t[23] = 11'b00000000110;
        x_t[24] = 11'b00000000111;
        x_t[25] = 11'b00000001000;
        x_t[26] = 11'b00000000100;
        x_t[27] = 11'b11111111110;
        x_t[28] = 11'b00000000111;
        x_t[29] = 11'b00000000011;
        x_t[30] = 11'b00000001111;
        x_t[31] = 11'b00000000110;
        x_t[32] = 11'b00000001101;
        x_t[33] = 11'b00000001000;
        x_t[34] = 11'b00000000011;
        x_t[35] = 11'b11111111110;
        x_t[36] = 11'b11111110110;
        x_t[37] = 11'b00000000000;
        x_t[38] = 11'b00000001110;
        x_t[39] = 11'b11111110011;
        x_t[40] = 11'b00000011110;
        x_t[41] = 11'b00000010010;
        x_t[42] = 11'b00000100001;
        x_t[43] = 11'b00000000110;
        x_t[44] = 11'b00000100111;
        x_t[45] = 11'b00000001111;
        x_t[46] = 11'b00000101101;
        x_t[47] = 11'b00000101001;
        x_t[48] = 11'b00000010111;
        x_t[49] = 11'b00000011111;
        x_t[50] = 11'b00000011100;
        x_t[51] = 11'b00000011011;
        x_t[52] = 11'b00000010100;
        x_t[53] = 11'b00000011000;
        x_t[54] = 11'b00000011010;
        x_t[55] = 11'b00000101011;
        x_t[56] = 11'b00000110000;
        x_t[57] = 11'b00000100110;
        x_t[58] = 11'b00000011110;
        x_t[59] = 11'b00000010110;
        x_t[60] = 11'b00000100110;
        x_t[61] = 11'b00000100101;
        x_t[62] = 11'b00000001100;
        x_t[63] = 11'b00000101010;
        
        h_t_prev[0] = 11'b00000000110;
        h_t_prev[1] = 11'b00000000111;
        h_t_prev[2] = 11'b00000001011;
        h_t_prev[3] = 11'b00000010001;
        h_t_prev[4] = 11'b00000001101;
        h_t_prev[5] = 11'b00000000000;
        h_t_prev[6] = 11'b11111111100;
        h_t_prev[7] = 11'b11111111111;
        h_t_prev[8] = 11'b00000001100;
        h_t_prev[9] = 11'b00000001111;
        h_t_prev[10] = 11'b00000010001;
        h_t_prev[11] = 11'b00000010010;
        h_t_prev[12] = 11'b00000001011;
        h_t_prev[13] = 11'b11111111100;
        h_t_prev[14] = 11'b00000011000;
        h_t_prev[15] = 11'b00000011100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 11 timeout!");
                $fdisplay(fd_cycles, "Test Vector  11: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  11: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 11");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 12
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000010101;
        x_t[1] = 11'b00000010000;
        x_t[2] = 11'b00000010000;
        x_t[3] = 11'b00000010001;
        x_t[4] = 11'b00000001101;
        x_t[5] = 11'b11111111101;
        x_t[6] = 11'b11111111011;
        x_t[7] = 11'b00000001101;
        x_t[8] = 11'b00000010100;
        x_t[9] = 11'b00000010001;
        x_t[10] = 11'b00000001110;
        x_t[11] = 11'b00000001111;
        x_t[12] = 11'b00000000110;
        x_t[13] = 11'b11111111011;
        x_t[14] = 11'b00000100000;
        x_t[15] = 11'b00000011111;
        x_t[16] = 11'b00000011000;
        x_t[17] = 11'b00000010001;
        x_t[18] = 11'b00000001011;
        x_t[19] = 11'b00000001100;
        x_t[20] = 11'b00000000110;
        x_t[21] = 11'b00000001011;
        x_t[22] = 11'b00000000100;
        x_t[23] = 11'b00000000100;
        x_t[24] = 11'b00000001100;
        x_t[25] = 11'b00000001101;
        x_t[26] = 11'b00000000110;
        x_t[27] = 11'b11111111111;
        x_t[28] = 11'b00000000100;
        x_t[29] = 11'b00000010000;
        x_t[30] = 11'b00000010001;
        x_t[31] = 11'b00000000111;
        x_t[32] = 11'b00000010010;
        x_t[33] = 11'b00000001110;
        x_t[34] = 11'b00000001000;
        x_t[35] = 11'b00000000011;
        x_t[36] = 11'b11111111000;
        x_t[37] = 11'b00000000010;
        x_t[38] = 11'b00000010011;
        x_t[39] = 11'b11111101110;
        x_t[40] = 11'b00000100110;
        x_t[41] = 11'b11111111000;
        x_t[42] = 11'b00000101101;
        x_t[43] = 11'b11111101010;
        x_t[44] = 11'b00000101000;
        x_t[45] = 11'b00000000000;
        x_t[46] = 11'b00000101010;
        x_t[47] = 11'b00000101001;
        x_t[48] = 11'b00000010111;
        x_t[49] = 11'b00000011011;
        x_t[50] = 11'b00000010110;
        x_t[51] = 11'b00000010100;
        x_t[52] = 11'b00000001011;
        x_t[53] = 11'b00000001110;
        x_t[54] = 11'b00000001100;
        x_t[55] = 11'b00000101010;
        x_t[56] = 11'b00000101110;
        x_t[57] = 11'b00000100011;
        x_t[58] = 11'b00000010110;
        x_t[59] = 11'b00000001010;
        x_t[60] = 11'b00000101011;
        x_t[61] = 11'b00000101000;
        x_t[62] = 11'b00000001100;
        x_t[63] = 11'b00000101111;
        
        h_t_prev[0] = 11'b00000010101;
        h_t_prev[1] = 11'b00000010000;
        h_t_prev[2] = 11'b00000010000;
        h_t_prev[3] = 11'b00000010001;
        h_t_prev[4] = 11'b00000001101;
        h_t_prev[5] = 11'b11111111101;
        h_t_prev[6] = 11'b11111111011;
        h_t_prev[7] = 11'b00000001101;
        h_t_prev[8] = 11'b00000010100;
        h_t_prev[9] = 11'b00000010001;
        h_t_prev[10] = 11'b00000001110;
        h_t_prev[11] = 11'b00000001111;
        h_t_prev[12] = 11'b00000000110;
        h_t_prev[13] = 11'b11111111011;
        h_t_prev[14] = 11'b00000100000;
        h_t_prev[15] = 11'b00000011111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 12 timeout!");
                $fdisplay(fd_cycles, "Test Vector  12: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  12: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 12");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 13
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000010101;
        x_t[1] = 11'b00000010010;
        x_t[2] = 11'b00000010001;
        x_t[3] = 11'b00000010010;
        x_t[4] = 11'b00000001010;
        x_t[5] = 11'b11111111001;
        x_t[6] = 11'b11111111000;
        x_t[7] = 11'b00000010000;
        x_t[8] = 11'b00000010010;
        x_t[9] = 11'b00000001110;
        x_t[10] = 11'b00000001101;
        x_t[11] = 11'b00000001101;
        x_t[12] = 11'b00000000000;
        x_t[13] = 11'b11111110010;
        x_t[14] = 11'b00000100000;
        x_t[15] = 11'b00000011100;
        x_t[16] = 11'b00000010100;
        x_t[17] = 11'b00000001100;
        x_t[18] = 11'b00000001001;
        x_t[19] = 11'b00000001001;
        x_t[20] = 11'b00000000000;
        x_t[21] = 11'b00000001100;
        x_t[22] = 11'b00000000001;
        x_t[23] = 11'b00000000010;
        x_t[24] = 11'b00000001111;
        x_t[25] = 11'b00000010000;
        x_t[26] = 11'b00000000100;
        x_t[27] = 11'b11111111110;
        x_t[28] = 11'b00000000100;
        x_t[29] = 11'b00000010110;
        x_t[30] = 11'b00000001011;
        x_t[31] = 11'b00000000110;
        x_t[32] = 11'b00000001111;
        x_t[33] = 11'b00000001001;
        x_t[34] = 11'b00000000011;
        x_t[35] = 11'b11111111100;
        x_t[36] = 11'b11111110111;
        x_t[37] = 11'b00000000010;
        x_t[38] = 11'b00000011000;
        x_t[39] = 11'b11111100111;
        x_t[40] = 11'b00000101011;
        x_t[41] = 11'b11111100010;
        x_t[42] = 11'b00000100110;
        x_t[43] = 11'b00000110000;
        x_t[44] = 11'b00000100111;
        x_t[45] = 11'b11111111101;
        x_t[46] = 11'b00000100101;
        x_t[47] = 11'b00000100010;
        x_t[48] = 11'b00000010010;
        x_t[49] = 11'b00000011000;
        x_t[50] = 11'b00000010101;
        x_t[51] = 11'b00000010011;
        x_t[52] = 11'b00000001010;
        x_t[53] = 11'b00000001011;
        x_t[54] = 11'b00000000100;
        x_t[55] = 11'b00000011101;
        x_t[56] = 11'b00000100100;
        x_t[57] = 11'b00000011100;
        x_t[58] = 11'b00000010000;
        x_t[59] = 11'b00000000010;
        x_t[60] = 11'b00000100100;
        x_t[61] = 11'b00000100001;
        x_t[62] = 11'b00000000100;
        x_t[63] = 11'b00000100000;
        
        h_t_prev[0] = 11'b00000010101;
        h_t_prev[1] = 11'b00000010010;
        h_t_prev[2] = 11'b00000010001;
        h_t_prev[3] = 11'b00000010010;
        h_t_prev[4] = 11'b00000001010;
        h_t_prev[5] = 11'b11111111001;
        h_t_prev[6] = 11'b11111111000;
        h_t_prev[7] = 11'b00000010000;
        h_t_prev[8] = 11'b00000010010;
        h_t_prev[9] = 11'b00000001110;
        h_t_prev[10] = 11'b00000001101;
        h_t_prev[11] = 11'b00000001101;
        h_t_prev[12] = 11'b00000000000;
        h_t_prev[13] = 11'b11111110010;
        h_t_prev[14] = 11'b00000100000;
        h_t_prev[15] = 11'b00000011100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 13 timeout!");
                $fdisplay(fd_cycles, "Test Vector  13: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  13: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 13");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 14
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000001111;
        x_t[1] = 11'b00000000110;
        x_t[2] = 11'b00000001000;
        x_t[3] = 11'b00000001101;
        x_t[4] = 11'b11111111110;
        x_t[5] = 11'b11111101101;
        x_t[6] = 11'b11111101110;
        x_t[7] = 11'b00000000001;
        x_t[8] = 11'b00000000111;
        x_t[9] = 11'b00000000110;
        x_t[10] = 11'b00000001000;
        x_t[11] = 11'b00000000100;
        x_t[12] = 11'b11111110101;
        x_t[13] = 11'b11111101100;
        x_t[14] = 11'b00000001111;
        x_t[15] = 11'b00000001111;
        x_t[16] = 11'b00000001001;
        x_t[17] = 11'b00000000101;
        x_t[18] = 11'b00000000010;
        x_t[19] = 11'b00000000001;
        x_t[20] = 11'b11111110111;
        x_t[21] = 11'b00000000111;
        x_t[22] = 11'b11111110101;
        x_t[23] = 11'b11111110111;
        x_t[24] = 11'b00000001011;
        x_t[25] = 11'b00000001100;
        x_t[26] = 11'b11111110100;
        x_t[27] = 11'b11111101110;
        x_t[28] = 11'b11111110111;
        x_t[29] = 11'b00000001110;
        x_t[30] = 11'b00000000101;
        x_t[31] = 11'b11111111001;
        x_t[32] = 11'b00000000100;
        x_t[33] = 11'b11111111001;
        x_t[34] = 11'b11111110010;
        x_t[35] = 11'b11111101111;
        x_t[36] = 11'b11111100101;
        x_t[37] = 11'b11111110101;
        x_t[38] = 11'b00000010110;
        x_t[39] = 11'b11111011010;
        x_t[40] = 11'b00000100100;
        x_t[41] = 11'b11111101001;
        x_t[42] = 11'b00000001100;
        x_t[43] = 11'b00000101011;
        x_t[44] = 11'b00000010000;
        x_t[45] = 11'b11111011001;
        x_t[46] = 11'b00000001110;
        x_t[47] = 11'b00000001111;
        x_t[48] = 11'b00000000010;
        x_t[49] = 11'b00000001001;
        x_t[50] = 11'b00000000111;
        x_t[51] = 11'b00000000101;
        x_t[52] = 11'b11111111011;
        x_t[53] = 11'b11111111000;
        x_t[54] = 11'b11111101011;
        x_t[55] = 11'b00000001100;
        x_t[56] = 11'b00000010011;
        x_t[57] = 11'b00000001111;
        x_t[58] = 11'b00000000010;
        x_t[59] = 11'b11111110110;
        x_t[60] = 11'b00000010101;
        x_t[61] = 11'b00000010000;
        x_t[62] = 11'b11111110100;
        x_t[63] = 11'b00000001000;
        
        h_t_prev[0] = 11'b00000001111;
        h_t_prev[1] = 11'b00000000110;
        h_t_prev[2] = 11'b00000001000;
        h_t_prev[3] = 11'b00000001101;
        h_t_prev[4] = 11'b11111111110;
        h_t_prev[5] = 11'b11111101101;
        h_t_prev[6] = 11'b11111101110;
        h_t_prev[7] = 11'b00000000001;
        h_t_prev[8] = 11'b00000000111;
        h_t_prev[9] = 11'b00000000110;
        h_t_prev[10] = 11'b00000001000;
        h_t_prev[11] = 11'b00000000100;
        h_t_prev[12] = 11'b11111110101;
        h_t_prev[13] = 11'b11111101100;
        h_t_prev[14] = 11'b00000001111;
        h_t_prev[15] = 11'b00000001111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 14 timeout!");
                $fdisplay(fd_cycles, "Test Vector  14: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  14: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 14");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 15
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000010100;
        x_t[1] = 11'b00000001011;
        x_t[2] = 11'b00000001011;
        x_t[3] = 11'b00000001110;
        x_t[4] = 11'b00000000001;
        x_t[5] = 11'b11111101110;
        x_t[6] = 11'b11111100111;
        x_t[7] = 11'b00000001101;
        x_t[8] = 11'b00000010000;
        x_t[9] = 11'b00000010001;
        x_t[10] = 11'b00000010011;
        x_t[11] = 11'b00000010001;
        x_t[12] = 11'b11111111101;
        x_t[13] = 11'b11111110000;
        x_t[14] = 11'b00000010101;
        x_t[15] = 11'b00000011001;
        x_t[16] = 11'b00000010011;
        x_t[17] = 11'b00000010001;
        x_t[18] = 11'b00000010000;
        x_t[19] = 11'b00000001110;
        x_t[20] = 11'b11111111111;
        x_t[21] = 11'b00000000011;
        x_t[22] = 11'b11111110111;
        x_t[23] = 11'b11111111011;
        x_t[24] = 11'b00000001001;
        x_t[25] = 11'b00000001011;
        x_t[26] = 11'b11111111101;
        x_t[27] = 11'b11111110011;
        x_t[28] = 11'b11111111011;
        x_t[29] = 11'b00000001111;
        x_t[30] = 11'b00000000111;
        x_t[31] = 11'b00000000100;
        x_t[32] = 11'b00000010010;
        x_t[33] = 11'b00000001011;
        x_t[34] = 11'b00000000010;
        x_t[35] = 11'b11111111110;
        x_t[36] = 11'b11111110010;
        x_t[37] = 11'b00000000110;
        x_t[38] = 11'b00000011100;
        x_t[39] = 11'b11111110000;
        x_t[40] = 11'b00000100000;
        x_t[41] = 11'b00000001100;
        x_t[42] = 11'b00000011001;
        x_t[43] = 11'b00000011011;
        x_t[44] = 11'b00000010111;
        x_t[45] = 11'b00000001100;
        x_t[46] = 11'b00000011001;
        x_t[47] = 11'b00000011101;
        x_t[48] = 11'b00000010001;
        x_t[49] = 11'b00000011010;
        x_t[50] = 11'b00000011011;
        x_t[51] = 11'b00000011001;
        x_t[52] = 11'b00000010001;
        x_t[53] = 11'b00000010000;
        x_t[54] = 11'b00000001101;
        x_t[55] = 11'b00000011000;
        x_t[56] = 11'b00000100001;
        x_t[57] = 11'b00000011101;
        x_t[58] = 11'b00000010010;
        x_t[59] = 11'b00000000101;
        x_t[60] = 11'b00000010001;
        x_t[61] = 11'b00000001111;
        x_t[62] = 11'b11111110011;
        x_t[63] = 11'b00000001000;
        
        h_t_prev[0] = 11'b00000010100;
        h_t_prev[1] = 11'b00000001011;
        h_t_prev[2] = 11'b00000001011;
        h_t_prev[3] = 11'b00000001110;
        h_t_prev[4] = 11'b00000000001;
        h_t_prev[5] = 11'b11111101110;
        h_t_prev[6] = 11'b11111100111;
        h_t_prev[7] = 11'b00000001101;
        h_t_prev[8] = 11'b00000010000;
        h_t_prev[9] = 11'b00000010001;
        h_t_prev[10] = 11'b00000010011;
        h_t_prev[11] = 11'b00000010001;
        h_t_prev[12] = 11'b11111111101;
        h_t_prev[13] = 11'b11111110000;
        h_t_prev[14] = 11'b00000010101;
        h_t_prev[15] = 11'b00000011001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 15 timeout!");
                $fdisplay(fd_cycles, "Test Vector  15: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  15: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 15");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 16
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000011010;
        x_t[1] = 11'b00000011001;
        x_t[2] = 11'b00000011100;
        x_t[3] = 11'b00000100000;
        x_t[4] = 11'b00000011001;
        x_t[5] = 11'b00000000101;
        x_t[6] = 11'b11111111101;
        x_t[7] = 11'b00000010111;
        x_t[8] = 11'b00000011101;
        x_t[9] = 11'b00000011110;
        x_t[10] = 11'b00000100011;
        x_t[11] = 11'b00000100100;
        x_t[12] = 11'b00000010111;
        x_t[13] = 11'b00000001001;
        x_t[14] = 11'b00000100101;
        x_t[15] = 11'b00000100100;
        x_t[16] = 11'b00000100011;
        x_t[17] = 11'b00000100001;
        x_t[18] = 11'b00000100001;
        x_t[19] = 11'b00000100000;
        x_t[20] = 11'b00000010011;
        x_t[21] = 11'b00000001000;
        x_t[22] = 11'b00000000001;
        x_t[23] = 11'b00000000010;
        x_t[24] = 11'b00000001001;
        x_t[25] = 11'b00000001100;
        x_t[26] = 11'b00000001000;
        x_t[27] = 11'b11111111100;
        x_t[28] = 11'b00000000000;
        x_t[29] = 11'b00000001110;
        x_t[30] = 11'b00000000111;
        x_t[31] = 11'b00000001011;
        x_t[32] = 11'b00000010110;
        x_t[33] = 11'b00000010000;
        x_t[34] = 11'b00000001010;
        x_t[35] = 11'b00000000010;
        x_t[36] = 11'b11111111000;
        x_t[37] = 11'b00000001011;
        x_t[38] = 11'b00000001101;
        x_t[39] = 11'b11111111000;
        x_t[40] = 11'b00000001111;
        x_t[41] = 11'b00000001100;
        x_t[42] = 11'b00000011001;
        x_t[43] = 11'b00000011110;
        x_t[44] = 11'b00000010101;
        x_t[45] = 11'b00000010101;
        x_t[46] = 11'b00000011111;
        x_t[47] = 11'b00000100010;
        x_t[48] = 11'b00000010010;
        x_t[49] = 11'b00000011110;
        x_t[50] = 11'b00000011110;
        x_t[51] = 11'b00000011101;
        x_t[52] = 11'b00000010111;
        x_t[53] = 11'b00000010011;
        x_t[54] = 11'b00000001010;
        x_t[55] = 11'b00000011101;
        x_t[56] = 11'b00000100101;
        x_t[57] = 11'b00000100000;
        x_t[58] = 11'b00000010110;
        x_t[59] = 11'b00000000110;
        x_t[60] = 11'b00000011001;
        x_t[61] = 11'b00000011001;
        x_t[62] = 11'b11111111111;
        x_t[63] = 11'b00000010101;
        
        h_t_prev[0] = 11'b00000011010;
        h_t_prev[1] = 11'b00000011001;
        h_t_prev[2] = 11'b00000011100;
        h_t_prev[3] = 11'b00000100000;
        h_t_prev[4] = 11'b00000011001;
        h_t_prev[5] = 11'b00000000101;
        h_t_prev[6] = 11'b11111111101;
        h_t_prev[7] = 11'b00000010111;
        h_t_prev[8] = 11'b00000011101;
        h_t_prev[9] = 11'b00000011110;
        h_t_prev[10] = 11'b00000100011;
        h_t_prev[11] = 11'b00000100100;
        h_t_prev[12] = 11'b00000010111;
        h_t_prev[13] = 11'b00000001001;
        h_t_prev[14] = 11'b00000100101;
        h_t_prev[15] = 11'b00000100100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 16 timeout!");
                $fdisplay(fd_cycles, "Test Vector  16: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  16: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 16");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 17
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000000101;
        x_t[1] = 11'b00000000111;
        x_t[2] = 11'b11111101000;
        x_t[3] = 11'b11111110000;
        x_t[4] = 11'b11111101101;
        x_t[5] = 11'b11111101001;
        x_t[6] = 11'b11111110100;
        x_t[7] = 11'b00000010001;
        x_t[8] = 11'b00000000001;
        x_t[9] = 11'b11111110100;
        x_t[10] = 11'b11111101100;
        x_t[11] = 11'b11111011111;
        x_t[12] = 11'b11111100010;
        x_t[13] = 11'b11111100110;
        x_t[14] = 11'b00000011000;
        x_t[15] = 11'b00000001001;
        x_t[16] = 11'b11111111000;
        x_t[17] = 11'b11111110000;
        x_t[18] = 11'b11111011111;
        x_t[19] = 11'b11111100000;
        x_t[20] = 11'b11111101010;
        x_t[21] = 11'b11111111111;
        x_t[22] = 11'b00000001000;
        x_t[23] = 11'b00000001010;
        x_t[24] = 11'b00000000110;
        x_t[25] = 11'b00000000101;
        x_t[26] = 11'b11111110001;
        x_t[27] = 11'b11111111000;
        x_t[28] = 11'b00000001111;
        x_t[29] = 11'b00000000011;
        x_t[30] = 11'b00000010010;
        x_t[31] = 11'b11111111110;
        x_t[32] = 11'b11111111001;
        x_t[33] = 11'b11111110101;
        x_t[34] = 11'b11111110011;
        x_t[35] = 11'b11111101110;
        x_t[36] = 11'b11111111110;
        x_t[37] = 11'b11111011001;
        x_t[38] = 11'b00000001001;
        x_t[39] = 11'b00000000100;
        x_t[40] = 11'b00000010001;
        x_t[41] = 11'b00000000111;
        x_t[42] = 11'b00000011000;
        x_t[43] = 11'b11111111110;
        x_t[44] = 11'b00000011100;
        x_t[45] = 11'b00000000000;
        x_t[46] = 11'b00000011011;
        x_t[47] = 11'b00000010110;
        x_t[48] = 11'b00000001110;
        x_t[49] = 11'b00000000101;
        x_t[50] = 11'b11111110101;
        x_t[51] = 11'b11111101111;
        x_t[52] = 11'b11111110001;
        x_t[53] = 11'b11111110111;
        x_t[54] = 11'b00000001010;
        x_t[55] = 11'b00000001110;
        x_t[56] = 11'b00000010101;
        x_t[57] = 11'b11111111010;
        x_t[58] = 11'b11111111001;
        x_t[59] = 11'b00000010101;
        x_t[60] = 11'b00000000011;
        x_t[61] = 11'b11111111010;
        x_t[62] = 11'b11111111101;
        x_t[63] = 11'b00000001000;
        
        h_t_prev[0] = 11'b00000000101;
        h_t_prev[1] = 11'b00000000111;
        h_t_prev[2] = 11'b11111101000;
        h_t_prev[3] = 11'b11111110000;
        h_t_prev[4] = 11'b11111101101;
        h_t_prev[5] = 11'b11111101001;
        h_t_prev[6] = 11'b11111110100;
        h_t_prev[7] = 11'b00000010001;
        h_t_prev[8] = 11'b00000000001;
        h_t_prev[9] = 11'b11111110100;
        h_t_prev[10] = 11'b11111101100;
        h_t_prev[11] = 11'b11111011111;
        h_t_prev[12] = 11'b11111100010;
        h_t_prev[13] = 11'b11111100110;
        h_t_prev[14] = 11'b00000011000;
        h_t_prev[15] = 11'b00000001001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 17 timeout!");
                $fdisplay(fd_cycles, "Test Vector  17: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  17: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 17");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 18
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000010101;
        x_t[1] = 11'b00000011000;
        x_t[2] = 11'b00000000000;
        x_t[3] = 11'b00000000101;
        x_t[4] = 11'b11111111101;
        x_t[5] = 11'b11111111001;
        x_t[6] = 11'b11111111110;
        x_t[7] = 11'b00000100110;
        x_t[8] = 11'b00000010010;
        x_t[9] = 11'b00000000111;
        x_t[10] = 11'b00000000000;
        x_t[11] = 11'b11111110110;
        x_t[12] = 11'b11111111000;
        x_t[13] = 11'b11111111011;
        x_t[14] = 11'b00000011000;
        x_t[15] = 11'b00000010100;
        x_t[16] = 11'b00000001000;
        x_t[17] = 11'b00000000110;
        x_t[18] = 11'b11111110110;
        x_t[19] = 11'b11111111010;
        x_t[20] = 11'b00000000000;
        x_t[21] = 11'b00000000001;
        x_t[22] = 11'b00000001010;
        x_t[23] = 11'b00000001101;
        x_t[24] = 11'b00000001011;
        x_t[25] = 11'b00000001011;
        x_t[26] = 11'b11111111100;
        x_t[27] = 11'b11111111111;
        x_t[28] = 11'b00000010000;
        x_t[29] = 11'b00000001111;
        x_t[30] = 11'b00000011110;
        x_t[31] = 11'b00000001000;
        x_t[32] = 11'b00000001001;
        x_t[33] = 11'b00000000010;
        x_t[34] = 11'b11111111101;
        x_t[35] = 11'b11111111011;
        x_t[36] = 11'b00000000010;
        x_t[37] = 11'b11111010101;
        x_t[38] = 11'b00000011101;
        x_t[39] = 11'b00000000110;
        x_t[40] = 11'b00000100111;
        x_t[41] = 11'b11111110011;
        x_t[42] = 11'b00000011001;
        x_t[43] = 11'b00000010100;
        x_t[44] = 11'b00000011100;
        x_t[45] = 11'b00000001010;
        x_t[46] = 11'b00000010000;
        x_t[47] = 11'b00000010011;
        x_t[48] = 11'b00000001110;
        x_t[49] = 11'b00000001001;
        x_t[50] = 11'b00000000010;
        x_t[51] = 11'b00000000001;
        x_t[52] = 11'b00000000010;
        x_t[53] = 11'b00000000100;
        x_t[54] = 11'b00000010010;
        x_t[55] = 11'b00000001001;
        x_t[56] = 11'b00000001111;
        x_t[57] = 11'b00000000000;
        x_t[58] = 11'b00000001010;
        x_t[59] = 11'b00000010110;
        x_t[60] = 11'b11111111100;
        x_t[61] = 11'b11111111101;
        x_t[62] = 11'b00000001001;
        x_t[63] = 11'b11111110111;
        
        h_t_prev[0] = 11'b00000010101;
        h_t_prev[1] = 11'b00000011000;
        h_t_prev[2] = 11'b00000000000;
        h_t_prev[3] = 11'b00000000101;
        h_t_prev[4] = 11'b11111111101;
        h_t_prev[5] = 11'b11111111001;
        h_t_prev[6] = 11'b11111111110;
        h_t_prev[7] = 11'b00000100110;
        h_t_prev[8] = 11'b00000010010;
        h_t_prev[9] = 11'b00000000111;
        h_t_prev[10] = 11'b00000000000;
        h_t_prev[11] = 11'b11111110110;
        h_t_prev[12] = 11'b11111111000;
        h_t_prev[13] = 11'b11111111011;
        h_t_prev[14] = 11'b00000011000;
        h_t_prev[15] = 11'b00000010100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 18 timeout!");
                $fdisplay(fd_cycles, "Test Vector  18: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  18: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 18");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 19
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000100101;
        x_t[1] = 11'b00000100001;
        x_t[2] = 11'b00000001010;
        x_t[3] = 11'b00000001011;
        x_t[4] = 11'b00000000001;
        x_t[5] = 11'b11111111101;
        x_t[6] = 11'b11111111101;
        x_t[7] = 11'b00000101010;
        x_t[8] = 11'b00000010100;
        x_t[9] = 11'b00000001100;
        x_t[10] = 11'b00000000100;
        x_t[11] = 11'b00000000001;
        x_t[12] = 11'b00000000010;
        x_t[13] = 11'b11111111011;
        x_t[14] = 11'b00000011100;
        x_t[15] = 11'b00000010110;
        x_t[16] = 11'b00000001011;
        x_t[17] = 11'b00000001101;
        x_t[18] = 11'b00000000101;
        x_t[19] = 11'b00000001011;
        x_t[20] = 11'b00000001110;
        x_t[21] = 11'b00000010100;
        x_t[22] = 11'b00000011001;
        x_t[23] = 11'b00000010110;
        x_t[24] = 11'b00000100100;
        x_t[25] = 11'b00000100010;
        x_t[26] = 11'b00000001000;
        x_t[27] = 11'b00000000110;
        x_t[28] = 11'b00000010011;
        x_t[29] = 11'b00000101000;
        x_t[30] = 11'b00000110111;
        x_t[31] = 11'b00000010101;
        x_t[32] = 11'b00000011000;
        x_t[33] = 11'b00000001111;
        x_t[34] = 11'b00000001001;
        x_t[35] = 11'b00000000110;
        x_t[36] = 11'b00000000011;
        x_t[37] = 11'b11111001110;
        x_t[38] = 11'b00000111001;
        x_t[39] = 11'b11111111110;
        x_t[40] = 11'b00000110111;
        x_t[41] = 11'b11111100001;
        x_t[42] = 11'b00000101110;
        x_t[43] = 11'b00000000001;
        x_t[44] = 11'b00000101001;
        x_t[45] = 11'b00000101010;
        x_t[46] = 11'b00000011110;
        x_t[47] = 11'b00000100000;
        x_t[48] = 11'b00000100000;
        x_t[49] = 11'b00000011011;
        x_t[50] = 11'b00000011100;
        x_t[51] = 11'b00000100011;
        x_t[52] = 11'b00000101000;
        x_t[53] = 11'b00000101001;
        x_t[54] = 11'b00000110000;
        x_t[55] = 11'b00000010111;
        x_t[56] = 11'b00000011101;
        x_t[57] = 11'b00000011100;
        x_t[58] = 11'b00000110000;
        x_t[59] = 11'b00000101110;
        x_t[60] = 11'b11111111100;
        x_t[61] = 11'b00000000100;
        x_t[62] = 11'b00000010000;
        x_t[63] = 11'b11111101000;
        
        h_t_prev[0] = 11'b00000100101;
        h_t_prev[1] = 11'b00000100001;
        h_t_prev[2] = 11'b00000001010;
        h_t_prev[3] = 11'b00000001011;
        h_t_prev[4] = 11'b00000000001;
        h_t_prev[5] = 11'b11111111101;
        h_t_prev[6] = 11'b11111111101;
        h_t_prev[7] = 11'b00000101010;
        h_t_prev[8] = 11'b00000010100;
        h_t_prev[9] = 11'b00000001100;
        h_t_prev[10] = 11'b00000000100;
        h_t_prev[11] = 11'b00000000001;
        h_t_prev[12] = 11'b00000000010;
        h_t_prev[13] = 11'b11111111011;
        h_t_prev[14] = 11'b00000011100;
        h_t_prev[15] = 11'b00000010110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 19 timeout!");
                $fdisplay(fd_cycles, "Test Vector  19: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  19: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 19");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 20
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000111001;
        x_t[1] = 11'b00000110110;
        x_t[2] = 11'b00000011111;
        x_t[3] = 11'b00000011100;
        x_t[4] = 11'b00000010111;
        x_t[5] = 11'b00000010110;
        x_t[6] = 11'b00000010000;
        x_t[7] = 11'b00000111011;
        x_t[8] = 11'b00000101010;
        x_t[9] = 11'b00000100101;
        x_t[10] = 11'b00000100001;
        x_t[11] = 11'b00000011101;
        x_t[12] = 11'b00000100110;
        x_t[13] = 11'b00000100000;
        x_t[14] = 11'b00000110001;
        x_t[15] = 11'b00000101111;
        x_t[16] = 11'b00000100101;
        x_t[17] = 11'b00000100111;
        x_t[18] = 11'b00000101010;
        x_t[19] = 11'b00000110011;
        x_t[20] = 11'b00000111001;
        x_t[21] = 11'b00000011000;
        x_t[22] = 11'b00000011001;
        x_t[23] = 11'b00000010110;
        x_t[24] = 11'b00000100011;
        x_t[25] = 11'b00000100011;
        x_t[26] = 11'b00000010000;
        x_t[27] = 11'b00000001011;
        x_t[28] = 11'b00000010100;
        x_t[29] = 11'b00000011111;
        x_t[30] = 11'b00000111000;
        x_t[31] = 11'b00000011001;
        x_t[32] = 11'b00000011010;
        x_t[33] = 11'b00000010100;
        x_t[34] = 11'b00000001111;
        x_t[35] = 11'b00000001011;
        x_t[36] = 11'b00000001011;
        x_t[37] = 11'b11111010110;
        x_t[38] = 11'b00000101101;
        x_t[39] = 11'b00000010011;
        x_t[40] = 11'b00000101101;
        x_t[41] = 11'b00000001110;
        x_t[42] = 11'b00000101001;
        x_t[43] = 11'b11111111110;
        x_t[44] = 11'b00000101100;
        x_t[45] = 11'b00001000011;
        x_t[46] = 11'b00000100110;
        x_t[47] = 11'b00000100100;
        x_t[48] = 11'b00000100011;
        x_t[49] = 11'b00000100011;
        x_t[50] = 11'b00000100110;
        x_t[51] = 11'b00000111000;
        x_t[52] = 11'b00000111101;
        x_t[53] = 11'b00000111110;
        x_t[54] = 11'b00001000000;
        x_t[55] = 11'b00000011001;
        x_t[56] = 11'b00000011100;
        x_t[57] = 11'b00000100111;
        x_t[58] = 11'b00001000100;
        x_t[59] = 11'b00000111010;
        x_t[60] = 11'b00000000100;
        x_t[61] = 11'b00000010101;
        x_t[62] = 11'b00000100001;
        x_t[63] = 11'b11111110100;
        
        h_t_prev[0] = 11'b00000111001;
        h_t_prev[1] = 11'b00000110110;
        h_t_prev[2] = 11'b00000011111;
        h_t_prev[3] = 11'b00000011100;
        h_t_prev[4] = 11'b00000010111;
        h_t_prev[5] = 11'b00000010110;
        h_t_prev[6] = 11'b00000010000;
        h_t_prev[7] = 11'b00000111011;
        h_t_prev[8] = 11'b00000101010;
        h_t_prev[9] = 11'b00000100101;
        h_t_prev[10] = 11'b00000100001;
        h_t_prev[11] = 11'b00000011101;
        h_t_prev[12] = 11'b00000100110;
        h_t_prev[13] = 11'b00000100000;
        h_t_prev[14] = 11'b00000110001;
        h_t_prev[15] = 11'b00000101111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 20 timeout!");
                $fdisplay(fd_cycles, "Test Vector  20: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  20: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 20");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 21
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000010111;
        x_t[1] = 11'b00000011001;
        x_t[2] = 11'b00000001000;
        x_t[3] = 11'b00000001001;
        x_t[4] = 11'b00000001101;
        x_t[5] = 11'b00000010000;
        x_t[6] = 11'b00000010101;
        x_t[7] = 11'b00000011010;
        x_t[8] = 11'b00000010000;
        x_t[9] = 11'b00000001110;
        x_t[10] = 11'b00000001110;
        x_t[11] = 11'b00000010000;
        x_t[12] = 11'b00000100100;
        x_t[13] = 11'b00000100110;
        x_t[14] = 11'b00000011000;
        x_t[15] = 11'b00000010111;
        x_t[16] = 11'b00000010010;
        x_t[17] = 11'b00000010111;
        x_t[18] = 11'b00000011101;
        x_t[19] = 11'b00000101011;
        x_t[20] = 11'b00000110110;
        x_t[21] = 11'b11111110111;
        x_t[22] = 11'b00000000001;
        x_t[23] = 11'b00000001011;
        x_t[24] = 11'b11111111010;
        x_t[25] = 11'b11111111010;
        x_t[26] = 11'b11111111001;
        x_t[27] = 11'b00000000001;
        x_t[28] = 11'b00000001101;
        x_t[29] = 11'b11111110110;
        x_t[30] = 11'b00000001001;
        x_t[31] = 11'b00000000111;
        x_t[32] = 11'b11111111011;
        x_t[33] = 11'b11111111011;
        x_t[34] = 11'b11111111110;
        x_t[35] = 11'b11111110111;
        x_t[36] = 11'b00000001011;
        x_t[37] = 11'b11111011100;
        x_t[38] = 11'b11111111101;
        x_t[39] = 11'b00000011000;
        x_t[40] = 11'b00000010011;
        x_t[41] = 11'b00000010111;
        x_t[42] = 11'b00000000100;
        x_t[43] = 11'b00000100111;
        x_t[44] = 11'b00000010001;
        x_t[45] = 11'b00000110001;
        x_t[46] = 11'b00000010010;
        x_t[47] = 11'b00000010010;
        x_t[48] = 11'b00000010001;
        x_t[49] = 11'b00000010011;
        x_t[50] = 11'b00000011011;
        x_t[51] = 11'b00000101101;
        x_t[52] = 11'b00000110000;
        x_t[53] = 11'b00000110001;
        x_t[54] = 11'b00000101010;
        x_t[55] = 11'b00000001111;
        x_t[56] = 11'b00000010011;
        x_t[57] = 11'b00000100001;
        x_t[58] = 11'b00000111001;
        x_t[59] = 11'b00000101110;
        x_t[60] = 11'b00000000111;
        x_t[61] = 11'b00000100010;
        x_t[62] = 11'b00000101101;
        x_t[63] = 11'b00000000011;
        
        h_t_prev[0] = 11'b00000010111;
        h_t_prev[1] = 11'b00000011001;
        h_t_prev[2] = 11'b00000001000;
        h_t_prev[3] = 11'b00000001001;
        h_t_prev[4] = 11'b00000001101;
        h_t_prev[5] = 11'b00000010000;
        h_t_prev[6] = 11'b00000010101;
        h_t_prev[7] = 11'b00000011010;
        h_t_prev[8] = 11'b00000010000;
        h_t_prev[9] = 11'b00000001110;
        h_t_prev[10] = 11'b00000001110;
        h_t_prev[11] = 11'b00000010000;
        h_t_prev[12] = 11'b00000100100;
        h_t_prev[13] = 11'b00000100110;
        h_t_prev[14] = 11'b00000011000;
        h_t_prev[15] = 11'b00000010111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 21 timeout!");
                $fdisplay(fd_cycles, "Test Vector  21: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  21: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 21");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 22
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000000110;
        x_t[1] = 11'b00000001011;
        x_t[2] = 11'b11111111101;
        x_t[3] = 11'b00000000010;
        x_t[4] = 11'b00000001001;
        x_t[5] = 11'b00000001110;
        x_t[6] = 11'b00000010101;
        x_t[7] = 11'b00000010110;
        x_t[8] = 11'b00000000111;
        x_t[9] = 11'b00000001000;
        x_t[10] = 11'b00000001011;
        x_t[11] = 11'b00000010000;
        x_t[12] = 11'b00000011111;
        x_t[13] = 11'b00000100111;
        x_t[14] = 11'b00000010110;
        x_t[15] = 11'b00000010011;
        x_t[16] = 11'b00000001110;
        x_t[17] = 11'b00000010101;
        x_t[18] = 11'b00000011001;
        x_t[19] = 11'b00000100100;
        x_t[20] = 11'b00000110001;
        x_t[21] = 11'b00000000011;
        x_t[22] = 11'b00000001010;
        x_t[23] = 11'b00000001110;
        x_t[24] = 11'b00000001101;
        x_t[25] = 11'b00000001011;
        x_t[26] = 11'b11111111110;
        x_t[27] = 11'b00000000100;
        x_t[28] = 11'b00000010001;
        x_t[29] = 11'b00000010000;
        x_t[30] = 11'b00000011111;
        x_t[31] = 11'b00000001110;
        x_t[32] = 11'b00000000101;
        x_t[33] = 11'b00000000100;
        x_t[34] = 11'b00000000011;
        x_t[35] = 11'b00000000000;
        x_t[36] = 11'b00000001101;
        x_t[37] = 11'b11111010100;
        x_t[38] = 11'b00000100001;
        x_t[39] = 11'b00000010000;
        x_t[40] = 11'b00000011100;
        x_t[41] = 11'b00000010000;
        x_t[42] = 11'b00000101111;
        x_t[43] = 11'b11111111110;
        x_t[44] = 11'b00000011110;
        x_t[45] = 11'b00000100011;
        x_t[46] = 11'b00000100100;
        x_t[47] = 11'b00000100100;
        x_t[48] = 11'b00000011111;
        x_t[49] = 11'b00000011111;
        x_t[50] = 11'b00000100010;
        x_t[51] = 11'b00000101111;
        x_t[52] = 11'b00000110000;
        x_t[53] = 11'b00000101101;
        x_t[54] = 11'b00000100111;
        x_t[55] = 11'b00000100101;
        x_t[56] = 11'b00000100111;
        x_t[57] = 11'b00000101011;
        x_t[58] = 11'b00000111010;
        x_t[59] = 11'b00000101110;
        x_t[60] = 11'b00000010001;
        x_t[61] = 11'b00000101100;
        x_t[62] = 11'b00000110010;
        x_t[63] = 11'b00000011010;
        
        h_t_prev[0] = 11'b00000000110;
        h_t_prev[1] = 11'b00000001011;
        h_t_prev[2] = 11'b11111111101;
        h_t_prev[3] = 11'b00000000010;
        h_t_prev[4] = 11'b00000001001;
        h_t_prev[5] = 11'b00000001110;
        h_t_prev[6] = 11'b00000010101;
        h_t_prev[7] = 11'b00000010110;
        h_t_prev[8] = 11'b00000000111;
        h_t_prev[9] = 11'b00000001000;
        h_t_prev[10] = 11'b00000001011;
        h_t_prev[11] = 11'b00000010000;
        h_t_prev[12] = 11'b00000011111;
        h_t_prev[13] = 11'b00000100111;
        h_t_prev[14] = 11'b00000010110;
        h_t_prev[15] = 11'b00000010011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 22 timeout!");
                $fdisplay(fd_cycles, "Test Vector  22: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  22: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 22");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 23
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000100110;
        x_t[1] = 11'b00000100001;
        x_t[2] = 11'b00000001011;
        x_t[3] = 11'b00000010001;
        x_t[4] = 11'b00000001101;
        x_t[5] = 11'b00000001110;
        x_t[6] = 11'b00000010100;
        x_t[7] = 11'b00000110110;
        x_t[8] = 11'b00000011101;
        x_t[9] = 11'b00000010110;
        x_t[10] = 11'b00000010101;
        x_t[11] = 11'b00000010011;
        x_t[12] = 11'b00000011001;
        x_t[13] = 11'b00000011100;
        x_t[14] = 11'b00000110001;
        x_t[15] = 11'b00000100100;
        x_t[16] = 11'b00000011100;
        x_t[17] = 11'b00000011101;
        x_t[18] = 11'b00000011011;
        x_t[19] = 11'b00000100010;
        x_t[20] = 11'b00000101001;
        x_t[21] = 11'b00000001110;
        x_t[22] = 11'b00000010101;
        x_t[23] = 11'b00000010111;
        x_t[24] = 11'b00000010111;
        x_t[25] = 11'b00000010111;
        x_t[26] = 11'b00000000011;
        x_t[27] = 11'b00000001010;
        x_t[28] = 11'b00000011110;
        x_t[29] = 11'b00000011010;
        x_t[30] = 11'b00000100111;
        x_t[31] = 11'b00000001100;
        x_t[32] = 11'b00000001001;
        x_t[33] = 11'b00000000110;
        x_t[34] = 11'b00000000011;
        x_t[35] = 11'b11111111111;
        x_t[36] = 11'b00000001100;
        x_t[37] = 11'b11111011111;
        x_t[38] = 11'b00000100001;
        x_t[39] = 11'b00000010010;
        x_t[40] = 11'b00000100111;
        x_t[41] = 11'b00000000110;
        x_t[42] = 11'b00000101110;
        x_t[43] = 11'b00000001100;
        x_t[44] = 11'b00000110110;
        x_t[45] = 11'b00000011010;
        x_t[46] = 11'b00000110100;
        x_t[47] = 11'b00000101011;
        x_t[48] = 11'b00000100010;
        x_t[49] = 11'b00000011111;
        x_t[50] = 11'b00000011111;
        x_t[51] = 11'b00000101001;
        x_t[52] = 11'b00000100111;
        x_t[53] = 11'b00000100101;
        x_t[54] = 11'b00000100101;
        x_t[55] = 11'b00000100111;
        x_t[56] = 11'b00000100101;
        x_t[57] = 11'b00000100101;
        x_t[58] = 11'b00000110100;
        x_t[59] = 11'b00000101100;
        x_t[60] = 11'b00000011011;
        x_t[61] = 11'b00000110011;
        x_t[62] = 11'b00000110010;
        x_t[63] = 11'b00000101010;
        
        h_t_prev[0] = 11'b00000100110;
        h_t_prev[1] = 11'b00000100001;
        h_t_prev[2] = 11'b00000001011;
        h_t_prev[3] = 11'b00000010001;
        h_t_prev[4] = 11'b00000001101;
        h_t_prev[5] = 11'b00000001110;
        h_t_prev[6] = 11'b00000010100;
        h_t_prev[7] = 11'b00000110110;
        h_t_prev[8] = 11'b00000011101;
        h_t_prev[9] = 11'b00000010110;
        h_t_prev[10] = 11'b00000010101;
        h_t_prev[11] = 11'b00000010011;
        h_t_prev[12] = 11'b00000011001;
        h_t_prev[13] = 11'b00000011100;
        h_t_prev[14] = 11'b00000110001;
        h_t_prev[15] = 11'b00000100100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 23 timeout!");
                $fdisplay(fd_cycles, "Test Vector  23: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  23: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 23");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 24
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000001001;
        x_t[1] = 11'b00000001110;
        x_t[2] = 11'b11111111111;
        x_t[3] = 11'b00000000111;
        x_t[4] = 11'b11111111111;
        x_t[5] = 11'b11111111100;
        x_t[6] = 11'b00000000011;
        x_t[7] = 11'b00000011010;
        x_t[8] = 11'b00000001011;
        x_t[9] = 11'b00000001100;
        x_t[10] = 11'b00000001100;
        x_t[11] = 11'b00000000001;
        x_t[12] = 11'b00000001000;
        x_t[13] = 11'b00000000011;
        x_t[14] = 11'b00000100100;
        x_t[15] = 11'b00000011000;
        x_t[16] = 11'b00000010010;
        x_t[17] = 11'b00000010101;
        x_t[18] = 11'b00000001111;
        x_t[19] = 11'b00000010101;
        x_t[20] = 11'b00000011000;
        x_t[21] = 11'b11111110101;
        x_t[22] = 11'b11111111110;
        x_t[23] = 11'b00000000101;
        x_t[24] = 11'b11111111010;
        x_t[25] = 11'b11111111010;
        x_t[26] = 11'b11111101111;
        x_t[27] = 11'b11111110101;
        x_t[28] = 11'b00000001010;
        x_t[29] = 11'b11111111000;
        x_t[30] = 11'b00000001101;
        x_t[31] = 11'b11111111100;
        x_t[32] = 11'b11111111010;
        x_t[33] = 11'b11111110110;
        x_t[34] = 11'b11111110010;
        x_t[35] = 11'b11111101011;
        x_t[36] = 11'b11111110100;
        x_t[37] = 11'b11111010101;
        x_t[38] = 11'b11111111111;
        x_t[39] = 11'b11111111011;
        x_t[40] = 11'b00000101010;
        x_t[41] = 11'b11111011101;
        x_t[42] = 11'b00000101001;
        x_t[43] = 11'b00000010001;
        x_t[44] = 11'b00000110110;
        x_t[45] = 11'b00000100100;
        x_t[46] = 11'b00000110001;
        x_t[47] = 11'b00000100111;
        x_t[48] = 11'b00000100001;
        x_t[49] = 11'b00000011110;
        x_t[50] = 11'b00000011100;
        x_t[51] = 11'b00000101000;
        x_t[52] = 11'b00000100111;
        x_t[53] = 11'b00000100110;
        x_t[54] = 11'b00000101101;
        x_t[55] = 11'b00000011111;
        x_t[56] = 11'b00000100001;
        x_t[57] = 11'b00000100011;
        x_t[58] = 11'b00000110110;
        x_t[59] = 11'b00000110011;
        x_t[60] = 11'b00000011011;
        x_t[61] = 11'b00000110011;
        x_t[62] = 11'b00000110000;
        x_t[63] = 11'b00000101001;
        
        h_t_prev[0] = 11'b00000001001;
        h_t_prev[1] = 11'b00000001110;
        h_t_prev[2] = 11'b11111111111;
        h_t_prev[3] = 11'b00000000111;
        h_t_prev[4] = 11'b11111111111;
        h_t_prev[5] = 11'b11111111100;
        h_t_prev[6] = 11'b00000000011;
        h_t_prev[7] = 11'b00000011010;
        h_t_prev[8] = 11'b00000001011;
        h_t_prev[9] = 11'b00000001100;
        h_t_prev[10] = 11'b00000001100;
        h_t_prev[11] = 11'b00000000001;
        h_t_prev[12] = 11'b00000001000;
        h_t_prev[13] = 11'b00000000011;
        h_t_prev[14] = 11'b00000100100;
        h_t_prev[15] = 11'b00000011000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 24 timeout!");
                $fdisplay(fd_cycles, "Test Vector  24: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  24: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 24");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 25
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000001001;
        x_t[1] = 11'b00000010010;
        x_t[2] = 11'b00000000100;
        x_t[3] = 11'b00000001010;
        x_t[4] = 11'b00000000000;
        x_t[5] = 11'b11111111001;
        x_t[6] = 11'b11111110101;
        x_t[7] = 11'b00000101010;
        x_t[8] = 11'b00000010110;
        x_t[9] = 11'b00000010110;
        x_t[10] = 11'b00000010100;
        x_t[11] = 11'b00000001010;
        x_t[12] = 11'b00000001011;
        x_t[13] = 11'b11111111111;
        x_t[14] = 11'b00000110001;
        x_t[15] = 11'b00000100111;
        x_t[16] = 11'b00000011100;
        x_t[17] = 11'b00000011111;
        x_t[18] = 11'b00000010110;
        x_t[19] = 11'b00000011001;
        x_t[20] = 11'b00000011101;
        x_t[21] = 11'b11111111110;
        x_t[22] = 11'b00000000001;
        x_t[23] = 11'b00000000101;
        x_t[24] = 11'b00000000111;
        x_t[25] = 11'b00000000101;
        x_t[26] = 11'b11111110111;
        x_t[27] = 11'b11111110110;
        x_t[28] = 11'b00000000100;
        x_t[29] = 11'b00000000000;
        x_t[30] = 11'b00000011000;
        x_t[31] = 11'b00000000100;
        x_t[32] = 11'b00000001000;
        x_t[33] = 11'b00000000100;
        x_t[34] = 11'b11111111011;
        x_t[35] = 11'b11111110111;
        x_t[36] = 11'b11111110111;
        x_t[37] = 11'b11111010100;
        x_t[38] = 11'b00000001011;
        x_t[39] = 11'b11111110111;
        x_t[40] = 11'b00000010011;
        x_t[41] = 11'b11111100100;
        x_t[42] = 11'b00000011110;
        x_t[43] = 11'b00000010100;
        x_t[44] = 11'b00000100011;
        x_t[45] = 11'b00000101001;
        x_t[46] = 11'b00000101011;
        x_t[47] = 11'b00000101011;
        x_t[48] = 11'b00000100111;
        x_t[49] = 11'b00000100101;
        x_t[50] = 11'b00000100100;
        x_t[51] = 11'b00000101010;
        x_t[52] = 11'b00000101001;
        x_t[53] = 11'b00000100111;
        x_t[54] = 11'b00000101010;
        x_t[55] = 11'b00000100011;
        x_t[56] = 11'b00000100011;
        x_t[57] = 11'b00000100011;
        x_t[58] = 11'b00000110100;
        x_t[59] = 11'b00000101110;
        x_t[60] = 11'b00000011001;
        x_t[61] = 11'b00000110000;
        x_t[62] = 11'b00000101100;
        x_t[63] = 11'b00000100011;
        
        h_t_prev[0] = 11'b00000001001;
        h_t_prev[1] = 11'b00000010010;
        h_t_prev[2] = 11'b00000000100;
        h_t_prev[3] = 11'b00000001010;
        h_t_prev[4] = 11'b00000000000;
        h_t_prev[5] = 11'b11111111001;
        h_t_prev[6] = 11'b11111110101;
        h_t_prev[7] = 11'b00000101010;
        h_t_prev[8] = 11'b00000010110;
        h_t_prev[9] = 11'b00000010110;
        h_t_prev[10] = 11'b00000010100;
        h_t_prev[11] = 11'b00000001010;
        h_t_prev[12] = 11'b00000001011;
        h_t_prev[13] = 11'b11111111111;
        h_t_prev[14] = 11'b00000110001;
        h_t_prev[15] = 11'b00000100111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 25 timeout!");
                $fdisplay(fd_cycles, "Test Vector  25: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  25: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 25");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 26
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000001010;
        x_t[1] = 11'b00000011001;
        x_t[2] = 11'b00000001110;
        x_t[3] = 11'b00000010110;
        x_t[4] = 11'b00000001010;
        x_t[5] = 11'b00000000110;
        x_t[6] = 11'b00000000011;
        x_t[7] = 11'b00000100001;
        x_t[8] = 11'b00000010111;
        x_t[9] = 11'b00000010111;
        x_t[10] = 11'b00000010101;
        x_t[11] = 11'b00000001111;
        x_t[12] = 11'b00000010001;
        x_t[13] = 11'b00000000110;
        x_t[14] = 11'b00000100000;
        x_t[15] = 11'b00000011011;
        x_t[16] = 11'b00000010110;
        x_t[17] = 11'b00000011100;
        x_t[18] = 11'b00000010100;
        x_t[19] = 11'b00000010110;
        x_t[20] = 11'b00000011010;
        x_t[21] = 11'b11111111000;
        x_t[22] = 11'b11111111111;
        x_t[23] = 11'b00000000100;
        x_t[24] = 11'b11111111100;
        x_t[25] = 11'b11111111101;
        x_t[26] = 11'b11111111100;
        x_t[27] = 11'b11111111010;
        x_t[28] = 11'b00000000110;
        x_t[29] = 11'b11111101011;
        x_t[30] = 11'b00000001100;
        x_t[31] = 11'b00000000011;
        x_t[32] = 11'b00000000110;
        x_t[33] = 11'b00000000100;
        x_t[34] = 11'b11111111101;
        x_t[35] = 11'b11111110101;
        x_t[36] = 11'b11111111011;
        x_t[37] = 11'b11111010111;
        x_t[38] = 11'b11111110101;
        x_t[39] = 11'b00000000001;
        x_t[40] = 11'b00000000001;
        x_t[41] = 11'b11111110110;
        x_t[42] = 11'b00000001100;
        x_t[43] = 11'b11111101111;
        x_t[44] = 11'b00000010010;
        x_t[45] = 11'b00000010101;
        x_t[46] = 11'b00000010010;
        x_t[47] = 11'b00000010010;
        x_t[48] = 11'b00000010101;
        x_t[49] = 11'b00000010001;
        x_t[50] = 11'b00000010101;
        x_t[51] = 11'b00000011010;
        x_t[52] = 11'b00000011001;
        x_t[53] = 11'b00000010111;
        x_t[54] = 11'b00000011001;
        x_t[55] = 11'b00000010000;
        x_t[56] = 11'b00000010010;
        x_t[57] = 11'b00000010010;
        x_t[58] = 11'b00000100100;
        x_t[59] = 11'b00000011111;
        x_t[60] = 11'b00000001111;
        x_t[61] = 11'b00000100011;
        x_t[62] = 11'b00000011101;
        x_t[63] = 11'b00000010000;
        
        h_t_prev[0] = 11'b00000001010;
        h_t_prev[1] = 11'b00000011001;
        h_t_prev[2] = 11'b00000001110;
        h_t_prev[3] = 11'b00000010110;
        h_t_prev[4] = 11'b00000001010;
        h_t_prev[5] = 11'b00000000110;
        h_t_prev[6] = 11'b00000000011;
        h_t_prev[7] = 11'b00000100001;
        h_t_prev[8] = 11'b00000010111;
        h_t_prev[9] = 11'b00000010111;
        h_t_prev[10] = 11'b00000010101;
        h_t_prev[11] = 11'b00000001111;
        h_t_prev[12] = 11'b00000010001;
        h_t_prev[13] = 11'b00000000110;
        h_t_prev[14] = 11'b00000100000;
        h_t_prev[15] = 11'b00000011011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 26 timeout!");
                $fdisplay(fd_cycles, "Test Vector  26: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  26: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 26");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 27
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111111010;
        x_t[1] = 11'b00000000110;
        x_t[2] = 11'b00000000001;
        x_t[3] = 11'b00000001001;
        x_t[4] = 11'b00000000000;
        x_t[5] = 11'b11111111110;
        x_t[6] = 11'b00000000001;
        x_t[7] = 11'b00000000101;
        x_t[8] = 11'b11111111111;
        x_t[9] = 11'b00000001000;
        x_t[10] = 11'b00000001001;
        x_t[11] = 11'b00000000001;
        x_t[12] = 11'b00000000110;
        x_t[13] = 11'b00000000011;
        x_t[14] = 11'b00000000101;
        x_t[15] = 11'b00000001001;
        x_t[16] = 11'b00000001000;
        x_t[17] = 11'b00000001111;
        x_t[18] = 11'b00000000110;
        x_t[19] = 11'b00000001001;
        x_t[20] = 11'b00000010011;
        x_t[21] = 11'b11111111110;
        x_t[22] = 11'b00000000100;
        x_t[23] = 11'b00000001010;
        x_t[24] = 11'b00000000001;
        x_t[25] = 11'b00000000001;
        x_t[26] = 11'b11111111011;
        x_t[27] = 11'b11111111101;
        x_t[28] = 11'b00000001100;
        x_t[29] = 11'b11111111011;
        x_t[30] = 11'b00000001100;
        x_t[31] = 11'b00000000010;
        x_t[32] = 11'b00000000000;
        x_t[33] = 11'b00000000000;
        x_t[34] = 11'b11111111001;
        x_t[35] = 11'b11111110010;
        x_t[36] = 11'b11111111111;
        x_t[37] = 11'b11111011111;
        x_t[38] = 11'b00000000100;
        x_t[39] = 11'b00000000111;
        x_t[40] = 11'b00000010101;
        x_t[41] = 11'b11111101111;
        x_t[42] = 11'b00000010010;
        x_t[43] = 11'b11111110101;
        x_t[44] = 11'b00000010001;
        x_t[45] = 11'b00000100100;
        x_t[46] = 11'b00000010000;
        x_t[47] = 11'b00000010000;
        x_t[48] = 11'b00000010101;
        x_t[49] = 11'b00000010000;
        x_t[50] = 11'b00000001111;
        x_t[51] = 11'b00000010011;
        x_t[52] = 11'b00000010010;
        x_t[53] = 11'b00000010010;
        x_t[54] = 11'b00000011110;
        x_t[55] = 11'b00000010001;
        x_t[56] = 11'b00000010111;
        x_t[57] = 11'b00000010001;
        x_t[58] = 11'b00000011101;
        x_t[59] = 11'b00000011100;
        x_t[60] = 11'b00000001001;
        x_t[61] = 11'b00000011010;
        x_t[62] = 11'b00000010001;
        x_t[63] = 11'b00000001000;
        
        h_t_prev[0] = 11'b11111111010;
        h_t_prev[1] = 11'b00000000110;
        h_t_prev[2] = 11'b00000000001;
        h_t_prev[3] = 11'b00000001001;
        h_t_prev[4] = 11'b00000000000;
        h_t_prev[5] = 11'b11111111110;
        h_t_prev[6] = 11'b00000000001;
        h_t_prev[7] = 11'b00000000101;
        h_t_prev[8] = 11'b11111111111;
        h_t_prev[9] = 11'b00000001000;
        h_t_prev[10] = 11'b00000001001;
        h_t_prev[11] = 11'b00000000001;
        h_t_prev[12] = 11'b00000000110;
        h_t_prev[13] = 11'b00000000011;
        h_t_prev[14] = 11'b00000000101;
        h_t_prev[15] = 11'b00000001001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 27 timeout!");
                $fdisplay(fd_cycles, "Test Vector  27: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  27: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 27");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 28
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000001001;
        x_t[1] = 11'b00000001001;
        x_t[2] = 11'b11111111110;
        x_t[3] = 11'b00000000001;
        x_t[4] = 11'b11111111000;
        x_t[5] = 11'b11111110111;
        x_t[6] = 11'b11111111100;
        x_t[7] = 11'b00000011000;
        x_t[8] = 11'b00000000110;
        x_t[9] = 11'b00000001001;
        x_t[10] = 11'b00000001001;
        x_t[11] = 11'b11111111011;
        x_t[12] = 11'b11111111101;
        x_t[13] = 11'b11111111001;
        x_t[14] = 11'b00000010011;
        x_t[15] = 11'b00000010001;
        x_t[16] = 11'b00000001100;
        x_t[17] = 11'b00000001111;
        x_t[18] = 11'b00000000000;
        x_t[19] = 11'b11111111111;
        x_t[20] = 11'b00000001010;
        x_t[21] = 11'b00000000101;
        x_t[22] = 11'b00000001010;
        x_t[23] = 11'b00000001110;
        x_t[24] = 11'b00000001011;
        x_t[25] = 11'b00000001011;
        x_t[26] = 11'b11111110111;
        x_t[27] = 11'b11111111010;
        x_t[28] = 11'b00000001000;
        x_t[29] = 11'b00000000010;
        x_t[30] = 11'b00000010101;
        x_t[31] = 11'b11111111010;
        x_t[32] = 11'b11111111010;
        x_t[33] = 11'b11111111001;
        x_t[34] = 11'b11111110010;
        x_t[35] = 11'b11111101100;
        x_t[36] = 11'b11111110110;
        x_t[37] = 11'b11111011100;
        x_t[38] = 11'b00000010000;
        x_t[39] = 11'b11111110110;
        x_t[40] = 11'b00000011010;
        x_t[41] = 11'b11111100100;
        x_t[42] = 11'b00000001111;
        x_t[43] = 11'b00000011000;
        x_t[44] = 11'b00000010110;
        x_t[45] = 11'b00000010000;
        x_t[46] = 11'b00000010110;
        x_t[47] = 11'b00000010100;
        x_t[48] = 11'b00000010101;
        x_t[49] = 11'b00000001111;
        x_t[50] = 11'b00000000101;
        x_t[51] = 11'b00000000011;
        x_t[52] = 11'b11111111110;
        x_t[53] = 11'b11111111101;
        x_t[54] = 11'b00000001010;
        x_t[55] = 11'b00000010110;
        x_t[56] = 11'b00000011001;
        x_t[57] = 11'b00000001001;
        x_t[58] = 11'b00000001001;
        x_t[59] = 11'b00000001000;
        x_t[60] = 11'b00000001010;
        x_t[61] = 11'b00000010110;
        x_t[62] = 11'b00000001010;
        x_t[63] = 11'b00000001001;
        
        h_t_prev[0] = 11'b00000001001;
        h_t_prev[1] = 11'b00000001001;
        h_t_prev[2] = 11'b11111111110;
        h_t_prev[3] = 11'b00000000001;
        h_t_prev[4] = 11'b11111111000;
        h_t_prev[5] = 11'b11111110111;
        h_t_prev[6] = 11'b11111111100;
        h_t_prev[7] = 11'b00000011000;
        h_t_prev[8] = 11'b00000000110;
        h_t_prev[9] = 11'b00000001001;
        h_t_prev[10] = 11'b00000001001;
        h_t_prev[11] = 11'b11111111011;
        h_t_prev[12] = 11'b11111111101;
        h_t_prev[13] = 11'b11111111001;
        h_t_prev[14] = 11'b00000010011;
        h_t_prev[15] = 11'b00000010001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 28 timeout!");
                $fdisplay(fd_cycles, "Test Vector  28: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  28: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 28");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 29
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000001010;
        x_t[1] = 11'b00000001010;
        x_t[2] = 11'b11111111011;
        x_t[3] = 11'b11111111101;
        x_t[4] = 11'b11111110000;
        x_t[5] = 11'b11111101001;
        x_t[6] = 11'b11111110000;
        x_t[7] = 11'b00000011011;
        x_t[8] = 11'b00000001101;
        x_t[9] = 11'b00000001000;
        x_t[10] = 11'b00000000011;
        x_t[11] = 11'b11111111010;
        x_t[12] = 11'b11111110000;
        x_t[13] = 11'b11111101010;
        x_t[14] = 11'b00000010110;
        x_t[15] = 11'b00000010000;
        x_t[16] = 11'b00000001011;
        x_t[17] = 11'b00000001010;
        x_t[18] = 11'b11111110111;
        x_t[19] = 11'b11111110010;
        x_t[20] = 11'b11111111001;
        x_t[21] = 11'b00000000001;
        x_t[22] = 11'b00000000111;
        x_t[23] = 11'b00000001001;
        x_t[24] = 11'b00000001001;
        x_t[25] = 11'b00000001001;
        x_t[26] = 11'b11111111010;
        x_t[27] = 11'b11111111000;
        x_t[28] = 11'b00000000011;
        x_t[29] = 11'b00000000111;
        x_t[30] = 11'b00000010011;
        x_t[31] = 11'b11111111111;
        x_t[32] = 11'b11111111111;
        x_t[33] = 11'b00000000000;
        x_t[34] = 11'b11111110111;
        x_t[35] = 11'b11111101111;
        x_t[36] = 11'b11111111000;
        x_t[37] = 11'b11111011100;
        x_t[38] = 11'b00000010011;
        x_t[39] = 11'b11111110111;
        x_t[40] = 11'b00000011101;
        x_t[41] = 11'b00000000101;
        x_t[42] = 11'b00000101100;
        x_t[43] = 11'b11111111010;
        x_t[44] = 11'b00000100101;
        x_t[45] = 11'b00000000100;
        x_t[46] = 11'b00000100010;
        x_t[47] = 11'b00000011011;
        x_t[48] = 11'b00000011010;
        x_t[49] = 11'b00000010011;
        x_t[50] = 11'b00000001010;
        x_t[51] = 11'b00000000000;
        x_t[52] = 11'b11111111100;
        x_t[53] = 11'b11111110111;
        x_t[54] = 11'b00000000001;
        x_t[55] = 11'b00000100001;
        x_t[56] = 11'b00000100001;
        x_t[57] = 11'b00000001010;
        x_t[58] = 11'b11111111110;
        x_t[59] = 11'b00000000000;
        x_t[60] = 11'b00000010010;
        x_t[61] = 11'b00000010110;
        x_t[62] = 11'b00000000001;
        x_t[63] = 11'b00000001100;
        
        h_t_prev[0] = 11'b00000001010;
        h_t_prev[1] = 11'b00000001010;
        h_t_prev[2] = 11'b11111111011;
        h_t_prev[3] = 11'b11111111101;
        h_t_prev[4] = 11'b11111110000;
        h_t_prev[5] = 11'b11111101001;
        h_t_prev[6] = 11'b11111110000;
        h_t_prev[7] = 11'b00000011011;
        h_t_prev[8] = 11'b00000001101;
        h_t_prev[9] = 11'b00000001000;
        h_t_prev[10] = 11'b00000000011;
        h_t_prev[11] = 11'b11111111010;
        h_t_prev[12] = 11'b11111110000;
        h_t_prev[13] = 11'b11111101010;
        h_t_prev[14] = 11'b00000010110;
        h_t_prev[15] = 11'b00000010000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 29 timeout!");
                $fdisplay(fd_cycles, "Test Vector  29: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  29: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 29");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 30
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000011000;
        x_t[1] = 11'b00000011100;
        x_t[2] = 11'b00000001101;
        x_t[3] = 11'b00000001111;
        x_t[4] = 11'b00000000111;
        x_t[5] = 11'b11111111101;
        x_t[6] = 11'b00000000110;
        x_t[7] = 11'b00000101101;
        x_t[8] = 11'b00000011101;
        x_t[9] = 11'b00000011001;
        x_t[10] = 11'b00000010101;
        x_t[11] = 11'b00000001001;
        x_t[12] = 11'b00000000000;
        x_t[13] = 11'b00000000111;
        x_t[14] = 11'b00000100001;
        x_t[15] = 11'b00000011100;
        x_t[16] = 11'b00000010110;
        x_t[17] = 11'b00000010111;
        x_t[18] = 11'b00000000100;
        x_t[19] = 11'b11111111010;
        x_t[20] = 11'b00000000010;
        x_t[21] = 11'b00000010011;
        x_t[22] = 11'b00000011001;
        x_t[23] = 11'b00000011000;
        x_t[24] = 11'b00000011100;
        x_t[25] = 11'b00000011100;
        x_t[26] = 11'b00000001110;
        x_t[27] = 11'b00000001011;
        x_t[28] = 11'b00000010100;
        x_t[29] = 11'b00000011110;
        x_t[30] = 11'b00000100011;
        x_t[31] = 11'b00000010001;
        x_t[32] = 11'b00000010010;
        x_t[33] = 11'b00000010100;
        x_t[34] = 11'b00000001100;
        x_t[35] = 11'b00000000011;
        x_t[36] = 11'b00000001010;
        x_t[37] = 11'b11111101011;
        x_t[38] = 11'b00000100100;
        x_t[39] = 11'b00000010001;
        x_t[40] = 11'b00000100101;
        x_t[41] = 11'b00000010001;
        x_t[42] = 11'b00000111101;
        x_t[43] = 11'b11111110101;
        x_t[44] = 11'b00000101111;
        x_t[45] = 11'b11111111011;
        x_t[46] = 11'b00000101100;
        x_t[47] = 11'b00000011111;
        x_t[48] = 11'b00000011011;
        x_t[49] = 11'b00000010010;
        x_t[50] = 11'b00000000100;
        x_t[51] = 11'b11111101110;
        x_t[52] = 11'b11111101010;
        x_t[53] = 11'b11111100001;
        x_t[54] = 11'b11111101100;
        x_t[55] = 11'b00000100100;
        x_t[56] = 11'b00000100000;
        x_t[57] = 11'b11111111011;
        x_t[58] = 11'b11111011011;
        x_t[59] = 11'b11111100110;
        x_t[60] = 11'b00000011000;
        x_t[61] = 11'b00000010010;
        x_t[62] = 11'b11111110000;
        x_t[63] = 11'b00000001101;
        
        h_t_prev[0] = 11'b00000011000;
        h_t_prev[1] = 11'b00000011100;
        h_t_prev[2] = 11'b00000001101;
        h_t_prev[3] = 11'b00000001111;
        h_t_prev[4] = 11'b00000000111;
        h_t_prev[5] = 11'b11111111101;
        h_t_prev[6] = 11'b00000000110;
        h_t_prev[7] = 11'b00000101101;
        h_t_prev[8] = 11'b00000011101;
        h_t_prev[9] = 11'b00000011001;
        h_t_prev[10] = 11'b00000010101;
        h_t_prev[11] = 11'b00000001001;
        h_t_prev[12] = 11'b00000000000;
        h_t_prev[13] = 11'b00000000111;
        h_t_prev[14] = 11'b00000100001;
        h_t_prev[15] = 11'b00000011100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 30 timeout!");
                $fdisplay(fd_cycles, "Test Vector  30: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  30: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 30");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 31
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000011111;
        x_t[1] = 11'b00000100000;
        x_t[2] = 11'b00000001110;
        x_t[3] = 11'b00000010111;
        x_t[4] = 11'b00000001011;
        x_t[5] = 11'b00000000000;
        x_t[6] = 11'b00000000000;
        x_t[7] = 11'b00000101001;
        x_t[8] = 11'b00000011001;
        x_t[9] = 11'b00000010110;
        x_t[10] = 11'b00000010010;
        x_t[11] = 11'b11111111111;
        x_t[12] = 11'b11111110111;
        x_t[13] = 11'b11111110010;
        x_t[14] = 11'b00000011110;
        x_t[15] = 11'b00000010011;
        x_t[16] = 11'b00000001100;
        x_t[17] = 11'b00000001001;
        x_t[18] = 11'b11111110101;
        x_t[19] = 11'b11111101000;
        x_t[20] = 11'b11111101001;
        x_t[21] = 11'b00000010100;
        x_t[22] = 11'b00000011010;
        x_t[23] = 11'b00000011011;
        x_t[24] = 11'b00000010111;
        x_t[25] = 11'b00000011000;
        x_t[26] = 11'b00000001100;
        x_t[27] = 11'b00000001010;
        x_t[28] = 11'b00000010011;
        x_t[29] = 11'b00000010111;
        x_t[30] = 11'b00000011001;
        x_t[31] = 11'b00000001010;
        x_t[32] = 11'b00000001101;
        x_t[33] = 11'b00000001110;
        x_t[34] = 11'b00000001000;
        x_t[35] = 11'b11111111110;
        x_t[36] = 11'b00000000100;
        x_t[37] = 11'b11111100010;
        x_t[38] = 11'b00000010100;
        x_t[39] = 11'b11111111111;
        x_t[40] = 11'b00000100010;
        x_t[41] = 11'b11111011000;
        x_t[42] = 11'b00000101001;
        x_t[43] = 11'b00000010100;
        x_t[44] = 11'b00000101010;
        x_t[45] = 11'b11111101011;
        x_t[46] = 11'b00000101000;
        x_t[47] = 11'b00000010010;
        x_t[48] = 11'b00000001000;
        x_t[49] = 11'b00000000001;
        x_t[50] = 11'b11111101111;
        x_t[51] = 11'b11111010101;
        x_t[52] = 11'b11111010000;
        x_t[53] = 11'b11111001100;
        x_t[54] = 11'b11111011111;
        x_t[55] = 11'b00000011011;
        x_t[56] = 11'b00000010101;
        x_t[57] = 11'b11111101010;
        x_t[58] = 11'b11111000011;
        x_t[59] = 11'b11111011000;
        x_t[60] = 11'b00000010101;
        x_t[61] = 11'b00000000101;
        x_t[62] = 11'b11111011010;
        x_t[63] = 11'b00000001101;
        
        h_t_prev[0] = 11'b00000011111;
        h_t_prev[1] = 11'b00000100000;
        h_t_prev[2] = 11'b00000001110;
        h_t_prev[3] = 11'b00000010111;
        h_t_prev[4] = 11'b00000001011;
        h_t_prev[5] = 11'b00000000000;
        h_t_prev[6] = 11'b00000000000;
        h_t_prev[7] = 11'b00000101001;
        h_t_prev[8] = 11'b00000011001;
        h_t_prev[9] = 11'b00000010110;
        h_t_prev[10] = 11'b00000010010;
        h_t_prev[11] = 11'b11111111111;
        h_t_prev[12] = 11'b11111110111;
        h_t_prev[13] = 11'b11111110010;
        h_t_prev[14] = 11'b00000011110;
        h_t_prev[15] = 11'b00000010011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 31 timeout!");
                $fdisplay(fd_cycles, "Test Vector  31: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  31: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 31");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 32
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000001100;
        x_t[1] = 11'b00000010101;
        x_t[2] = 11'b11111111110;
        x_t[3] = 11'b00000010010;
        x_t[4] = 11'b00000000110;
        x_t[5] = 11'b11111111000;
        x_t[6] = 11'b11111111011;
        x_t[7] = 11'b00000011101;
        x_t[8] = 11'b00000001110;
        x_t[9] = 11'b00000001101;
        x_t[10] = 11'b00000001001;
        x_t[11] = 11'b11111111011;
        x_t[12] = 11'b11111111000;
        x_t[13] = 11'b11111101101;
        x_t[14] = 11'b00000010110;
        x_t[15] = 11'b00000001011;
        x_t[16] = 11'b00000000010;
        x_t[17] = 11'b11111111111;
        x_t[18] = 11'b11111110001;
        x_t[19] = 11'b11111101100;
        x_t[20] = 11'b11111101111;
        x_t[21] = 11'b00000001000;
        x_t[22] = 11'b00000010000;
        x_t[23] = 11'b00000010011;
        x_t[24] = 11'b00000001110;
        x_t[25] = 11'b00000001110;
        x_t[26] = 11'b00000000101;
        x_t[27] = 11'b00000000010;
        x_t[28] = 11'b00000001101;
        x_t[29] = 11'b00000000101;
        x_t[30] = 11'b00000001111;
        x_t[31] = 11'b00000001000;
        x_t[32] = 11'b00000001010;
        x_t[33] = 11'b00000001110;
        x_t[34] = 11'b00000000101;
        x_t[35] = 11'b11111111000;
        x_t[36] = 11'b00000000011;
        x_t[37] = 11'b11111011100;
        x_t[38] = 11'b11111111111;
        x_t[39] = 11'b00000000110;
        x_t[40] = 11'b00000010011;
        x_t[41] = 11'b11111101100;
        x_t[42] = 11'b00000011010;
        x_t[43] = 11'b11111110000;
        x_t[44] = 11'b00000011000;
        x_t[45] = 11'b11111111101;
        x_t[46] = 11'b00000011000;
        x_t[47] = 11'b00000001101;
        x_t[48] = 11'b00000001000;
        x_t[49] = 11'b11111111010;
        x_t[50] = 11'b11111101110;
        x_t[51] = 11'b11111011011;
        x_t[52] = 11'b11111011001;
        x_t[53] = 11'b11111010101;
        x_t[54] = 11'b11111100011;
        x_t[55] = 11'b00000010110;
        x_t[56] = 11'b00000001111;
        x_t[57] = 11'b11111100101;
        x_t[58] = 11'b11111001001;
        x_t[59] = 11'b11111011001;
        x_t[60] = 11'b00000001111;
        x_t[61] = 11'b11111111000;
        x_t[62] = 11'b11111001110;
        x_t[63] = 11'b00000001011;
        
        h_t_prev[0] = 11'b00000001100;
        h_t_prev[1] = 11'b00000010101;
        h_t_prev[2] = 11'b11111111110;
        h_t_prev[3] = 11'b00000010010;
        h_t_prev[4] = 11'b00000000110;
        h_t_prev[5] = 11'b11111111000;
        h_t_prev[6] = 11'b11111111011;
        h_t_prev[7] = 11'b00000011101;
        h_t_prev[8] = 11'b00000001110;
        h_t_prev[9] = 11'b00000001101;
        h_t_prev[10] = 11'b00000001001;
        h_t_prev[11] = 11'b11111111011;
        h_t_prev[12] = 11'b11111111000;
        h_t_prev[13] = 11'b11111101101;
        h_t_prev[14] = 11'b00000010110;
        h_t_prev[15] = 11'b00000001011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 32 timeout!");
                $fdisplay(fd_cycles, "Test Vector  32: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  32: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 32");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 33
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111110101;
        x_t[1] = 11'b11111110101;
        x_t[2] = 11'b11111110000;
        x_t[3] = 11'b11111110001;
        x_t[4] = 11'b11111101100;
        x_t[5] = 11'b11111011100;
        x_t[6] = 11'b11111011000;
        x_t[7] = 11'b11111111101;
        x_t[8] = 11'b11111110001;
        x_t[9] = 11'b11111101101;
        x_t[10] = 11'b11111101100;
        x_t[11] = 11'b11111100101;
        x_t[12] = 11'b11111011101;
        x_t[13] = 11'b11111001000;
        x_t[14] = 11'b11111111101;
        x_t[15] = 11'b11111110011;
        x_t[16] = 11'b11111101110;
        x_t[17] = 11'b11111101001;
        x_t[18] = 11'b11111101001;
        x_t[19] = 11'b11111100101;
        x_t[20] = 11'b11111100001;
        x_t[21] = 11'b11111110110;
        x_t[22] = 11'b11111101010;
        x_t[23] = 11'b11111110001;
        x_t[24] = 11'b11111110101;
        x_t[25] = 11'b11111110110;
        x_t[26] = 11'b11111100110;
        x_t[27] = 11'b11111101010;
        x_t[28] = 11'b11111101010;
        x_t[29] = 11'b11111110111;
        x_t[30] = 11'b11111101001;
        x_t[31] = 11'b11111110110;
        x_t[32] = 11'b11111110001;
        x_t[33] = 11'b11111101001;
        x_t[34] = 11'b11111100011;
        x_t[35] = 11'b11111011110;
        x_t[36] = 11'b11111011100;
        x_t[37] = 11'b11111000011;
        x_t[38] = 11'b11111110001;
        x_t[39] = 11'b11111000111;
        x_t[40] = 11'b11111110000;
        x_t[41] = 11'b11111010101;
        x_t[42] = 11'b11111111100;
        x_t[43] = 11'b11111110110;
        x_t[44] = 11'b11111011100;
        x_t[45] = 11'b11111011000;
        x_t[46] = 11'b11111111110;
        x_t[47] = 11'b11111111000;
        x_t[48] = 11'b11111110011;
        x_t[49] = 11'b11111111010;
        x_t[50] = 11'b11111110001;
        x_t[51] = 11'b11111110010;
        x_t[52] = 11'b11111110010;
        x_t[53] = 11'b11111101000;
        x_t[54] = 11'b11111100100;
        x_t[55] = 11'b11111111000;
        x_t[56] = 11'b11111111110;
        x_t[57] = 11'b11111111110;
        x_t[58] = 11'b00000000010;
        x_t[59] = 11'b00000000001;
        x_t[60] = 11'b11111110110;
        x_t[61] = 11'b11111101110;
        x_t[62] = 11'b11111110100;
        x_t[63] = 11'b11111100001;
        
        h_t_prev[0] = 11'b11111110101;
        h_t_prev[1] = 11'b11111110101;
        h_t_prev[2] = 11'b11111110000;
        h_t_prev[3] = 11'b11111110001;
        h_t_prev[4] = 11'b11111101100;
        h_t_prev[5] = 11'b11111011100;
        h_t_prev[6] = 11'b11111011000;
        h_t_prev[7] = 11'b11111111101;
        h_t_prev[8] = 11'b11111110001;
        h_t_prev[9] = 11'b11111101101;
        h_t_prev[10] = 11'b11111101100;
        h_t_prev[11] = 11'b11111100101;
        h_t_prev[12] = 11'b11111011101;
        h_t_prev[13] = 11'b11111001000;
        h_t_prev[14] = 11'b11111111101;
        h_t_prev[15] = 11'b11111110011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 33 timeout!");
                $fdisplay(fd_cycles, "Test Vector  33: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  33: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 33");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 34
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111100100;
        x_t[1] = 11'b11111100100;
        x_t[2] = 11'b11111011111;
        x_t[3] = 11'b11111011101;
        x_t[4] = 11'b11111011011;
        x_t[5] = 11'b11111001111;
        x_t[6] = 11'b11111001111;
        x_t[7] = 11'b11111110101;
        x_t[8] = 11'b11111101000;
        x_t[9] = 11'b11111100010;
        x_t[10] = 11'b11111100010;
        x_t[11] = 11'b11111100000;
        x_t[12] = 11'b11111011110;
        x_t[13] = 11'b11111010001;
        x_t[14] = 11'b11111110110;
        x_t[15] = 11'b11111101110;
        x_t[16] = 11'b11111101001;
        x_t[17] = 11'b11111100101;
        x_t[18] = 11'b11111101010;
        x_t[19] = 11'b11111101101;
        x_t[20] = 11'b11111101010;
        x_t[21] = 11'b11111101010;
        x_t[22] = 11'b11111011111;
        x_t[23] = 11'b11111100110;
        x_t[24] = 11'b11111101011;
        x_t[25] = 11'b11111101011;
        x_t[26] = 11'b11111010110;
        x_t[27] = 11'b11111011011;
        x_t[28] = 11'b11111011110;
        x_t[29] = 11'b11111101000;
        x_t[30] = 11'b11111011010;
        x_t[31] = 11'b11111101000;
        x_t[32] = 11'b11111100000;
        x_t[33] = 11'b11111011000;
        x_t[34] = 11'b11111010011;
        x_t[35] = 11'b11111001101;
        x_t[36] = 11'b11111001111;
        x_t[37] = 11'b11111000100;
        x_t[38] = 11'b11111100011;
        x_t[39] = 11'b11111001100;
        x_t[40] = 11'b11111100100;
        x_t[41] = 11'b11111100110;
        x_t[42] = 11'b11111100001;
        x_t[43] = 11'b11111001010;
        x_t[44] = 11'b11111001111;
        x_t[45] = 11'b11111101001;
        x_t[46] = 11'b11111110010;
        x_t[47] = 11'b11111111000;
        x_t[48] = 11'b11111111001;
        x_t[49] = 11'b00000000100;
        x_t[50] = 11'b11111111001;
        x_t[51] = 11'b11111111111;
        x_t[52] = 11'b00000000000;
        x_t[53] = 11'b11111110111;
        x_t[54] = 11'b11111110101;
        x_t[55] = 11'b11111111110;
        x_t[56] = 11'b00000000110;
        x_t[57] = 11'b00000001011;
        x_t[58] = 11'b00000001111;
        x_t[59] = 11'b00000010000;
        x_t[60] = 11'b11111111010;
        x_t[61] = 11'b11111110111;
        x_t[62] = 11'b00000000001;
        x_t[63] = 11'b11111101101;
        
        h_t_prev[0] = 11'b11111100100;
        h_t_prev[1] = 11'b11111100100;
        h_t_prev[2] = 11'b11111011111;
        h_t_prev[3] = 11'b11111011101;
        h_t_prev[4] = 11'b11111011011;
        h_t_prev[5] = 11'b11111001111;
        h_t_prev[6] = 11'b11111001111;
        h_t_prev[7] = 11'b11111110101;
        h_t_prev[8] = 11'b11111101000;
        h_t_prev[9] = 11'b11111100010;
        h_t_prev[10] = 11'b11111100010;
        h_t_prev[11] = 11'b11111100000;
        h_t_prev[12] = 11'b11111011110;
        h_t_prev[13] = 11'b11111010001;
        h_t_prev[14] = 11'b11111110110;
        h_t_prev[15] = 11'b11111101110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 34 timeout!");
                $fdisplay(fd_cycles, "Test Vector  34: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  34: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 34");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 35
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111100010;
        x_t[1] = 11'b11111100001;
        x_t[2] = 11'b11111011011;
        x_t[3] = 11'b11111011101;
        x_t[4] = 11'b11111011011;
        x_t[5] = 11'b11111010011;
        x_t[6] = 11'b11111001110;
        x_t[7] = 11'b11111110001;
        x_t[8] = 11'b11111101000;
        x_t[9] = 11'b11111100111;
        x_t[10] = 11'b11111101101;
        x_t[11] = 11'b11111101111;
        x_t[12] = 11'b11111101010;
        x_t[13] = 11'b11111100010;
        x_t[14] = 11'b11111101110;
        x_t[15] = 11'b11111110001;
        x_t[16] = 11'b11111110001;
        x_t[17] = 11'b11111101111;
        x_t[18] = 11'b11111110101;
        x_t[19] = 11'b11111111010;
        x_t[20] = 11'b11111111000;
        x_t[21] = 11'b11111100111;
        x_t[22] = 11'b11111011011;
        x_t[23] = 11'b11111100011;
        x_t[24] = 11'b11111101000;
        x_t[25] = 11'b11111101001;
        x_t[26] = 11'b11111011000;
        x_t[27] = 11'b11111011011;
        x_t[28] = 11'b11111011001;
        x_t[29] = 11'b11111100111;
        x_t[30] = 11'b11111011010;
        x_t[31] = 11'b11111101111;
        x_t[32] = 11'b11111101000;
        x_t[33] = 11'b11111100010;
        x_t[34] = 11'b11111011100;
        x_t[35] = 11'b11111010110;
        x_t[36] = 11'b11111011000;
        x_t[37] = 11'b11111000110;
        x_t[38] = 11'b11111101010;
        x_t[39] = 11'b11111011011;
        x_t[40] = 11'b11111110011;
        x_t[41] = 11'b11111111110;
        x_t[42] = 11'b11111110101;
        x_t[43] = 11'b11110111011;
        x_t[44] = 11'b11111011011;
        x_t[45] = 11'b11111110001;
        x_t[46] = 11'b00000000000;
        x_t[47] = 11'b00000000101;
        x_t[48] = 11'b00000000111;
        x_t[49] = 11'b00000010101;
        x_t[50] = 11'b00000001001;
        x_t[51] = 11'b00000001011;
        x_t[52] = 11'b00000001010;
        x_t[53] = 11'b00000000011;
        x_t[54] = 11'b00000000100;
        x_t[55] = 11'b00000001111;
        x_t[56] = 11'b00000011000;
        x_t[57] = 11'b00000011011;
        x_t[58] = 11'b00000010111;
        x_t[59] = 11'b00000011100;
        x_t[60] = 11'b00000001010;
        x_t[61] = 11'b00000001000;
        x_t[62] = 11'b00000010001;
        x_t[63] = 11'b00000000011;
        
        h_t_prev[0] = 11'b11111100010;
        h_t_prev[1] = 11'b11111100001;
        h_t_prev[2] = 11'b11111011011;
        h_t_prev[3] = 11'b11111011101;
        h_t_prev[4] = 11'b11111011011;
        h_t_prev[5] = 11'b11111010011;
        h_t_prev[6] = 11'b11111001110;
        h_t_prev[7] = 11'b11111110001;
        h_t_prev[8] = 11'b11111101000;
        h_t_prev[9] = 11'b11111100111;
        h_t_prev[10] = 11'b11111101101;
        h_t_prev[11] = 11'b11111101111;
        h_t_prev[12] = 11'b11111101010;
        h_t_prev[13] = 11'b11111100010;
        h_t_prev[14] = 11'b11111101110;
        h_t_prev[15] = 11'b11111110001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 35 timeout!");
                $fdisplay(fd_cycles, "Test Vector  35: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  35: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 35");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 36
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111101101;
        x_t[1] = 11'b11111110101;
        x_t[2] = 11'b11111110011;
        x_t[3] = 11'b11111110100;
        x_t[4] = 11'b11111110011;
        x_t[5] = 11'b11111101100;
        x_t[6] = 11'b11111100111;
        x_t[7] = 11'b00000000101;
        x_t[8] = 11'b11111111110;
        x_t[9] = 11'b11111111110;
        x_t[10] = 11'b00000000100;
        x_t[11] = 11'b00000000110;
        x_t[12] = 11'b11111111111;
        x_t[13] = 11'b11111110011;
        x_t[14] = 11'b00000001000;
        x_t[15] = 11'b00000001000;
        x_t[16] = 11'b00000001000;
        x_t[17] = 11'b00000000101;
        x_t[18] = 11'b00000001010;
        x_t[19] = 11'b00000001100;
        x_t[20] = 11'b00000001001;
        x_t[21] = 11'b11111110011;
        x_t[22] = 11'b11111100111;
        x_t[23] = 11'b11111101100;
        x_t[24] = 11'b11111110011;
        x_t[25] = 11'b11111110100;
        x_t[26] = 11'b11111101100;
        x_t[27] = 11'b11111101101;
        x_t[28] = 11'b11111100110;
        x_t[29] = 11'b11111110010;
        x_t[30] = 11'b11111101000;
        x_t[31] = 11'b00000000010;
        x_t[32] = 11'b11111111111;
        x_t[33] = 11'b11111111000;
        x_t[34] = 11'b11111110000;
        x_t[35] = 11'b11111101110;
        x_t[36] = 11'b11111101111;
        x_t[37] = 11'b11111010011;
        x_t[38] = 11'b11111111111;
        x_t[39] = 11'b11111101000;
        x_t[40] = 11'b00000000110;
        x_t[41] = 11'b11111111100;
        x_t[42] = 11'b00000001010;
        x_t[43] = 11'b11111110110;
        x_t[44] = 11'b11111110010;
        x_t[45] = 11'b11111111101;
        x_t[46] = 11'b00000011000;
        x_t[47] = 11'b00000011101;
        x_t[48] = 11'b00000011100;
        x_t[49] = 11'b00000101001;
        x_t[50] = 11'b00000011111;
        x_t[51] = 11'b00000011011;
        x_t[52] = 11'b00000010111;
        x_t[53] = 11'b00000001110;
        x_t[54] = 11'b00000010011;
        x_t[55] = 11'b00000100100;
        x_t[56] = 11'b00000101100;
        x_t[57] = 11'b00000101111;
        x_t[58] = 11'b00000100010;
        x_t[59] = 11'b00000100011;
        x_t[60] = 11'b00000100011;
        x_t[61] = 11'b00000100001;
        x_t[62] = 11'b00000100001;
        x_t[63] = 11'b00000011110;
        
        h_t_prev[0] = 11'b11111101101;
        h_t_prev[1] = 11'b11111110101;
        h_t_prev[2] = 11'b11111110011;
        h_t_prev[3] = 11'b11111110100;
        h_t_prev[4] = 11'b11111110011;
        h_t_prev[5] = 11'b11111101100;
        h_t_prev[6] = 11'b11111100111;
        h_t_prev[7] = 11'b00000000101;
        h_t_prev[8] = 11'b11111111110;
        h_t_prev[9] = 11'b11111111110;
        h_t_prev[10] = 11'b00000000100;
        h_t_prev[11] = 11'b00000000110;
        h_t_prev[12] = 11'b11111111111;
        h_t_prev[13] = 11'b11111110011;
        h_t_prev[14] = 11'b00000001000;
        h_t_prev[15] = 11'b00000001000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 36 timeout!");
                $fdisplay(fd_cycles, "Test Vector  36: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  36: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 36");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 37
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111111100;
        x_t[1] = 11'b00000000110;
        x_t[2] = 11'b11111111111;
        x_t[3] = 11'b11111111100;
        x_t[4] = 11'b11111111000;
        x_t[5] = 11'b11111110001;
        x_t[6] = 11'b11111101111;
        x_t[7] = 11'b00000011000;
        x_t[8] = 11'b00000001011;
        x_t[9] = 11'b00000001000;
        x_t[10] = 11'b00000001010;
        x_t[11] = 11'b00000000010;
        x_t[12] = 11'b11111111101;
        x_t[13] = 11'b11111100111;
        x_t[14] = 11'b00000010111;
        x_t[15] = 11'b00000010011;
        x_t[16] = 11'b00000010000;
        x_t[17] = 11'b00000001011;
        x_t[18] = 11'b00000001101;
        x_t[19] = 11'b00000001010;
        x_t[20] = 11'b00000000001;
        x_t[21] = 11'b11111110011;
        x_t[22] = 11'b11111101011;
        x_t[23] = 11'b11111101110;
        x_t[24] = 11'b11111110100;
        x_t[25] = 11'b11111110110;
        x_t[26] = 11'b11111101101;
        x_t[27] = 11'b11111110000;
        x_t[28] = 11'b11111101010;
        x_t[29] = 11'b11111111111;
        x_t[30] = 11'b11111100001;
        x_t[31] = 11'b00000000100;
        x_t[32] = 11'b11111111110;
        x_t[33] = 11'b11111110100;
        x_t[34] = 11'b11111101101;
        x_t[35] = 11'b11111101011;
        x_t[36] = 11'b11111110000;
        x_t[37] = 11'b11111010100;
        x_t[38] = 11'b00000000100;
        x_t[39] = 11'b11111100011;
        x_t[40] = 11'b00000001110;
        x_t[41] = 11'b11111101010;
        x_t[42] = 11'b00000000111;
        x_t[43] = 11'b11111100011;
        x_t[44] = 11'b11111110111;
        x_t[45] = 11'b11111110101;
        x_t[46] = 11'b00000011111;
        x_t[47] = 11'b00000100010;
        x_t[48] = 11'b00000100010;
        x_t[49] = 11'b00000101010;
        x_t[50] = 11'b00000100000;
        x_t[51] = 11'b00000011010;
        x_t[52] = 11'b00000010100;
        x_t[53] = 11'b00000000111;
        x_t[54] = 11'b00000000100;
        x_t[55] = 11'b00000101100;
        x_t[56] = 11'b00000110010;
        x_t[57] = 11'b00000110110;
        x_t[58] = 11'b00000100000;
        x_t[59] = 11'b00000011011;
        x_t[60] = 11'b00000110111;
        x_t[61] = 11'b00000110001;
        x_t[62] = 11'b00000100111;
        x_t[63] = 11'b00000101100;
        
        h_t_prev[0] = 11'b11111111100;
        h_t_prev[1] = 11'b00000000110;
        h_t_prev[2] = 11'b11111111111;
        h_t_prev[3] = 11'b11111111100;
        h_t_prev[4] = 11'b11111111000;
        h_t_prev[5] = 11'b11111110001;
        h_t_prev[6] = 11'b11111101111;
        h_t_prev[7] = 11'b00000011000;
        h_t_prev[8] = 11'b00000001011;
        h_t_prev[9] = 11'b00000001000;
        h_t_prev[10] = 11'b00000001010;
        h_t_prev[11] = 11'b00000000010;
        h_t_prev[12] = 11'b11111111101;
        h_t_prev[13] = 11'b11111100111;
        h_t_prev[14] = 11'b00000010111;
        h_t_prev[15] = 11'b00000010011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 37 timeout!");
                $fdisplay(fd_cycles, "Test Vector  37: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  37: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 37");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 38
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000000010;
        x_t[1] = 11'b00000000010;
        x_t[2] = 11'b11111111001;
        x_t[3] = 11'b11111110010;
        x_t[4] = 11'b11111101110;
        x_t[5] = 11'b11111101000;
        x_t[6] = 11'b11111101001;
        x_t[7] = 11'b00000011001;
        x_t[8] = 11'b00000001010;
        x_t[9] = 11'b00000000011;
        x_t[10] = 11'b11111111111;
        x_t[11] = 11'b11111110011;
        x_t[12] = 11'b11111110011;
        x_t[13] = 11'b11111100011;
        x_t[14] = 11'b00000011100;
        x_t[15] = 11'b00000010101;
        x_t[16] = 11'b00000001110;
        x_t[17] = 11'b00000001000;
        x_t[18] = 11'b00000001000;
        x_t[19] = 11'b00000000100;
        x_t[20] = 11'b11111111111;
        x_t[21] = 11'b11111110101;
        x_t[22] = 11'b11111101101;
        x_t[23] = 11'b11111110001;
        x_t[24] = 11'b11111111000;
        x_t[25] = 11'b11111111010;
        x_t[26] = 11'b11111101101;
        x_t[27] = 11'b11111110010;
        x_t[28] = 11'b11111101110;
        x_t[29] = 11'b00000000111;
        x_t[30] = 11'b11111101101;
        x_t[31] = 11'b00000000100;
        x_t[32] = 11'b00000000000;
        x_t[33] = 11'b11111110111;
        x_t[34] = 11'b11111101111;
        x_t[35] = 11'b11111101110;
        x_t[36] = 11'b11111110001;
        x_t[37] = 11'b11111010110;
        x_t[38] = 11'b00000011000;
        x_t[39] = 11'b11111101100;
        x_t[40] = 11'b00000011101;
        x_t[41] = 11'b00000000110;
        x_t[42] = 11'b00000011000;
        x_t[43] = 11'b11111010100;
        x_t[44] = 11'b00000000001;
        x_t[45] = 11'b11111110100;
        x_t[46] = 11'b00000101110;
        x_t[47] = 11'b00000101110;
        x_t[48] = 11'b00000101100;
        x_t[49] = 11'b00000110011;
        x_t[50] = 11'b00000100101;
        x_t[51] = 11'b00000011110;
        x_t[52] = 11'b00000011001;
        x_t[53] = 11'b00000001011;
        x_t[54] = 11'b00000000100;
        x_t[55] = 11'b00000111001;
        x_t[56] = 11'b00000111100;
        x_t[57] = 11'b00000111110;
        x_t[58] = 11'b00000100011;
        x_t[59] = 11'b00000011110;
        x_t[60] = 11'b00001000011;
        x_t[61] = 11'b00000111001;
        x_t[62] = 11'b00000100110;
        x_t[63] = 11'b00000101110;
        
        h_t_prev[0] = 11'b00000000010;
        h_t_prev[1] = 11'b00000000010;
        h_t_prev[2] = 11'b11111111001;
        h_t_prev[3] = 11'b11111110010;
        h_t_prev[4] = 11'b11111101110;
        h_t_prev[5] = 11'b11111101000;
        h_t_prev[6] = 11'b11111101001;
        h_t_prev[7] = 11'b00000011001;
        h_t_prev[8] = 11'b00000001010;
        h_t_prev[9] = 11'b00000000011;
        h_t_prev[10] = 11'b11111111111;
        h_t_prev[11] = 11'b11111110011;
        h_t_prev[12] = 11'b11111110011;
        h_t_prev[13] = 11'b11111100011;
        h_t_prev[14] = 11'b00000011100;
        h_t_prev[15] = 11'b00000010101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 38 timeout!");
                $fdisplay(fd_cycles, "Test Vector  38: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  38: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 38");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 39
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000010011;
        x_t[1] = 11'b00000010010;
        x_t[2] = 11'b00000000110;
        x_t[3] = 11'b11111111101;
        x_t[4] = 11'b11111111000;
        x_t[5] = 11'b11111101111;
        x_t[6] = 11'b11111101110;
        x_t[7] = 11'b00000101101;
        x_t[8] = 11'b00000011101;
        x_t[9] = 11'b00000010011;
        x_t[10] = 11'b00000001011;
        x_t[11] = 11'b11111111101;
        x_t[12] = 11'b11111111011;
        x_t[13] = 11'b11111101110;
        x_t[14] = 11'b00000110000;
        x_t[15] = 11'b00000101000;
        x_t[16] = 11'b00000011101;
        x_t[17] = 11'b00000010100;
        x_t[18] = 11'b00000010010;
        x_t[19] = 11'b00000001110;
        x_t[20] = 11'b00000001001;
        x_t[21] = 11'b11111111100;
        x_t[22] = 11'b11111110001;
        x_t[23] = 11'b11111110100;
        x_t[24] = 11'b11111111110;
        x_t[25] = 11'b11111111111;
        x_t[26] = 11'b11111110011;
        x_t[27] = 11'b11111110101;
        x_t[28] = 11'b11111101101;
        x_t[29] = 11'b00000001101;
        x_t[30] = 11'b11111111001;
        x_t[31] = 11'b00000001001;
        x_t[32] = 11'b00000001000;
        x_t[33] = 11'b11111111110;
        x_t[34] = 11'b11111110110;
        x_t[35] = 11'b11111110011;
        x_t[36] = 11'b11111101101;
        x_t[37] = 11'b11111010001;
        x_t[38] = 11'b00000011100;
        x_t[39] = 11'b11111100101;
        x_t[40] = 11'b00000011100;
        x_t[41] = 11'b11111110011;
        x_t[42] = 11'b00000001110;
        x_t[43] = 11'b11111011011;
        x_t[44] = 11'b00000001111;
        x_t[45] = 11'b11111111000;
        x_t[46] = 11'b00000110110;
        x_t[47] = 11'b00000110111;
        x_t[48] = 11'b00000110101;
        x_t[49] = 11'b00000111100;
        x_t[50] = 11'b00000101101;
        x_t[51] = 11'b00000100101;
        x_t[52] = 11'b00000100000;
        x_t[53] = 11'b00000010011;
        x_t[54] = 11'b00000001101;
        x_t[55] = 11'b00000111101;
        x_t[56] = 11'b00001000000;
        x_t[57] = 11'b00001000001;
        x_t[58] = 11'b00000101000;
        x_t[59] = 11'b00000100101;
        x_t[60] = 11'b00001001000;
        x_t[61] = 11'b00000111110;
        x_t[62] = 11'b00000101001;
        x_t[63] = 11'b00000110011;
        
        h_t_prev[0] = 11'b00000010011;
        h_t_prev[1] = 11'b00000010010;
        h_t_prev[2] = 11'b00000000110;
        h_t_prev[3] = 11'b11111111101;
        h_t_prev[4] = 11'b11111111000;
        h_t_prev[5] = 11'b11111101111;
        h_t_prev[6] = 11'b11111101110;
        h_t_prev[7] = 11'b00000101101;
        h_t_prev[8] = 11'b00000011101;
        h_t_prev[9] = 11'b00000010011;
        h_t_prev[10] = 11'b00000001011;
        h_t_prev[11] = 11'b11111111101;
        h_t_prev[12] = 11'b11111111011;
        h_t_prev[13] = 11'b11111101110;
        h_t_prev[14] = 11'b00000110000;
        h_t_prev[15] = 11'b00000101000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 39 timeout!");
                $fdisplay(fd_cycles, "Test Vector  39: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  39: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 39");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 40
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000001111;
        x_t[1] = 11'b00000010011;
        x_t[2] = 11'b00000000110;
        x_t[3] = 11'b00000000001;
        x_t[4] = 11'b11111111011;
        x_t[5] = 11'b11111110000;
        x_t[6] = 11'b11111110000;
        x_t[7] = 11'b00000101001;
        x_t[8] = 11'b00000100000;
        x_t[9] = 11'b00000010110;
        x_t[10] = 11'b00000010100;
        x_t[11] = 11'b00000000110;
        x_t[12] = 11'b00000000011;
        x_t[13] = 11'b11111110011;
        x_t[14] = 11'b00000101011;
        x_t[15] = 11'b00000101010;
        x_t[16] = 11'b00000100011;
        x_t[17] = 11'b00000011001;
        x_t[18] = 11'b00000010111;
        x_t[19] = 11'b00000010010;
        x_t[20] = 11'b00000001100;
        x_t[21] = 11'b11111110111;
        x_t[22] = 11'b11111101011;
        x_t[23] = 11'b11111101110;
        x_t[24] = 11'b11111110111;
        x_t[25] = 11'b11111111001;
        x_t[26] = 11'b11111101010;
        x_t[27] = 11'b11111101101;
        x_t[28] = 11'b11111100110;
        x_t[29] = 11'b00000000011;
        x_t[30] = 11'b11111110011;
        x_t[31] = 11'b00000000010;
        x_t[32] = 11'b11111111101;
        x_t[33] = 11'b11111110011;
        x_t[34] = 11'b11111101101;
        x_t[35] = 11'b11111100111;
        x_t[36] = 11'b11111100110;
        x_t[37] = 11'b11111001110;
        x_t[38] = 11'b00000001111;
        x_t[39] = 11'b11111100000;
        x_t[40] = 11'b00000001100;
        x_t[41] = 11'b11111110101;
        x_t[42] = 11'b00000010100;
        x_t[43] = 11'b11111000110;
        x_t[44] = 11'b00000001110;
        x_t[45] = 11'b11111110001;
        x_t[46] = 11'b00000101000;
        x_t[47] = 11'b00000101110;
        x_t[48] = 11'b00000101111;
        x_t[49] = 11'b00000111000;
        x_t[50] = 11'b00000101001;
        x_t[51] = 11'b00000011111;
        x_t[52] = 11'b00000011010;
        x_t[53] = 11'b00000001100;
        x_t[54] = 11'b00000001100;
        x_t[55] = 11'b00000110111;
        x_t[56] = 11'b00000111011;
        x_t[57] = 11'b00000111011;
        x_t[58] = 11'b00000100010;
        x_t[59] = 11'b00000011111;
        x_t[60] = 11'b00001001000;
        x_t[61] = 11'b00000111111;
        x_t[62] = 11'b00000101111;
        x_t[63] = 11'b00000111010;
        
        h_t_prev[0] = 11'b00000001111;
        h_t_prev[1] = 11'b00000010011;
        h_t_prev[2] = 11'b00000000110;
        h_t_prev[3] = 11'b00000000001;
        h_t_prev[4] = 11'b11111111011;
        h_t_prev[5] = 11'b11111110000;
        h_t_prev[6] = 11'b11111110000;
        h_t_prev[7] = 11'b00000101001;
        h_t_prev[8] = 11'b00000100000;
        h_t_prev[9] = 11'b00000010110;
        h_t_prev[10] = 11'b00000010100;
        h_t_prev[11] = 11'b00000000110;
        h_t_prev[12] = 11'b00000000011;
        h_t_prev[13] = 11'b11111110011;
        h_t_prev[14] = 11'b00000101011;
        h_t_prev[15] = 11'b00000101010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 40 timeout!");
                $fdisplay(fd_cycles, "Test Vector  40: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  40: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 40");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 41
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000000011;
        x_t[1] = 11'b00000001001;
        x_t[2] = 11'b00000000010;
        x_t[3] = 11'b11111111101;
        x_t[4] = 11'b11111111001;
        x_t[5] = 11'b11111101101;
        x_t[6] = 11'b11111101011;
        x_t[7] = 11'b00000011011;
        x_t[8] = 11'b00000011001;
        x_t[9] = 11'b00000010100;
        x_t[10] = 11'b00000010101;
        x_t[11] = 11'b00000001001;
        x_t[12] = 11'b11111111110;
        x_t[13] = 11'b11111100100;
        x_t[14] = 11'b00000100101;
        x_t[15] = 11'b00000100110;
        x_t[16] = 11'b00000100000;
        x_t[17] = 11'b00000010101;
        x_t[18] = 11'b00000010011;
        x_t[19] = 11'b00000001010;
        x_t[20] = 11'b11111111100;
        x_t[21] = 11'b11111111000;
        x_t[22] = 11'b11111101101;
        x_t[23] = 11'b11111101111;
        x_t[24] = 11'b11111111001;
        x_t[25] = 11'b11111111011;
        x_t[26] = 11'b11111101101;
        x_t[27] = 11'b11111110000;
        x_t[28] = 11'b11111101011;
        x_t[29] = 11'b00000000110;
        x_t[30] = 11'b11111110111;
        x_t[31] = 11'b00000000111;
        x_t[32] = 11'b00000000101;
        x_t[33] = 11'b11111111100;
        x_t[34] = 11'b11111110100;
        x_t[35] = 11'b11111110001;
        x_t[36] = 11'b11111101101;
        x_t[37] = 11'b11111011011;
        x_t[38] = 11'b00000010000;
        x_t[39] = 11'b11111100111;
        x_t[40] = 11'b00000010100;
        x_t[41] = 11'b11111101001;
        x_t[42] = 11'b00000011011;
        x_t[43] = 11'b11111101000;
        x_t[44] = 11'b00000001101;
        x_t[45] = 11'b11111101110;
        x_t[46] = 11'b00000100110;
        x_t[47] = 11'b00000101101;
        x_t[48] = 11'b00000101110;
        x_t[49] = 11'b00000110100;
        x_t[50] = 11'b00000101000;
        x_t[51] = 11'b00000011010;
        x_t[52] = 11'b00000010011;
        x_t[53] = 11'b00000000011;
        x_t[54] = 11'b00000000100;
        x_t[55] = 11'b00000111001;
        x_t[56] = 11'b00000111100;
        x_t[57] = 11'b00000111000;
        x_t[58] = 11'b00000011011;
        x_t[59] = 11'b00000011001;
        x_t[60] = 11'b00001000011;
        x_t[61] = 11'b00000111001;
        x_t[62] = 11'b00000101110;
        x_t[63] = 11'b00000110011;
        
        h_t_prev[0] = 11'b00000000011;
        h_t_prev[1] = 11'b00000001001;
        h_t_prev[2] = 11'b00000000010;
        h_t_prev[3] = 11'b11111111101;
        h_t_prev[4] = 11'b11111111001;
        h_t_prev[5] = 11'b11111101101;
        h_t_prev[6] = 11'b11111101011;
        h_t_prev[7] = 11'b00000011011;
        h_t_prev[8] = 11'b00000011001;
        h_t_prev[9] = 11'b00000010100;
        h_t_prev[10] = 11'b00000010101;
        h_t_prev[11] = 11'b00000001001;
        h_t_prev[12] = 11'b11111111110;
        h_t_prev[13] = 11'b11111100100;
        h_t_prev[14] = 11'b00000100101;
        h_t_prev[15] = 11'b00000100110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 41 timeout!");
                $fdisplay(fd_cycles, "Test Vector  41: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  41: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 41");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 42
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000010001;
        x_t[1] = 11'b00000011101;
        x_t[2] = 11'b00000010111;
        x_t[3] = 11'b00000010011;
        x_t[4] = 11'b00000001011;
        x_t[5] = 11'b11111111011;
        x_t[6] = 11'b11111101111;
        x_t[7] = 11'b00000110010;
        x_t[8] = 11'b00000101100;
        x_t[9] = 11'b00000100111;
        x_t[10] = 11'b00000100010;
        x_t[11] = 11'b00000010111;
        x_t[12] = 11'b00000000110;
        x_t[13] = 11'b11111100011;
        x_t[14] = 11'b00000111100;
        x_t[15] = 11'b00000110100;
        x_t[16] = 11'b00000101101;
        x_t[17] = 11'b00000100001;
        x_t[18] = 11'b00000011101;
        x_t[19] = 11'b00000010010;
        x_t[20] = 11'b00000000001;
        x_t[21] = 11'b11111111001;
        x_t[22] = 11'b11111110000;
        x_t[23] = 11'b11111110100;
        x_t[24] = 11'b11111111110;
        x_t[25] = 11'b00000000000;
        x_t[26] = 11'b11111111010;
        x_t[27] = 11'b11111111010;
        x_t[28] = 11'b11111110010;
        x_t[29] = 11'b00000001110;
        x_t[30] = 11'b00000000000;
        x_t[31] = 11'b00000010110;
        x_t[32] = 11'b00000010011;
        x_t[33] = 11'b00000001011;
        x_t[34] = 11'b00000000011;
        x_t[35] = 11'b11111111101;
        x_t[36] = 11'b11111110110;
        x_t[37] = 11'b11111100000;
        x_t[38] = 11'b00000010101;
        x_t[39] = 11'b11111101011;
        x_t[40] = 11'b00000010011;
        x_t[41] = 11'b11111100111;
        x_t[42] = 11'b00000011111;
        x_t[43] = 11'b11111110010;
        x_t[44] = 11'b00000011100;
        x_t[45] = 11'b00000000001;
        x_t[46] = 11'b00000110111;
        x_t[47] = 11'b00000111100;
        x_t[48] = 11'b00000110111;
        x_t[49] = 11'b00001000000;
        x_t[50] = 11'b00000110011;
        x_t[51] = 11'b00000100111;
        x_t[52] = 11'b00000100010;
        x_t[53] = 11'b00000010001;
        x_t[54] = 11'b00000010001;
        x_t[55] = 11'b00001000011;
        x_t[56] = 11'b00001000110;
        x_t[57] = 11'b00001000001;
        x_t[58] = 11'b00000100011;
        x_t[59] = 11'b00000100000;
        x_t[60] = 11'b00001000011;
        x_t[61] = 11'b00000111000;
        x_t[62] = 11'b00000110000;
        x_t[63] = 11'b00000110100;
        
        h_t_prev[0] = 11'b00000010001;
        h_t_prev[1] = 11'b00000011101;
        h_t_prev[2] = 11'b00000010111;
        h_t_prev[3] = 11'b00000010011;
        h_t_prev[4] = 11'b00000001011;
        h_t_prev[5] = 11'b11111111011;
        h_t_prev[6] = 11'b11111101111;
        h_t_prev[7] = 11'b00000110010;
        h_t_prev[8] = 11'b00000101100;
        h_t_prev[9] = 11'b00000100111;
        h_t_prev[10] = 11'b00000100010;
        h_t_prev[11] = 11'b00000010111;
        h_t_prev[12] = 11'b00000000110;
        h_t_prev[13] = 11'b11111100011;
        h_t_prev[14] = 11'b00000111100;
        h_t_prev[15] = 11'b00000110100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 42 timeout!");
                $fdisplay(fd_cycles, "Test Vector  42: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  42: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 42");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 43
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000010110;
        x_t[1] = 11'b00000011011;
        x_t[2] = 11'b00000010101;
        x_t[3] = 11'b00000010101;
        x_t[4] = 11'b00000001110;
        x_t[5] = 11'b00000000001;
        x_t[6] = 11'b11111111100;
        x_t[7] = 11'b00000100111;
        x_t[8] = 11'b00000100011;
        x_t[9] = 11'b00000100000;
        x_t[10] = 11'b00000011111;
        x_t[11] = 11'b00000011001;
        x_t[12] = 11'b00000001101;
        x_t[13] = 11'b11111111000;
        x_t[14] = 11'b00000101100;
        x_t[15] = 11'b00000101001;
        x_t[16] = 11'b00000100111;
        x_t[17] = 11'b00000011101;
        x_t[18] = 11'b00000100001;
        x_t[19] = 11'b00000011100;
        x_t[20] = 11'b00000010010;
        x_t[21] = 11'b11111110110;
        x_t[22] = 11'b11111101100;
        x_t[23] = 11'b11111110010;
        x_t[24] = 11'b11111111001;
        x_t[25] = 11'b11111111011;
        x_t[26] = 11'b11111110011;
        x_t[27] = 11'b11111110111;
        x_t[28] = 11'b11111110001;
        x_t[29] = 11'b00000001110;
        x_t[30] = 11'b11111111101;
        x_t[31] = 11'b00000001111;
        x_t[32] = 11'b00000000111;
        x_t[33] = 11'b00000000010;
        x_t[34] = 11'b11111111100;
        x_t[35] = 11'b11111110110;
        x_t[36] = 11'b11111110011;
        x_t[37] = 11'b11111100001;
        x_t[38] = 11'b00000011100;
        x_t[39] = 11'b11111111000;
        x_t[40] = 11'b00000101001;
        x_t[41] = 11'b00000011011;
        x_t[42] = 11'b00000101101;
        x_t[43] = 11'b11111110101;
        x_t[44] = 11'b00000011110;
        x_t[45] = 11'b00000001101;
        x_t[46] = 11'b00000101100;
        x_t[47] = 11'b00000101101;
        x_t[48] = 11'b00000100110;
        x_t[49] = 11'b00000110101;
        x_t[50] = 11'b00000101000;
        x_t[51] = 11'b00000100010;
        x_t[52] = 11'b00000100001;
        x_t[53] = 11'b00000010101;
        x_t[54] = 11'b00000010110;
        x_t[55] = 11'b00000110100;
        x_t[56] = 11'b00000111001;
        x_t[57] = 11'b00000110111;
        x_t[58] = 11'b00000100001;
        x_t[59] = 11'b00000100000;
        x_t[60] = 11'b00001000010;
        x_t[61] = 11'b00000111001;
        x_t[62] = 11'b00000110001;
        x_t[63] = 11'b00000110101;
        
        h_t_prev[0] = 11'b00000010110;
        h_t_prev[1] = 11'b00000011011;
        h_t_prev[2] = 11'b00000010101;
        h_t_prev[3] = 11'b00000010101;
        h_t_prev[4] = 11'b00000001110;
        h_t_prev[5] = 11'b00000000001;
        h_t_prev[6] = 11'b11111111100;
        h_t_prev[7] = 11'b00000100111;
        h_t_prev[8] = 11'b00000100011;
        h_t_prev[9] = 11'b00000100000;
        h_t_prev[10] = 11'b00000011111;
        h_t_prev[11] = 11'b00000011001;
        h_t_prev[12] = 11'b00000001101;
        h_t_prev[13] = 11'b11111111000;
        h_t_prev[14] = 11'b00000101100;
        h_t_prev[15] = 11'b00000101001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 43 timeout!");
                $fdisplay(fd_cycles, "Test Vector  43: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  43: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 43");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 44
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000010100;
        x_t[1] = 11'b00000010101;
        x_t[2] = 11'b00000001110;
        x_t[3] = 11'b00000001111;
        x_t[4] = 11'b00000001001;
        x_t[5] = 11'b00000000000;
        x_t[6] = 11'b00000001000;
        x_t[7] = 11'b00000011110;
        x_t[8] = 11'b00000011010;
        x_t[9] = 11'b00000010111;
        x_t[10] = 11'b00000011001;
        x_t[11] = 11'b00000011010;
        x_t[12] = 11'b00000010010;
        x_t[13] = 11'b00000001101;
        x_t[14] = 11'b00000011111;
        x_t[15] = 11'b00000011111;
        x_t[16] = 11'b00000011110;
        x_t[17] = 11'b00000011001;
        x_t[18] = 11'b00000100001;
        x_t[19] = 11'b00000100000;
        x_t[20] = 11'b00000100010;
        x_t[21] = 11'b11111111010;
        x_t[22] = 11'b11111110000;
        x_t[23] = 11'b11111110100;
        x_t[24] = 11'b11111111111;
        x_t[25] = 11'b00000000000;
        x_t[26] = 11'b11111111001;
        x_t[27] = 11'b11111111010;
        x_t[28] = 11'b11111110010;
        x_t[29] = 11'b00000010100;
        x_t[30] = 11'b00000000011;
        x_t[31] = 11'b00000010100;
        x_t[32] = 11'b00000001111;
        x_t[33] = 11'b00000001001;
        x_t[34] = 11'b00000000011;
        x_t[35] = 11'b11111111111;
        x_t[36] = 11'b11111111100;
        x_t[37] = 11'b11111101001;
        x_t[38] = 11'b00000011110;
        x_t[39] = 11'b00000001010;
        x_t[40] = 11'b00000100100;
        x_t[41] = 11'b00000101011;
        x_t[42] = 11'b00000101101;
        x_t[43] = 11'b00000000110;
        x_t[44] = 11'b00000010010;
        x_t[45] = 11'b00000011011;
        x_t[46] = 11'b00000100111;
        x_t[47] = 11'b00000101010;
        x_t[48] = 11'b00000100101;
        x_t[49] = 11'b00000110011;
        x_t[50] = 11'b00000101001;
        x_t[51] = 11'b00000100110;
        x_t[52] = 11'b00000101001;
        x_t[53] = 11'b00000100001;
        x_t[54] = 11'b00000100011;
        x_t[55] = 11'b00000101111;
        x_t[56] = 11'b00000110011;
        x_t[57] = 11'b00000110100;
        x_t[58] = 11'b00000100101;
        x_t[59] = 11'b00000100110;
        x_t[60] = 11'b00000111011;
        x_t[61] = 11'b00000110101;
        x_t[62] = 11'b00000110011;
        x_t[63] = 11'b00000110000;
        
        h_t_prev[0] = 11'b00000010100;
        h_t_prev[1] = 11'b00000010101;
        h_t_prev[2] = 11'b00000001110;
        h_t_prev[3] = 11'b00000001111;
        h_t_prev[4] = 11'b00000001001;
        h_t_prev[5] = 11'b00000000000;
        h_t_prev[6] = 11'b00000001000;
        h_t_prev[7] = 11'b00000011110;
        h_t_prev[8] = 11'b00000011010;
        h_t_prev[9] = 11'b00000010111;
        h_t_prev[10] = 11'b00000011001;
        h_t_prev[11] = 11'b00000011010;
        h_t_prev[12] = 11'b00000010010;
        h_t_prev[13] = 11'b00000001101;
        h_t_prev[14] = 11'b00000011111;
        h_t_prev[15] = 11'b00000011111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 44 timeout!");
                $fdisplay(fd_cycles, "Test Vector  44: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  44: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 44");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 45
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000011100;
        x_t[1] = 11'b00000100000;
        x_t[2] = 11'b00000011100;
        x_t[3] = 11'b00000011010;
        x_t[4] = 11'b00000010011;
        x_t[5] = 11'b00000001100;
        x_t[6] = 11'b00000010010;
        x_t[7] = 11'b00000101001;
        x_t[8] = 11'b00000100110;
        x_t[9] = 11'b00000100001;
        x_t[10] = 11'b00000100001;
        x_t[11] = 11'b00000011111;
        x_t[12] = 11'b00000011100;
        x_t[13] = 11'b00000010000;
        x_t[14] = 11'b00000101000;
        x_t[15] = 11'b00000100100;
        x_t[16] = 11'b00000100001;
        x_t[17] = 11'b00000011101;
        x_t[18] = 11'b00000100010;
        x_t[19] = 11'b00000100010;
        x_t[20] = 11'b00000100100;
        x_t[21] = 11'b11111111011;
        x_t[22] = 11'b11111101111;
        x_t[23] = 11'b11111110001;
        x_t[24] = 11'b11111111110;
        x_t[25] = 11'b00000000001;
        x_t[26] = 11'b11111111100;
        x_t[27] = 11'b11111111101;
        x_t[28] = 11'b11111110001;
        x_t[29] = 11'b00000001111;
        x_t[30] = 11'b00000000110;
        x_t[31] = 11'b00000011011;
        x_t[32] = 11'b00000010010;
        x_t[33] = 11'b00000001011;
        x_t[34] = 11'b00000000110;
        x_t[35] = 11'b00000000010;
        x_t[36] = 11'b00000000010;
        x_t[37] = 11'b11111110011;
        x_t[38] = 11'b00000100010;
        x_t[39] = 11'b00000000111;
        x_t[40] = 11'b00000101010;
        x_t[41] = 11'b00000010101;
        x_t[42] = 11'b00000011100;
        x_t[43] = 11'b00000010110;
        x_t[44] = 11'b00000010001;
        x_t[45] = 11'b00000011100;
        x_t[46] = 11'b00000100011;
        x_t[47] = 11'b00000100011;
        x_t[48] = 11'b00000011110;
        x_t[49] = 11'b00000101001;
        x_t[50] = 11'b00000100000;
        x_t[51] = 11'b00000011100;
        x_t[52] = 11'b00000011110;
        x_t[53] = 11'b00000010111;
        x_t[54] = 11'b00000011001;
        x_t[55] = 11'b00000100001;
        x_t[56] = 11'b00000100101;
        x_t[57] = 11'b00000100011;
        x_t[58] = 11'b00000011000;
        x_t[59] = 11'b00000010101;
        x_t[60] = 11'b00000101010;
        x_t[61] = 11'b00000011111;
        x_t[62] = 11'b00000100100;
        x_t[63] = 11'b00000010111;
        
        h_t_prev[0] = 11'b00000011100;
        h_t_prev[1] = 11'b00000100000;
        h_t_prev[2] = 11'b00000011100;
        h_t_prev[3] = 11'b00000011010;
        h_t_prev[4] = 11'b00000010011;
        h_t_prev[5] = 11'b00000001100;
        h_t_prev[6] = 11'b00000010010;
        h_t_prev[7] = 11'b00000101001;
        h_t_prev[8] = 11'b00000100110;
        h_t_prev[9] = 11'b00000100001;
        h_t_prev[10] = 11'b00000100001;
        h_t_prev[11] = 11'b00000011111;
        h_t_prev[12] = 11'b00000011100;
        h_t_prev[13] = 11'b00000010000;
        h_t_prev[14] = 11'b00000101000;
        h_t_prev[15] = 11'b00000100100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 45 timeout!");
                $fdisplay(fd_cycles, "Test Vector  45: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  45: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 45");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 46
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000011010;
        x_t[1] = 11'b00000100001;
        x_t[2] = 11'b00000011010;
        x_t[3] = 11'b00000010111;
        x_t[4] = 11'b00000010000;
        x_t[5] = 11'b00000001010;
        x_t[6] = 11'b00000001110;
        x_t[7] = 11'b00000101101;
        x_t[8] = 11'b00000100111;
        x_t[9] = 11'b00000100011;
        x_t[10] = 11'b00000100011;
        x_t[11] = 11'b00000011011;
        x_t[12] = 11'b00000011010;
        x_t[13] = 11'b00000001100;
        x_t[14] = 11'b00000110000;
        x_t[15] = 11'b00000101000;
        x_t[16] = 11'b00000100011;
        x_t[17] = 11'b00000011110;
        x_t[18] = 11'b00000100010;
        x_t[19] = 11'b00000100001;
        x_t[20] = 11'b00000100001;
        x_t[21] = 11'b11111111011;
        x_t[22] = 11'b11111110001;
        x_t[23] = 11'b11111110000;
        x_t[24] = 11'b11111111110;
        x_t[25] = 11'b00000000001;
        x_t[26] = 11'b11111111101;
        x_t[27] = 11'b11111111111;
        x_t[28] = 11'b11111110011;
        x_t[29] = 11'b00000001110;
        x_t[30] = 11'b00000001011;
        x_t[31] = 11'b00000011011;
        x_t[32] = 11'b00000010110;
        x_t[33] = 11'b00000001101;
        x_t[34] = 11'b00000000110;
        x_t[35] = 11'b00000000011;
        x_t[36] = 11'b00000000000;
        x_t[37] = 11'b11111110101;
        x_t[38] = 11'b00000101001;
        x_t[39] = 11'b00000000101;
        x_t[40] = 11'b00000100101;
        x_t[41] = 11'b00000001100;
        x_t[42] = 11'b00000011111;
        x_t[43] = 11'b00000100011;
        x_t[44] = 11'b00000010110;
        x_t[45] = 11'b00000101011;
        x_t[46] = 11'b00000101010;
        x_t[47] = 11'b00000101010;
        x_t[48] = 11'b00000100100;
        x_t[49] = 11'b00000110000;
        x_t[50] = 11'b00000101001;
        x_t[51] = 11'b00000101000;
        x_t[52] = 11'b00000101001;
        x_t[53] = 11'b00000100011;
        x_t[54] = 11'b00000101000;
        x_t[55] = 11'b00000100011;
        x_t[56] = 11'b00000101000;
        x_t[57] = 11'b00000101010;
        x_t[58] = 11'b00000100011;
        x_t[59] = 11'b00000100000;
        x_t[60] = 11'b00000100000;
        x_t[61] = 11'b00000010011;
        x_t[62] = 11'b00000011100;
        x_t[63] = 11'b00000001101;
        
        h_t_prev[0] = 11'b00000011010;
        h_t_prev[1] = 11'b00000100001;
        h_t_prev[2] = 11'b00000011010;
        h_t_prev[3] = 11'b00000010111;
        h_t_prev[4] = 11'b00000010000;
        h_t_prev[5] = 11'b00000001010;
        h_t_prev[6] = 11'b00000001110;
        h_t_prev[7] = 11'b00000101101;
        h_t_prev[8] = 11'b00000100111;
        h_t_prev[9] = 11'b00000100011;
        h_t_prev[10] = 11'b00000100011;
        h_t_prev[11] = 11'b00000011011;
        h_t_prev[12] = 11'b00000011010;
        h_t_prev[13] = 11'b00000001100;
        h_t_prev[14] = 11'b00000110000;
        h_t_prev[15] = 11'b00000101000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 46 timeout!");
                $fdisplay(fd_cycles, "Test Vector  46: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  46: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 46");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 47
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000100110;
        x_t[1] = 11'b00000101100;
        x_t[2] = 11'b00000100011;
        x_t[3] = 11'b00000100100;
        x_t[4] = 11'b00000011010;
        x_t[5] = 11'b00000001110;
        x_t[6] = 11'b00000001101;
        x_t[7] = 11'b00000110100;
        x_t[8] = 11'b00000101101;
        x_t[9] = 11'b00000110001;
        x_t[10] = 11'b00000110000;
        x_t[11] = 11'b00000101011;
        x_t[12] = 11'b00000100010;
        x_t[13] = 11'b00000010001;
        x_t[14] = 11'b00000101011;
        x_t[15] = 11'b00000101101;
        x_t[16] = 11'b00000101101;
        x_t[17] = 11'b00000101010;
        x_t[18] = 11'b00000110000;
        x_t[19] = 11'b00000101101;
        x_t[20] = 11'b00000100111;
        x_t[21] = 11'b11111111011;
        x_t[22] = 11'b11111110011;
        x_t[23] = 11'b11111110011;
        x_t[24] = 11'b11111111110;
        x_t[25] = 11'b00000000001;
        x_t[26] = 11'b00000000010;
        x_t[27] = 11'b00000000000;
        x_t[28] = 11'b11111110101;
        x_t[29] = 11'b00000010111;
        x_t[30] = 11'b00000000011;
        x_t[31] = 11'b00000011010;
        x_t[32] = 11'b00000011000;
        x_t[33] = 11'b00000010000;
        x_t[34] = 11'b00000001000;
        x_t[35] = 11'b00000000010;
        x_t[36] = 11'b11111111101;
        x_t[37] = 11'b11111101110;
        x_t[38] = 11'b00000011011;
        x_t[39] = 11'b00000000011;
        x_t[40] = 11'b00000001001;
        x_t[41] = 11'b00000010100;
        x_t[42] = 11'b00000101110;
        x_t[43] = 11'b00000100000;
        x_t[44] = 11'b00000010010;
        x_t[45] = 11'b00000100110;
        x_t[46] = 11'b00000100001;
        x_t[47] = 11'b00000100010;
        x_t[48] = 11'b00000011111;
        x_t[49] = 11'b00000101001;
        x_t[50] = 11'b00000101000;
        x_t[51] = 11'b00000101001;
        x_t[52] = 11'b00000101001;
        x_t[53] = 11'b00000100001;
        x_t[54] = 11'b00000100010;
        x_t[55] = 11'b00000011011;
        x_t[56] = 11'b00000100100;
        x_t[57] = 11'b00000101000;
        x_t[58] = 11'b00000100101;
        x_t[59] = 11'b00000100001;
        x_t[60] = 11'b00000011100;
        x_t[61] = 11'b00000010011;
        x_t[62] = 11'b00000011110;
        x_t[63] = 11'b00000010011;
        
        h_t_prev[0] = 11'b00000100110;
        h_t_prev[1] = 11'b00000101100;
        h_t_prev[2] = 11'b00000100011;
        h_t_prev[3] = 11'b00000100100;
        h_t_prev[4] = 11'b00000011010;
        h_t_prev[5] = 11'b00000001110;
        h_t_prev[6] = 11'b00000001101;
        h_t_prev[7] = 11'b00000110100;
        h_t_prev[8] = 11'b00000101101;
        h_t_prev[9] = 11'b00000110001;
        h_t_prev[10] = 11'b00000110000;
        h_t_prev[11] = 11'b00000101011;
        h_t_prev[12] = 11'b00000100010;
        h_t_prev[13] = 11'b00000010001;
        h_t_prev[14] = 11'b00000101011;
        h_t_prev[15] = 11'b00000101101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 47 timeout!");
                $fdisplay(fd_cycles, "Test Vector  47: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  47: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 47");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 48
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000010101;
        x_t[1] = 11'b00000011100;
        x_t[2] = 11'b00000011001;
        x_t[3] = 11'b00000100000;
        x_t[4] = 11'b00000011001;
        x_t[5] = 11'b00000001100;
        x_t[6] = 11'b00000001111;
        x_t[7] = 11'b00000010111;
        x_t[8] = 11'b00000100000;
        x_t[9] = 11'b00000100100;
        x_t[10] = 11'b00000100110;
        x_t[11] = 11'b00000100010;
        x_t[12] = 11'b00000100001;
        x_t[13] = 11'b00000010000;
        x_t[14] = 11'b00000011101;
        x_t[15] = 11'b00000100010;
        x_t[16] = 11'b00000100100;
        x_t[17] = 11'b00000100001;
        x_t[18] = 11'b00000101011;
        x_t[19] = 11'b00000101000;
        x_t[20] = 11'b00000100011;
        x_t[21] = 11'b11111111010;
        x_t[22] = 11'b11111110010;
        x_t[23] = 11'b11111110011;
        x_t[24] = 11'b11111111100;
        x_t[25] = 11'b11111111110;
        x_t[26] = 11'b11111111111;
        x_t[27] = 11'b00000000000;
        x_t[28] = 11'b11111110100;
        x_t[29] = 11'b00000010011;
        x_t[30] = 11'b11111111111;
        x_t[31] = 11'b00000011001;
        x_t[32] = 11'b00000010000;
        x_t[33] = 11'b00000001011;
        x_t[34] = 11'b00000000110;
        x_t[35] = 11'b11111111111;
        x_t[36] = 11'b11111111111;
        x_t[37] = 11'b11111110100;
        x_t[38] = 11'b00000010111;
        x_t[39] = 11'b00000001000;
        x_t[40] = 11'b00000011100;
        x_t[41] = 11'b00000100000;
        x_t[42] = 11'b00000110001;
        x_t[43] = 11'b11111110101;
        x_t[44] = 11'b00000011010;
        x_t[45] = 11'b00000100111;
        x_t[46] = 11'b00000011011;
        x_t[47] = 11'b00000100010;
        x_t[48] = 11'b00000011111;
        x_t[49] = 11'b00000101010;
        x_t[50] = 11'b00000101001;
        x_t[51] = 11'b00000101111;
        x_t[52] = 11'b00000101101;
        x_t[53] = 11'b00000100111;
        x_t[54] = 11'b00000101000;
        x_t[55] = 11'b00000011101;
        x_t[56] = 11'b00000100111;
        x_t[57] = 11'b00000110000;
        x_t[58] = 11'b00000110000;
        x_t[59] = 11'b00000101101;
        x_t[60] = 11'b00000011110;
        x_t[61] = 11'b00000011101;
        x_t[62] = 11'b00000101011;
        x_t[63] = 11'b00000100011;
        
        h_t_prev[0] = 11'b00000010101;
        h_t_prev[1] = 11'b00000011100;
        h_t_prev[2] = 11'b00000011001;
        h_t_prev[3] = 11'b00000100000;
        h_t_prev[4] = 11'b00000011001;
        h_t_prev[5] = 11'b00000001100;
        h_t_prev[6] = 11'b00000001111;
        h_t_prev[7] = 11'b00000010111;
        h_t_prev[8] = 11'b00000100000;
        h_t_prev[9] = 11'b00000100100;
        h_t_prev[10] = 11'b00000100110;
        h_t_prev[11] = 11'b00000100010;
        h_t_prev[12] = 11'b00000100001;
        h_t_prev[13] = 11'b00000010000;
        h_t_prev[14] = 11'b00000011101;
        h_t_prev[15] = 11'b00000100010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 48 timeout!");
                $fdisplay(fd_cycles, "Test Vector  48: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  48: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 48");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 49
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111100111;
        x_t[1] = 11'b11111011000;
        x_t[2] = 11'b11111000111;
        x_t[3] = 11'b11110111000;
        x_t[4] = 11'b11110111100;
        x_t[5] = 11'b11110111000;
        x_t[6] = 11'b11111000110;
        x_t[7] = 11'b11111101111;
        x_t[8] = 11'b11111000110;
        x_t[9] = 11'b11111000010;
        x_t[10] = 11'b11110111101;
        x_t[11] = 11'b11110110101;
        x_t[12] = 11'b11111000000;
        x_t[13] = 11'b11110110111;
        x_t[14] = 11'b11111010010;
        x_t[15] = 11'b11111001100;
        x_t[16] = 11'b11111000100;
        x_t[17] = 11'b11111000000;
        x_t[18] = 11'b11111001011;
        x_t[19] = 11'b11111001111;
        x_t[20] = 11'b11111001011;
        x_t[21] = 11'b11111101011;
        x_t[22] = 11'b11111011010;
        x_t[23] = 11'b11111011001;
        x_t[24] = 11'b11111111001;
        x_t[25] = 11'b11111110111;
        x_t[26] = 11'b11111000010;
        x_t[27] = 11'b11110111111;
        x_t[28] = 11'b11111010100;
        x_t[29] = 11'b11111101110;
        x_t[30] = 11'b11111100101;
        x_t[31] = 11'b11110111101;
        x_t[32] = 11'b11111000001;
        x_t[33] = 11'b11110111001;
        x_t[34] = 11'b11110110110;
        x_t[35] = 11'b11111000000;
        x_t[36] = 11'b11110111010;
        x_t[37] = 11'b11111101000;
        x_t[38] = 11'b11111011110;
        x_t[39] = 11'b11110110101;
        x_t[40] = 11'b11111001101;
        x_t[41] = 11'b11110110110;
        x_t[42] = 11'b11111010110;
        x_t[43] = 11'b11111100011;
        x_t[44] = 11'b11111011010;
        x_t[45] = 11'b11111100001;
        x_t[46] = 11'b11111011001;
        x_t[47] = 11'b11111010101;
        x_t[48] = 11'b11111010010;
        x_t[49] = 11'b11111001111;
        x_t[50] = 11'b11111001001;
        x_t[51] = 11'b11111011010;
        x_t[52] = 11'b11111100000;
        x_t[53] = 11'b11111101010;
        x_t[54] = 11'b11111100000;
        x_t[55] = 11'b11111110100;
        x_t[56] = 11'b11111100010;
        x_t[57] = 11'b11111100101;
        x_t[58] = 11'b11111110010;
        x_t[59] = 11'b11111110100;
        x_t[60] = 11'b00000000111;
        x_t[61] = 11'b11111110110;
        x_t[62] = 11'b00000000100;
        x_t[63] = 11'b00000001001;
        
        h_t_prev[0] = 11'b11111100111;
        h_t_prev[1] = 11'b11111011000;
        h_t_prev[2] = 11'b11111000111;
        h_t_prev[3] = 11'b11110111000;
        h_t_prev[4] = 11'b11110111100;
        h_t_prev[5] = 11'b11110111000;
        h_t_prev[6] = 11'b11111000110;
        h_t_prev[7] = 11'b11111101111;
        h_t_prev[8] = 11'b11111000110;
        h_t_prev[9] = 11'b11111000010;
        h_t_prev[10] = 11'b11110111101;
        h_t_prev[11] = 11'b11110110101;
        h_t_prev[12] = 11'b11111000000;
        h_t_prev[13] = 11'b11110110111;
        h_t_prev[14] = 11'b11111010010;
        h_t_prev[15] = 11'b11111001100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 49 timeout!");
                $fdisplay(fd_cycles, "Test Vector  49: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  49: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 49");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 50
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111010111;
        x_t[1] = 11'b11111001010;
        x_t[2] = 11'b11110110101;
        x_t[3] = 11'b11110100100;
        x_t[4] = 11'b11110100100;
        x_t[5] = 11'b11110011100;
        x_t[6] = 11'b11110110011;
        x_t[7] = 11'b11111100000;
        x_t[8] = 11'b11110111001;
        x_t[9] = 11'b11110110100;
        x_t[10] = 11'b11110101110;
        x_t[11] = 11'b11110101001;
        x_t[12] = 11'b11110101001;
        x_t[13] = 11'b11110101011;
        x_t[14] = 11'b11111001001;
        x_t[15] = 11'b11111000001;
        x_t[16] = 11'b11110111010;
        x_t[17] = 11'b11110110110;
        x_t[18] = 11'b11110111110;
        x_t[19] = 11'b11110111111;
        x_t[20] = 11'b11110111110;
        x_t[21] = 11'b11111100110;
        x_t[22] = 11'b11111010111;
        x_t[23] = 11'b11111010111;
        x_t[24] = 11'b11111110111;
        x_t[25] = 11'b11111110110;
        x_t[26] = 11'b11110111001;
        x_t[27] = 11'b11110110111;
        x_t[28] = 11'b11111010010;
        x_t[29] = 11'b11111101110;
        x_t[30] = 11'b11111100100;
        x_t[31] = 11'b11110110011;
        x_t[32] = 11'b11110111000;
        x_t[33] = 11'b11110101110;
        x_t[34] = 11'b11110101011;
        x_t[35] = 11'b11110110101;
        x_t[36] = 11'b11110110000;
        x_t[37] = 11'b11111100101;
        x_t[38] = 11'b11111100000;
        x_t[39] = 11'b11110110001;
        x_t[40] = 11'b11111010001;
        x_t[41] = 11'b11110101000;
        x_t[42] = 11'b11111101110;
        x_t[43] = 11'b11111000011;
        x_t[44] = 11'b11111100100;
        x_t[45] = 11'b11111011101;
        x_t[46] = 11'b11111100010;
        x_t[47] = 11'b11111011001;
        x_t[48] = 11'b11111010101;
        x_t[49] = 11'b11111010101;
        x_t[50] = 11'b11111001111;
        x_t[51] = 11'b11111011111;
        x_t[52] = 11'b11111100010;
        x_t[53] = 11'b11111101010;
        x_t[54] = 11'b11111100011;
        x_t[55] = 11'b11111110111;
        x_t[56] = 11'b11111100110;
        x_t[57] = 11'b11111110000;
        x_t[58] = 11'b11111110011;
        x_t[59] = 11'b11111110010;
        x_t[60] = 11'b11111111100;
        x_t[61] = 11'b11111101111;
        x_t[62] = 11'b11111111001;
        x_t[63] = 11'b11111110011;
        
        h_t_prev[0] = 11'b11111010111;
        h_t_prev[1] = 11'b11111001010;
        h_t_prev[2] = 11'b11110110101;
        h_t_prev[3] = 11'b11110100100;
        h_t_prev[4] = 11'b11110100100;
        h_t_prev[5] = 11'b11110011100;
        h_t_prev[6] = 11'b11110110011;
        h_t_prev[7] = 11'b11111100000;
        h_t_prev[8] = 11'b11110111001;
        h_t_prev[9] = 11'b11110110100;
        h_t_prev[10] = 11'b11110101110;
        h_t_prev[11] = 11'b11110101001;
        h_t_prev[12] = 11'b11110101001;
        h_t_prev[13] = 11'b11110101011;
        h_t_prev[14] = 11'b11111001001;
        h_t_prev[15] = 11'b11111000001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 50 timeout!");
                $fdisplay(fd_cycles, "Test Vector  50: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  50: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 50");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 51
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111011001;
        x_t[1] = 11'b11111001001;
        x_t[2] = 11'b11110111001;
        x_t[3] = 11'b11110101010;
        x_t[4] = 11'b11110101001;
        x_t[5] = 11'b11110100110;
        x_t[6] = 11'b11110111010;
        x_t[7] = 11'b11111100101;
        x_t[8] = 11'b11111000100;
        x_t[9] = 11'b11110111111;
        x_t[10] = 11'b11110111100;
        x_t[11] = 11'b11110110111;
        x_t[12] = 11'b11110110000;
        x_t[13] = 11'b11110110010;
        x_t[14] = 11'b11111011000;
        x_t[15] = 11'b11111001111;
        x_t[16] = 11'b11111001010;
        x_t[17] = 11'b11111000110;
        x_t[18] = 11'b11111001100;
        x_t[19] = 11'b11111001011;
        x_t[20] = 11'b11111000101;
        x_t[21] = 11'b11111101010;
        x_t[22] = 11'b11111011011;
        x_t[23] = 11'b11111011011;
        x_t[24] = 11'b11111111100;
        x_t[25] = 11'b11111111011;
        x_t[26] = 11'b11111000010;
        x_t[27] = 11'b11110111111;
        x_t[28] = 11'b11111010101;
        x_t[29] = 11'b11111110110;
        x_t[30] = 11'b11111101101;
        x_t[31] = 11'b11111000001;
        x_t[32] = 11'b11111000100;
        x_t[33] = 11'b11110111001;
        x_t[34] = 11'b11110111000;
        x_t[35] = 11'b11111000011;
        x_t[36] = 11'b11110111101;
        x_t[37] = 11'b11111110011;
        x_t[38] = 11'b11111110011;
        x_t[39] = 11'b11111000111;
        x_t[40] = 11'b11111110111;
        x_t[41] = 11'b11111000001;
        x_t[42] = 11'b11111110101;
        x_t[43] = 11'b11111001101;
        x_t[44] = 11'b11111110111;
        x_t[45] = 11'b11111110100;
        x_t[46] = 11'b11111110010;
        x_t[47] = 11'b11111101010;
        x_t[48] = 11'b11111100111;
        x_t[49] = 11'b11111101010;
        x_t[50] = 11'b11111100111;
        x_t[51] = 11'b11111110010;
        x_t[52] = 11'b11111110010;
        x_t[53] = 11'b11111110111;
        x_t[54] = 11'b11111110010;
        x_t[55] = 11'b11111111010;
        x_t[56] = 11'b11111101110;
        x_t[57] = 11'b00000000000;
        x_t[58] = 11'b11111111101;
        x_t[59] = 11'b11111110101;
        x_t[60] = 11'b11111111000;
        x_t[61] = 11'b11111110001;
        x_t[62] = 11'b11111111001;
        x_t[63] = 11'b11111101111;
        
        h_t_prev[0] = 11'b11111011001;
        h_t_prev[1] = 11'b11111001001;
        h_t_prev[2] = 11'b11110111001;
        h_t_prev[3] = 11'b11110101010;
        h_t_prev[4] = 11'b11110101001;
        h_t_prev[5] = 11'b11110100110;
        h_t_prev[6] = 11'b11110111010;
        h_t_prev[7] = 11'b11111100101;
        h_t_prev[8] = 11'b11111000100;
        h_t_prev[9] = 11'b11110111111;
        h_t_prev[10] = 11'b11110111100;
        h_t_prev[11] = 11'b11110110111;
        h_t_prev[12] = 11'b11110110000;
        h_t_prev[13] = 11'b11110110010;
        h_t_prev[14] = 11'b11111011000;
        h_t_prev[15] = 11'b11111001111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 51 timeout!");
                $fdisplay(fd_cycles, "Test Vector  51: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  51: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 51");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 52
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111101101;
        x_t[1] = 11'b11111100001;
        x_t[2] = 11'b11111010000;
        x_t[3] = 11'b11111000000;
        x_t[4] = 11'b11111000000;
        x_t[5] = 11'b11110111110;
        x_t[6] = 11'b11111010110;
        x_t[7] = 11'b00000000110;
        x_t[8] = 11'b11111011111;
        x_t[9] = 11'b11111011110;
        x_t[10] = 11'b11111011010;
        x_t[11] = 11'b11111001100;
        x_t[12] = 11'b11111001011;
        x_t[13] = 11'b11111001001;
        x_t[14] = 11'b11111110110;
        x_t[15] = 11'b11111101011;
        x_t[16] = 11'b11111100101;
        x_t[17] = 11'b11111100011;
        x_t[18] = 11'b11111100101;
        x_t[19] = 11'b11111100010;
        x_t[20] = 11'b11111010111;
        x_t[21] = 11'b11111110000;
        x_t[22] = 11'b11111100010;
        x_t[23] = 11'b11111100001;
        x_t[24] = 11'b00000000011;
        x_t[25] = 11'b00000000010;
        x_t[26] = 11'b11111001010;
        x_t[27] = 11'b11111001000;
        x_t[28] = 11'b11111011011;
        x_t[29] = 11'b11111111111;
        x_t[30] = 11'b11111110101;
        x_t[31] = 11'b11111001011;
        x_t[32] = 11'b11111010011;
        x_t[33] = 11'b11111001000;
        x_t[34] = 11'b11111000101;
        x_t[35] = 11'b11111010001;
        x_t[36] = 11'b11111001110;
        x_t[37] = 11'b11111111110;
        x_t[38] = 11'b00000000010;
        x_t[39] = 11'b11111010110;
        x_t[40] = 11'b11111111000;
        x_t[41] = 11'b11111100000;
        x_t[42] = 11'b11111110111;
        x_t[43] = 11'b00000000000;
        x_t[44] = 11'b11111111110;
        x_t[45] = 11'b11111111000;
        x_t[46] = 11'b11111101101;
        x_t[47] = 11'b11111101110;
        x_t[48] = 11'b11111101101;
        x_t[49] = 11'b11111110000;
        x_t[50] = 11'b11111110011;
        x_t[51] = 11'b11111111000;
        x_t[52] = 11'b11111110111;
        x_t[53] = 11'b11111111000;
        x_t[54] = 11'b11111101111;
        x_t[55] = 11'b11111110100;
        x_t[56] = 11'b11111101011;
        x_t[57] = 11'b00000000001;
        x_t[58] = 11'b11111111001;
        x_t[59] = 11'b11111101010;
        x_t[60] = 11'b11111110101;
        x_t[61] = 11'b11111110001;
        x_t[62] = 11'b11111111011;
        x_t[63] = 11'b11111101110;
        
        h_t_prev[0] = 11'b11111101101;
        h_t_prev[1] = 11'b11111100001;
        h_t_prev[2] = 11'b11111010000;
        h_t_prev[3] = 11'b11111000000;
        h_t_prev[4] = 11'b11111000000;
        h_t_prev[5] = 11'b11110111110;
        h_t_prev[6] = 11'b11111010110;
        h_t_prev[7] = 11'b00000000110;
        h_t_prev[8] = 11'b11111011111;
        h_t_prev[9] = 11'b11111011110;
        h_t_prev[10] = 11'b11111011010;
        h_t_prev[11] = 11'b11111001100;
        h_t_prev[12] = 11'b11111001011;
        h_t_prev[13] = 11'b11111001001;
        h_t_prev[14] = 11'b11111110110;
        h_t_prev[15] = 11'b11111101011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 52 timeout!");
                $fdisplay(fd_cycles, "Test Vector  52: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  52: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 52");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 53
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111111101;
        x_t[1] = 11'b11111110000;
        x_t[2] = 11'b11111100001;
        x_t[3] = 11'b11111010110;
        x_t[4] = 11'b11111010110;
        x_t[5] = 11'b11111010010;
        x_t[6] = 11'b11111101001;
        x_t[7] = 11'b00000001101;
        x_t[8] = 11'b11111100110;
        x_t[9] = 11'b11111101100;
        x_t[10] = 11'b11111101100;
        x_t[11] = 11'b11111011011;
        x_t[12] = 11'b11111011101;
        x_t[13] = 11'b11111011001;
        x_t[14] = 11'b11111101110;
        x_t[15] = 11'b11111101101;
        x_t[16] = 11'b11111101101;
        x_t[17] = 11'b11111101100;
        x_t[18] = 11'b11111101101;
        x_t[19] = 11'b11111101001;
        x_t[20] = 11'b11111011111;
        x_t[21] = 11'b11111110100;
        x_t[22] = 11'b11111101000;
        x_t[23] = 11'b11111101001;
        x_t[24] = 11'b00000000110;
        x_t[25] = 11'b00000000101;
        x_t[26] = 11'b11111010100;
        x_t[27] = 11'b11111010011;
        x_t[28] = 11'b11111100101;
        x_t[29] = 11'b00000000010;
        x_t[30] = 11'b11111111110;
        x_t[31] = 11'b11111011001;
        x_t[32] = 11'b11111011100;
        x_t[33] = 11'b11111010100;
        x_t[34] = 11'b11111010001;
        x_t[35] = 11'b11111011100;
        x_t[36] = 11'b11111011100;
        x_t[37] = 11'b00000000111;
        x_t[38] = 11'b00000000001;
        x_t[39] = 11'b11111100001;
        x_t[40] = 11'b11111110011;
        x_t[41] = 11'b11111011101;
        x_t[42] = 11'b00000001111;
        x_t[43] = 11'b11111111011;
        x_t[44] = 11'b00000000101;
        x_t[45] = 11'b11111101111;
        x_t[46] = 11'b11111101101;
        x_t[47] = 11'b11111101010;
        x_t[48] = 11'b11111101001;
        x_t[49] = 11'b11111101110;
        x_t[50] = 11'b11111110011;
        x_t[51] = 11'b11111110110;
        x_t[52] = 11'b11111110011;
        x_t[53] = 11'b11111110011;
        x_t[54] = 11'b11111100000;
        x_t[55] = 11'b11111101100;
        x_t[56] = 11'b11111100011;
        x_t[57] = 11'b11111111010;
        x_t[58] = 11'b11111101101;
        x_t[59] = 11'b11111011110;
        x_t[60] = 11'b11111101101;
        x_t[61] = 11'b11111101001;
        x_t[62] = 11'b11111110001;
        x_t[63] = 11'b11111100111;
        
        h_t_prev[0] = 11'b11111111101;
        h_t_prev[1] = 11'b11111110000;
        h_t_prev[2] = 11'b11111100001;
        h_t_prev[3] = 11'b11111010110;
        h_t_prev[4] = 11'b11111010110;
        h_t_prev[5] = 11'b11111010010;
        h_t_prev[6] = 11'b11111101001;
        h_t_prev[7] = 11'b00000001101;
        h_t_prev[8] = 11'b11111100110;
        h_t_prev[9] = 11'b11111101100;
        h_t_prev[10] = 11'b11111101100;
        h_t_prev[11] = 11'b11111011011;
        h_t_prev[12] = 11'b11111011101;
        h_t_prev[13] = 11'b11111011001;
        h_t_prev[14] = 11'b11111101110;
        h_t_prev[15] = 11'b11111101101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 53 timeout!");
                $fdisplay(fd_cycles, "Test Vector  53: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  53: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 53");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 54
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111111011;
        x_t[1] = 11'b11111101111;
        x_t[2] = 11'b11111100010;
        x_t[3] = 11'b11111011010;
        x_t[4] = 11'b11111011001;
        x_t[5] = 11'b11111010100;
        x_t[6] = 11'b11111100110;
        x_t[7] = 11'b00000001000;
        x_t[8] = 11'b11111100100;
        x_t[9] = 11'b11111101000;
        x_t[10] = 11'b11111100110;
        x_t[11] = 11'b11111010110;
        x_t[12] = 11'b11111011011;
        x_t[13] = 11'b11111011100;
        x_t[14] = 11'b11111101101;
        x_t[15] = 11'b11111101001;
        x_t[16] = 11'b11111101001;
        x_t[17] = 11'b11111100101;
        x_t[18] = 11'b11111100101;
        x_t[19] = 11'b11111100001;
        x_t[20] = 11'b11111011000;
        x_t[21] = 11'b11111110101;
        x_t[22] = 11'b11111101001;
        x_t[23] = 11'b11111101100;
        x_t[24] = 11'b00000000110;
        x_t[25] = 11'b00000000101;
        x_t[26] = 11'b11111010100;
        x_t[27] = 11'b11111010111;
        x_t[28] = 11'b11111101000;
        x_t[29] = 11'b00000000011;
        x_t[30] = 11'b11111111111;
        x_t[31] = 11'b11111011010;
        x_t[32] = 11'b11111011011;
        x_t[33] = 11'b11111010010;
        x_t[34] = 11'b11111010001;
        x_t[35] = 11'b11111011101;
        x_t[36] = 11'b11111011100;
        x_t[37] = 11'b00000001101;
        x_t[38] = 11'b11111111111;
        x_t[39] = 11'b11111100010;
        x_t[40] = 11'b00000001011;
        x_t[41] = 11'b11111011000;
        x_t[42] = 11'b00000001001;
        x_t[43] = 11'b11111001011;
        x_t[44] = 11'b00000010100;
        x_t[45] = 11'b11111011001;
        x_t[46] = 11'b11111110001;
        x_t[47] = 11'b11111101011;
        x_t[48] = 11'b11111100111;
        x_t[49] = 11'b11111101000;
        x_t[50] = 11'b11111100111;
        x_t[51] = 11'b11111100101;
        x_t[52] = 11'b11111100001;
        x_t[53] = 11'b11111100000;
        x_t[54] = 11'b11111010001;
        x_t[55] = 11'b11111100110;
        x_t[56] = 11'b11111011101;
        x_t[57] = 11'b11111101110;
        x_t[58] = 11'b11111011000;
        x_t[59] = 11'b11111001111;
        x_t[60] = 11'b11111100010;
        x_t[61] = 11'b11111011010;
        x_t[62] = 11'b11111011011;
        x_t[63] = 11'b11111011110;
        
        h_t_prev[0] = 11'b11111111011;
        h_t_prev[1] = 11'b11111101111;
        h_t_prev[2] = 11'b11111100010;
        h_t_prev[3] = 11'b11111011010;
        h_t_prev[4] = 11'b11111011001;
        h_t_prev[5] = 11'b11111010100;
        h_t_prev[6] = 11'b11111100110;
        h_t_prev[7] = 11'b00000001000;
        h_t_prev[8] = 11'b11111100100;
        h_t_prev[9] = 11'b11111101000;
        h_t_prev[10] = 11'b11111100110;
        h_t_prev[11] = 11'b11111010110;
        h_t_prev[12] = 11'b11111011011;
        h_t_prev[13] = 11'b11111011100;
        h_t_prev[14] = 11'b11111101101;
        h_t_prev[15] = 11'b11111101001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 54 timeout!");
                $fdisplay(fd_cycles, "Test Vector  54: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  54: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 54");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 55
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111111010;
        x_t[1] = 11'b11111101100;
        x_t[2] = 11'b11111011100;
        x_t[3] = 11'b11111010001;
        x_t[4] = 11'b11111010001;
        x_t[5] = 11'b11111001101;
        x_t[6] = 11'b11111011101;
        x_t[7] = 11'b00000000111;
        x_t[8] = 11'b11111100110;
        x_t[9] = 11'b11111100010;
        x_t[10] = 11'b11111011100;
        x_t[11] = 11'b11111001010;
        x_t[12] = 11'b11111010100;
        x_t[13] = 11'b11111010000;
        x_t[14] = 11'b11111111000;
        x_t[15] = 11'b11111101000;
        x_t[16] = 11'b11111100010;
        x_t[17] = 11'b11111011010;
        x_t[18] = 11'b11111011011;
        x_t[19] = 11'b11111010111;
        x_t[20] = 11'b11111001111;
        x_t[21] = 11'b11111110100;
        x_t[22] = 11'b11111100111;
        x_t[23] = 11'b11111100111;
        x_t[24] = 11'b00000000110;
        x_t[25] = 11'b00000000101;
        x_t[26] = 11'b11111010000;
        x_t[27] = 11'b11111010001;
        x_t[28] = 11'b11111100011;
        x_t[29] = 11'b00000000100;
        x_t[30] = 11'b11111111010;
        x_t[31] = 11'b11111010010;
        x_t[32] = 11'b11111010111;
        x_t[33] = 11'b11111001100;
        x_t[34] = 11'b11111001010;
        x_t[35] = 11'b11111010111;
        x_t[36] = 11'b11111010001;
        x_t[37] = 11'b00000000001;
        x_t[38] = 11'b00000001001;
        x_t[39] = 11'b11111001110;
        x_t[40] = 11'b00000010110;
        x_t[41] = 11'b11110100110;
        x_t[42] = 11'b00000010001;
        x_t[43] = 11'b11111110111;
        x_t[44] = 11'b00000010011;
        x_t[45] = 11'b11111100100;
        x_t[46] = 11'b11111101111;
        x_t[47] = 11'b11111101001;
        x_t[48] = 11'b11111100011;
        x_t[49] = 11'b11111100000;
        x_t[50] = 11'b11111011101;
        x_t[51] = 11'b11111011000;
        x_t[52] = 11'b11111011000;
        x_t[53] = 11'b11111011100;
        x_t[54] = 11'b11111010111;
        x_t[55] = 11'b11111100010;
        x_t[56] = 11'b11111011010;
        x_t[57] = 11'b11111100011;
        x_t[58] = 11'b11111010000;
        x_t[59] = 11'b11111001111;
        x_t[60] = 11'b11111011001;
        x_t[61] = 11'b11111001111;
        x_t[62] = 11'b11111001001;
        x_t[63] = 11'b11111011010;
        
        h_t_prev[0] = 11'b11111111010;
        h_t_prev[1] = 11'b11111101100;
        h_t_prev[2] = 11'b11111011100;
        h_t_prev[3] = 11'b11111010001;
        h_t_prev[4] = 11'b11111010001;
        h_t_prev[5] = 11'b11111001101;
        h_t_prev[6] = 11'b11111011101;
        h_t_prev[7] = 11'b00000000111;
        h_t_prev[8] = 11'b11111100110;
        h_t_prev[9] = 11'b11111100010;
        h_t_prev[10] = 11'b11111011100;
        h_t_prev[11] = 11'b11111001010;
        h_t_prev[12] = 11'b11111010100;
        h_t_prev[13] = 11'b11111010000;
        h_t_prev[14] = 11'b11111111000;
        h_t_prev[15] = 11'b11111101000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 55 timeout!");
                $fdisplay(fd_cycles, "Test Vector  55: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  55: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 55");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 56
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111110111;
        x_t[1] = 11'b11111100111;
        x_t[2] = 11'b11111010110;
        x_t[3] = 11'b11111001110;
        x_t[4] = 11'b11111001101;
        x_t[5] = 11'b11111001010;
        x_t[6] = 11'b11111010011;
        x_t[7] = 11'b00000000001;
        x_t[8] = 11'b11111100000;
        x_t[9] = 11'b11111011011;
        x_t[10] = 11'b11111011000;
        x_t[11] = 11'b11111001001;
        x_t[12] = 11'b11111010000;
        x_t[13] = 11'b11111000000;
        x_t[14] = 11'b11111110010;
        x_t[15] = 11'b11111100011;
        x_t[16] = 11'b11111011100;
        x_t[17] = 11'b11111010100;
        x_t[18] = 11'b11111011000;
        x_t[19] = 11'b11111010100;
        x_t[20] = 11'b11111001101;
        x_t[21] = 11'b11111110000;
        x_t[22] = 11'b11111100011;
        x_t[23] = 11'b11111100010;
        x_t[24] = 11'b00000000100;
        x_t[25] = 11'b00000000100;
        x_t[26] = 11'b11111001110;
        x_t[27] = 11'b11111001101;
        x_t[28] = 11'b11111100001;
        x_t[29] = 11'b00000000100;
        x_t[30] = 11'b11111111011;
        x_t[31] = 11'b11111010001;
        x_t[32] = 11'b11111010001;
        x_t[33] = 11'b11111001001;
        x_t[34] = 11'b11111000111;
        x_t[35] = 11'b11111010011;
        x_t[36] = 11'b11111001110;
        x_t[37] = 11'b11111111010;
        x_t[38] = 11'b00000000001;
        x_t[39] = 11'b11111001011;
        x_t[40] = 11'b00000001001;
        x_t[41] = 11'b11111000100;
        x_t[42] = 11'b00000001100;
        x_t[43] = 11'b11111110101;
        x_t[44] = 11'b00000000101;
        x_t[45] = 11'b11111110010;
        x_t[46] = 11'b11111110101;
        x_t[47] = 11'b11111101010;
        x_t[48] = 11'b11111100010;
        x_t[49] = 11'b11111011110;
        x_t[50] = 11'b11111011100;
        x_t[51] = 11'b11111011011;
        x_t[52] = 11'b11111011111;
        x_t[53] = 11'b11111100111;
        x_t[54] = 11'b11111101001;
        x_t[55] = 11'b11111100011;
        x_t[56] = 11'b11111011100;
        x_t[57] = 11'b11111100110;
        x_t[58] = 11'b11111100001;
        x_t[59] = 11'b11111100110;
        x_t[60] = 11'b11111010111;
        x_t[61] = 11'b11111010001;
        x_t[62] = 11'b11111001011;
        x_t[63] = 11'b11111100011;
        
        h_t_prev[0] = 11'b11111110111;
        h_t_prev[1] = 11'b11111100111;
        h_t_prev[2] = 11'b11111010110;
        h_t_prev[3] = 11'b11111001110;
        h_t_prev[4] = 11'b11111001101;
        h_t_prev[5] = 11'b11111001010;
        h_t_prev[6] = 11'b11111010011;
        h_t_prev[7] = 11'b00000000001;
        h_t_prev[8] = 11'b11111100000;
        h_t_prev[9] = 11'b11111011011;
        h_t_prev[10] = 11'b11111011000;
        h_t_prev[11] = 11'b11111001001;
        h_t_prev[12] = 11'b11111010000;
        h_t_prev[13] = 11'b11111000000;
        h_t_prev[14] = 11'b11111110010;
        h_t_prev[15] = 11'b11111100011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 56 timeout!");
                $fdisplay(fd_cycles, "Test Vector  56: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  56: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 56");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 57
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111110110;
        x_t[1] = 11'b11111011111;
        x_t[2] = 11'b11111010000;
        x_t[3] = 11'b11111000111;
        x_t[4] = 11'b11111001000;
        x_t[5] = 11'b11111001010;
        x_t[6] = 11'b11111011001;
        x_t[7] = 11'b00000000000;
        x_t[8] = 11'b11111011010;
        x_t[9] = 11'b11111011000;
        x_t[10] = 11'b11111010101;
        x_t[11] = 11'b11111001001;
        x_t[12] = 11'b11111010010;
        x_t[13] = 11'b11111001100;
        x_t[14] = 11'b11111110001;
        x_t[15] = 11'b11111100100;
        x_t[16] = 11'b11111011100;
        x_t[17] = 11'b11111010101;
        x_t[18] = 11'b11111011011;
        x_t[19] = 11'b11111011001;
        x_t[20] = 11'b11111010011;
        x_t[21] = 11'b11111101100;
        x_t[22] = 11'b11111100001;
        x_t[23] = 11'b11111100000;
        x_t[24] = 11'b00000000001;
        x_t[25] = 11'b00000000000;
        x_t[26] = 11'b11111001100;
        x_t[27] = 11'b11111001100;
        x_t[28] = 11'b11111011111;
        x_t[29] = 11'b00000000011;
        x_t[30] = 11'b11111110110;
        x_t[31] = 11'b11111001111;
        x_t[32] = 11'b11111001101;
        x_t[33] = 11'b11111001000;
        x_t[34] = 11'b11111000111;
        x_t[35] = 11'b11111010010;
        x_t[36] = 11'b11111010011;
        x_t[37] = 11'b11111111001;
        x_t[38] = 11'b11111111011;
        x_t[39] = 11'b11111011001;
        x_t[40] = 11'b11111111101;
        x_t[41] = 11'b11111011111;
        x_t[42] = 11'b11111110101;
        x_t[43] = 11'b11111011101;
        x_t[44] = 11'b00000000010;
        x_t[45] = 11'b11111101001;
        x_t[46] = 11'b11111110011;
        x_t[47] = 11'b11111110000;
        x_t[48] = 11'b11111100111;
        x_t[49] = 11'b11111101001;
        x_t[50] = 11'b11111100011;
        x_t[51] = 11'b11111101100;
        x_t[52] = 11'b11111110000;
        x_t[53] = 11'b11111111011;
        x_t[54] = 11'b11111111100;
        x_t[55] = 11'b11111110000;
        x_t[56] = 11'b11111101010;
        x_t[57] = 11'b11111110101;
        x_t[58] = 11'b11111111111;
        x_t[59] = 11'b00000001100;
        x_t[60] = 11'b11111100100;
        x_t[61] = 11'b11111100110;
        x_t[62] = 11'b11111101001;
        x_t[63] = 11'b11111111001;
        
        h_t_prev[0] = 11'b11111110110;
        h_t_prev[1] = 11'b11111011111;
        h_t_prev[2] = 11'b11111010000;
        h_t_prev[3] = 11'b11111000111;
        h_t_prev[4] = 11'b11111001000;
        h_t_prev[5] = 11'b11111001010;
        h_t_prev[6] = 11'b11111011001;
        h_t_prev[7] = 11'b00000000000;
        h_t_prev[8] = 11'b11111011010;
        h_t_prev[9] = 11'b11111011000;
        h_t_prev[10] = 11'b11111010101;
        h_t_prev[11] = 11'b11111001001;
        h_t_prev[12] = 11'b11111010010;
        h_t_prev[13] = 11'b11111001100;
        h_t_prev[14] = 11'b11111110001;
        h_t_prev[15] = 11'b11111100100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 57 timeout!");
                $fdisplay(fd_cycles, "Test Vector  57: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  57: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 57");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 58
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111101111;
        x_t[1] = 11'b11111011011;
        x_t[2] = 11'b11111001101;
        x_t[3] = 11'b11111000011;
        x_t[4] = 11'b11111001000;
        x_t[5] = 11'b11111001001;
        x_t[6] = 11'b11111011000;
        x_t[7] = 11'b11111111011;
        x_t[8] = 11'b11111011010;
        x_t[9] = 11'b11111011000;
        x_t[10] = 11'b11111010111;
        x_t[11] = 11'b11111001011;
        x_t[12] = 11'b11111010101;
        x_t[13] = 11'b11111010000;
        x_t[14] = 11'b11111110000;
        x_t[15] = 11'b11111101000;
        x_t[16] = 11'b11111100010;
        x_t[17] = 11'b11111010111;
        x_t[18] = 11'b11111100011;
        x_t[19] = 11'b11111100001;
        x_t[20] = 11'b11111011010;
        x_t[21] = 11'b11111101010;
        x_t[22] = 11'b11111011100;
        x_t[23] = 11'b11111011011;
        x_t[24] = 11'b11111111011;
        x_t[25] = 11'b11111111011;
        x_t[26] = 11'b11111000101;
        x_t[27] = 11'b11111000101;
        x_t[28] = 11'b11111011001;
        x_t[29] = 11'b11111110111;
        x_t[30] = 11'b11111101110;
        x_t[31] = 11'b11111000111;
        x_t[32] = 11'b11111001000;
        x_t[33] = 11'b11111000010;
        x_t[34] = 11'b11111000010;
        x_t[35] = 11'b11111001011;
        x_t[36] = 11'b11111001010;
        x_t[37] = 11'b11111101110;
        x_t[38] = 11'b11111111010;
        x_t[39] = 11'b11111001011;
        x_t[40] = 11'b11111110011;
        x_t[41] = 11'b11110110111;
        x_t[42] = 11'b11111111000;
        x_t[43] = 11'b11111101010;
        x_t[44] = 11'b00000000001;
        x_t[45] = 11'b11111111010;
        x_t[46] = 11'b11111110010;
        x_t[47] = 11'b11111110101;
        x_t[48] = 11'b11111110000;
        x_t[49] = 11'b11111110010;
        x_t[50] = 11'b11111101010;
        x_t[51] = 11'b11111111101;
        x_t[52] = 11'b00000000010;
        x_t[53] = 11'b00000010010;
        x_t[54] = 11'b00000011001;
        x_t[55] = 11'b11111111110;
        x_t[56] = 11'b11111110111;
        x_t[57] = 11'b00000000011;
        x_t[58] = 11'b00000011111;
        x_t[59] = 11'b00000110100;
        x_t[60] = 11'b11111111001;
        x_t[61] = 11'b00000000111;
        x_t[62] = 11'b00000011000;
        x_t[63] = 11'b00000010100;
        
        h_t_prev[0] = 11'b11111101111;
        h_t_prev[1] = 11'b11111011011;
        h_t_prev[2] = 11'b11111001101;
        h_t_prev[3] = 11'b11111000011;
        h_t_prev[4] = 11'b11111001000;
        h_t_prev[5] = 11'b11111001001;
        h_t_prev[6] = 11'b11111011000;
        h_t_prev[7] = 11'b11111111011;
        h_t_prev[8] = 11'b11111011010;
        h_t_prev[9] = 11'b11111011000;
        h_t_prev[10] = 11'b11111010111;
        h_t_prev[11] = 11'b11111001011;
        h_t_prev[12] = 11'b11111010101;
        h_t_prev[13] = 11'b11111010000;
        h_t_prev[14] = 11'b11111110000;
        h_t_prev[15] = 11'b11111101000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 58 timeout!");
                $fdisplay(fd_cycles, "Test Vector  58: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  58: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 58");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 59
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111101110;
        x_t[1] = 11'b11111100000;
        x_t[2] = 11'b11111001101;
        x_t[3] = 11'b11111000011;
        x_t[4] = 11'b11111000110;
        x_t[5] = 11'b11111000101;
        x_t[6] = 11'b11111001101;
        x_t[7] = 11'b11111111010;
        x_t[8] = 11'b11111011111;
        x_t[9] = 11'b11111011011;
        x_t[10] = 11'b11111011010;
        x_t[11] = 11'b11111001110;
        x_t[12] = 11'b11111010011;
        x_t[13] = 11'b11111000101;
        x_t[14] = 11'b11111110100;
        x_t[15] = 11'b11111101100;
        x_t[16] = 11'b11111100111;
        x_t[17] = 11'b11111011010;
        x_t[18] = 11'b11111100111;
        x_t[19] = 11'b11111100111;
        x_t[20] = 11'b11111100000;
        x_t[21] = 11'b11111101111;
        x_t[22] = 11'b11111100001;
        x_t[23] = 11'b11111100001;
        x_t[24] = 11'b00000000001;
        x_t[25] = 11'b00000000000;
        x_t[26] = 11'b11111001101;
        x_t[27] = 11'b11111001011;
        x_t[28] = 11'b11111011101;
        x_t[29] = 11'b00000000000;
        x_t[30] = 11'b11111110101;
        x_t[31] = 11'b11111010000;
        x_t[32] = 11'b11111010001;
        x_t[33] = 11'b11111000111;
        x_t[34] = 11'b11111000110;
        x_t[35] = 11'b11111010010;
        x_t[36] = 11'b11111001010;
        x_t[37] = 11'b11111101011;
        x_t[38] = 11'b00000000100;
        x_t[39] = 11'b11111000110;
        x_t[40] = 11'b00000000101;
        x_t[41] = 11'b11110111000;
        x_t[42] = 11'b00000010101;
        x_t[43] = 11'b11111100001;
        x_t[44] = 11'b00000010101;
        x_t[45] = 11'b00000010000;
        x_t[46] = 11'b00000000011;
        x_t[47] = 11'b00000000001;
        x_t[48] = 11'b11111111001;
        x_t[49] = 11'b11111110100;
        x_t[50] = 11'b11111101011;
        x_t[51] = 11'b00000000001;
        x_t[52] = 11'b00000001010;
        x_t[53] = 11'b00000011110;
        x_t[54] = 11'b00000101000;
        x_t[55] = 11'b00000001111;
        x_t[56] = 11'b00000000010;
        x_t[57] = 11'b00000000011;
        x_t[58] = 11'b00000101001;
        x_t[59] = 11'b00001000100;
        x_t[60] = 11'b00000001110;
        x_t[61] = 11'b00000100000;
        x_t[62] = 11'b00000111101;
        x_t[63] = 11'b00000101001;
        
        h_t_prev[0] = 11'b11111101110;
        h_t_prev[1] = 11'b11111100000;
        h_t_prev[2] = 11'b11111001101;
        h_t_prev[3] = 11'b11111000011;
        h_t_prev[4] = 11'b11111000110;
        h_t_prev[5] = 11'b11111000101;
        h_t_prev[6] = 11'b11111001101;
        h_t_prev[7] = 11'b11111111010;
        h_t_prev[8] = 11'b11111011111;
        h_t_prev[9] = 11'b11111011011;
        h_t_prev[10] = 11'b11111011010;
        h_t_prev[11] = 11'b11111001110;
        h_t_prev[12] = 11'b11111010011;
        h_t_prev[13] = 11'b11111000101;
        h_t_prev[14] = 11'b11111110100;
        h_t_prev[15] = 11'b11111101100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 59 timeout!");
                $fdisplay(fd_cycles, "Test Vector  59: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  59: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 59");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 60
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111111101;
        x_t[1] = 11'b11111110000;
        x_t[2] = 11'b11111011010;
        x_t[3] = 11'b11111001111;
        x_t[4] = 11'b11111001011;
        x_t[5] = 11'b11111001001;
        x_t[6] = 11'b11111010010;
        x_t[7] = 11'b00000001000;
        x_t[8] = 11'b11111101010;
        x_t[9] = 11'b11111100010;
        x_t[10] = 11'b11111011111;
        x_t[11] = 11'b11111010001;
        x_t[12] = 11'b11111011001;
        x_t[13] = 11'b11111001111;
        x_t[14] = 11'b00000000000;
        x_t[15] = 11'b11111110000;
        x_t[16] = 11'b11111101001;
        x_t[17] = 11'b11111011101;
        x_t[18] = 11'b11111101001;
        x_t[19] = 11'b11111101100;
        x_t[20] = 11'b11111101010;
        x_t[21] = 11'b11111110001;
        x_t[22] = 11'b11111100000;
        x_t[23] = 11'b11111011111;
        x_t[24] = 11'b00000000100;
        x_t[25] = 11'b00000000010;
        x_t[26] = 11'b11111010000;
        x_t[27] = 11'b11111001000;
        x_t[28] = 11'b11111011000;
        x_t[29] = 11'b00000000101;
        x_t[30] = 11'b11111111011;
        x_t[31] = 11'b11111001110;
        x_t[32] = 11'b11111010111;
        x_t[33] = 11'b11111001100;
        x_t[34] = 11'b11111000110;
        x_t[35] = 11'b11111010010;
        x_t[36] = 11'b11111000100;
        x_t[37] = 11'b11111101000;
        x_t[38] = 11'b00000000110;
        x_t[39] = 11'b11111000111;
        x_t[40] = 11'b00000010011;
        x_t[41] = 11'b11111001001;
        x_t[42] = 11'b00000010010;
        x_t[43] = 11'b11111011111;
        x_t[44] = 11'b00000010110;
        x_t[45] = 11'b11111111100;
        x_t[46] = 11'b00000001010;
        x_t[47] = 11'b00000000011;
        x_t[48] = 11'b11111111000;
        x_t[49] = 11'b11111110010;
        x_t[50] = 11'b11111101000;
        x_t[51] = 11'b00000000001;
        x_t[52] = 11'b00000001011;
        x_t[53] = 11'b00000011110;
        x_t[54] = 11'b00000100101;
        x_t[55] = 11'b00000010101;
        x_t[56] = 11'b00000000100;
        x_t[57] = 11'b00000000010;
        x_t[58] = 11'b00000101011;
        x_t[59] = 11'b00001000111;
        x_t[60] = 11'b00000011011;
        x_t[61] = 11'b00000100111;
        x_t[62] = 11'b00001001010;
        x_t[63] = 11'b00000101011;
        
        h_t_prev[0] = 11'b11111111101;
        h_t_prev[1] = 11'b11111110000;
        h_t_prev[2] = 11'b11111011010;
        h_t_prev[3] = 11'b11111001111;
        h_t_prev[4] = 11'b11111001011;
        h_t_prev[5] = 11'b11111001001;
        h_t_prev[6] = 11'b11111010010;
        h_t_prev[7] = 11'b00000001000;
        h_t_prev[8] = 11'b11111101010;
        h_t_prev[9] = 11'b11111100010;
        h_t_prev[10] = 11'b11111011111;
        h_t_prev[11] = 11'b11111010001;
        h_t_prev[12] = 11'b11111011001;
        h_t_prev[13] = 11'b11111001111;
        h_t_prev[14] = 11'b00000000000;
        h_t_prev[15] = 11'b11111110000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 60 timeout!");
                $fdisplay(fd_cycles, "Test Vector  60: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  60: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 60");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 61
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111111101;
        x_t[1] = 11'b11111101011;
        x_t[2] = 11'b11111010111;
        x_t[3] = 11'b11111001010;
        x_t[4] = 11'b11111000101;
        x_t[5] = 11'b11111000010;
        x_t[6] = 11'b11111001000;
        x_t[7] = 11'b00000000110;
        x_t[8] = 11'b11111100110;
        x_t[9] = 11'b11111100000;
        x_t[10] = 11'b11111011111;
        x_t[11] = 11'b11111001101;
        x_t[12] = 11'b11111010111;
        x_t[13] = 11'b11111010000;
        x_t[14] = 11'b00000000001;
        x_t[15] = 11'b11111101101;
        x_t[16] = 11'b11111101000;
        x_t[17] = 11'b11111011111;
        x_t[18] = 11'b11111101101;
        x_t[19] = 11'b11111110000;
        x_t[20] = 11'b11111110000;
        x_t[21] = 11'b11111101000;
        x_t[22] = 11'b11111010110;
        x_t[23] = 11'b11111010100;
        x_t[24] = 11'b11111111101;
        x_t[25] = 11'b11111111011;
        x_t[26] = 11'b11111000101;
        x_t[27] = 11'b11110111011;
        x_t[28] = 11'b11111001110;
        x_t[29] = 11'b00000001010;
        x_t[30] = 11'b11111110010;
        x_t[31] = 11'b11111000111;
        x_t[32] = 11'b11111001111;
        x_t[33] = 11'b11111000011;
        x_t[34] = 11'b11110111011;
        x_t[35] = 11'b11111000110;
        x_t[36] = 11'b11110111100;
        x_t[37] = 11'b11111100111;
        x_t[38] = 11'b00000001100;
        x_t[39] = 11'b11110111111;
        x_t[40] = 11'b00000010101;
        x_t[41] = 11'b11111000110;
        x_t[42] = 11'b00000001110;
        x_t[43] = 11'b00000010000;
        x_t[44] = 11'b00000100000;
        x_t[45] = 11'b00000001110;
        x_t[46] = 11'b00000011011;
        x_t[47] = 11'b00000010010;
        x_t[48] = 11'b00000000100;
        x_t[49] = 11'b11111111111;
        x_t[50] = 11'b11111110110;
        x_t[51] = 11'b00000001111;
        x_t[52] = 11'b00000011000;
        x_t[53] = 11'b00000101100;
        x_t[54] = 11'b00000110011;
        x_t[55] = 11'b00000101001;
        x_t[56] = 11'b00000010110;
        x_t[57] = 11'b00000001111;
        x_t[58] = 11'b00000110101;
        x_t[59] = 11'b00001001011;
        x_t[60] = 11'b00000100110;
        x_t[61] = 11'b00000101000;
        x_t[62] = 11'b00001001001;
        x_t[63] = 11'b00000101101;
        
        h_t_prev[0] = 11'b11111111101;
        h_t_prev[1] = 11'b11111101011;
        h_t_prev[2] = 11'b11111010111;
        h_t_prev[3] = 11'b11111001010;
        h_t_prev[4] = 11'b11111000101;
        h_t_prev[5] = 11'b11111000010;
        h_t_prev[6] = 11'b11111001000;
        h_t_prev[7] = 11'b00000000110;
        h_t_prev[8] = 11'b11111100110;
        h_t_prev[9] = 11'b11111100000;
        h_t_prev[10] = 11'b11111011111;
        h_t_prev[11] = 11'b11111001101;
        h_t_prev[12] = 11'b11111010111;
        h_t_prev[13] = 11'b11111010000;
        h_t_prev[14] = 11'b00000000001;
        h_t_prev[15] = 11'b11111101101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 61 timeout!");
                $fdisplay(fd_cycles, "Test Vector  61: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  61: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 61");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 62
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000000101;
        x_t[1] = 11'b11111110010;
        x_t[2] = 11'b11111011100;
        x_t[3] = 11'b11111000110;
        x_t[4] = 11'b11111000100;
        x_t[5] = 11'b11111000010;
        x_t[6] = 11'b11111001111;
        x_t[7] = 11'b00000010101;
        x_t[8] = 11'b11111110011;
        x_t[9] = 11'b11111101101;
        x_t[10] = 11'b11111101010;
        x_t[11] = 11'b11111010100;
        x_t[12] = 11'b11111011011;
        x_t[13] = 11'b11111011101;
        x_t[14] = 11'b00000010011;
        x_t[15] = 11'b00000000010;
        x_t[16] = 11'b11111111010;
        x_t[17] = 11'b11111101110;
        x_t[18] = 11'b11111111010;
        x_t[19] = 11'b11111111100;
        x_t[20] = 11'b11111111110;
        x_t[21] = 11'b11111101011;
        x_t[22] = 11'b11111011000;
        x_t[23] = 11'b11111011000;
        x_t[24] = 11'b11111111111;
        x_t[25] = 11'b11111111101;
        x_t[26] = 11'b11111000110;
        x_t[27] = 11'b11110111100;
        x_t[28] = 11'b11111010011;
        x_t[29] = 11'b00000001001;
        x_t[30] = 11'b11111110110;
        x_t[31] = 11'b11111000111;
        x_t[32] = 11'b11111010010;
        x_t[33] = 11'b11111000010;
        x_t[34] = 11'b11110111010;
        x_t[35] = 11'b11111000110;
        x_t[36] = 11'b11111000000;
        x_t[37] = 11'b11111110000;
        x_t[38] = 11'b00000010001;
        x_t[39] = 11'b11111001001;
        x_t[40] = 11'b00000001111;
        x_t[41] = 11'b11111001001;
        x_t[42] = 11'b00000100100;
        x_t[43] = 11'b11111110110;
        x_t[44] = 11'b00000110110;
        x_t[45] = 11'b00000011011;
        x_t[46] = 11'b00000110101;
        x_t[47] = 11'b00000100010;
        x_t[48] = 11'b00000001111;
        x_t[49] = 11'b00000001010;
        x_t[50] = 11'b11111111111;
        x_t[51] = 11'b00000010001;
        x_t[52] = 11'b00000010110;
        x_t[53] = 11'b00000101000;
        x_t[54] = 11'b00000101110;
        x_t[55] = 11'b00000111000;
        x_t[56] = 11'b00000100001;
        x_t[57] = 11'b00000010101;
        x_t[58] = 11'b00000101111;
        x_t[59] = 11'b00001000001;
        x_t[60] = 11'b00000110010;
        x_t[61] = 11'b00000101011;
        x_t[62] = 11'b00001000011;
        x_t[63] = 11'b00000111000;
        
        h_t_prev[0] = 11'b00000000101;
        h_t_prev[1] = 11'b11111110010;
        h_t_prev[2] = 11'b11111011100;
        h_t_prev[3] = 11'b11111000110;
        h_t_prev[4] = 11'b11111000100;
        h_t_prev[5] = 11'b11111000010;
        h_t_prev[6] = 11'b11111001111;
        h_t_prev[7] = 11'b00000010101;
        h_t_prev[8] = 11'b11111110011;
        h_t_prev[9] = 11'b11111101101;
        h_t_prev[10] = 11'b11111101010;
        h_t_prev[11] = 11'b11111010100;
        h_t_prev[12] = 11'b11111011011;
        h_t_prev[13] = 11'b11111011101;
        h_t_prev[14] = 11'b00000010011;
        h_t_prev[15] = 11'b00000000010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 62 timeout!");
                $fdisplay(fd_cycles, "Test Vector  62: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  62: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 62");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 63
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000000001;
        x_t[1] = 11'b11111110111;
        x_t[2] = 11'b11111100001;
        x_t[3] = 11'b11111001011;
        x_t[4] = 11'b11111000001;
        x_t[5] = 11'b11110111010;
        x_t[6] = 11'b11111001010;
        x_t[7] = 11'b00000010100;
        x_t[8] = 11'b11111110101;
        x_t[9] = 11'b11111110010;
        x_t[10] = 11'b11111101011;
        x_t[11] = 11'b11111001100;
        x_t[12] = 11'b11111001011;
        x_t[13] = 11'b11111010000;
        x_t[14] = 11'b00000011100;
        x_t[15] = 11'b00000000101;
        x_t[16] = 11'b11111111100;
        x_t[17] = 11'b11111101111;
        x_t[18] = 11'b11111110101;
        x_t[19] = 11'b11111110001;
        x_t[20] = 11'b11111101101;
        x_t[21] = 11'b11111101111;
        x_t[22] = 11'b11111011100;
        x_t[23] = 11'b11111011011;
        x_t[24] = 11'b00000000100;
        x_t[25] = 11'b00000000010;
        x_t[26] = 11'b11111001010;
        x_t[27] = 11'b11110111110;
        x_t[28] = 11'b11111001111;
        x_t[29] = 11'b00000001111;
        x_t[30] = 11'b11111111010;
        x_t[31] = 11'b11111001010;
        x_t[32] = 11'b11111011001;
        x_t[33] = 11'b11111001010;
        x_t[34] = 11'b11111000000;
        x_t[35] = 11'b11111001011;
        x_t[36] = 11'b11111000001;
        x_t[37] = 11'b11111110000;
        x_t[38] = 11'b00000010010;
        x_t[39] = 11'b11111001010;
        x_t[40] = 11'b00000011011;
        x_t[41] = 11'b11111011100;
        x_t[42] = 11'b00000101100;
        x_t[43] = 11'b11111101011;
        x_t[44] = 11'b00000110110;
        x_t[45] = 11'b00000000101;
        x_t[46] = 11'b00000110000;
        x_t[47] = 11'b00000100001;
        x_t[48] = 11'b00000001101;
        x_t[49] = 11'b00000001001;
        x_t[50] = 11'b11111111011;
        x_t[51] = 11'b00000000111;
        x_t[52] = 11'b00000001011;
        x_t[53] = 11'b00000010111;
        x_t[54] = 11'b00000011100;
        x_t[55] = 11'b00000110111;
        x_t[56] = 11'b00000100000;
        x_t[57] = 11'b00000010001;
        x_t[58] = 11'b00000011110;
        x_t[59] = 11'b00000100011;
        x_t[60] = 11'b00000110110;
        x_t[61] = 11'b00000100011;
        x_t[62] = 11'b00000110100;
        x_t[63] = 11'b00000110100;
        
        h_t_prev[0] = 11'b00000000001;
        h_t_prev[1] = 11'b11111110111;
        h_t_prev[2] = 11'b11111100001;
        h_t_prev[3] = 11'b11111001011;
        h_t_prev[4] = 11'b11111000001;
        h_t_prev[5] = 11'b11110111010;
        h_t_prev[6] = 11'b11111001010;
        h_t_prev[7] = 11'b00000010100;
        h_t_prev[8] = 11'b11111110101;
        h_t_prev[9] = 11'b11111110010;
        h_t_prev[10] = 11'b11111101011;
        h_t_prev[11] = 11'b11111001100;
        h_t_prev[12] = 11'b11111001011;
        h_t_prev[13] = 11'b11111010000;
        h_t_prev[14] = 11'b00000011100;
        h_t_prev[15] = 11'b00000000101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 63 timeout!");
                $fdisplay(fd_cycles, "Test Vector  63: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  63: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 63");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 64
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000000111;
        x_t[1] = 11'b11111111011;
        x_t[2] = 11'b11111100100;
        x_t[3] = 11'b11111001111;
        x_t[4] = 11'b11111000111;
        x_t[5] = 11'b11110111101;
        x_t[6] = 11'b11111001011;
        x_t[7] = 11'b00000010111;
        x_t[8] = 11'b11111110110;
        x_t[9] = 11'b11111110001;
        x_t[10] = 11'b11111100101;
        x_t[11] = 11'b11111001100;
        x_t[12] = 11'b11111000111;
        x_t[13] = 11'b11111010000;
        x_t[14] = 11'b00000010111;
        x_t[15] = 11'b00000000011;
        x_t[16] = 11'b11111111001;
        x_t[17] = 11'b11111101101;
        x_t[18] = 11'b11111110001;
        x_t[19] = 11'b11111101001;
        x_t[20] = 11'b11111100101;
        x_t[21] = 11'b11111110101;
        x_t[22] = 11'b11111100011;
        x_t[23] = 11'b11111100011;
        x_t[24] = 11'b00000001000;
        x_t[25] = 11'b00000000111;
        x_t[26] = 11'b11111010001;
        x_t[27] = 11'b11111000111;
        x_t[28] = 11'b11111011101;
        x_t[29] = 11'b00000010100;
        x_t[30] = 11'b11111111011;
        x_t[31] = 11'b11111010100;
        x_t[32] = 11'b11111011010;
        x_t[33] = 11'b11111001101;
        x_t[34] = 11'b11111000111;
        x_t[35] = 11'b11111010000;
        x_t[36] = 11'b11111000111;
        x_t[37] = 11'b11111110100;
        x_t[38] = 11'b00000011000;
        x_t[39] = 11'b11111010101;
        x_t[40] = 11'b00000101010;
        x_t[41] = 11'b11111101011;
        x_t[42] = 11'b00000101110;
        x_t[43] = 11'b11111100100;
        x_t[44] = 11'b00000110110;
        x_t[45] = 11'b11111111110;
        x_t[46] = 11'b00000101010;
        x_t[47] = 11'b00000011011;
        x_t[48] = 11'b00000001010;
        x_t[49] = 11'b00000001000;
        x_t[50] = 11'b11111111101;
        x_t[51] = 11'b00000000101;
        x_t[52] = 11'b00000000110;
        x_t[53] = 11'b00000001100;
        x_t[54] = 11'b00000001101;
        x_t[55] = 11'b00000110000;
        x_t[56] = 11'b00000011011;
        x_t[57] = 11'b00000010000;
        x_t[58] = 11'b00000010110;
        x_t[59] = 11'b00000010001;
        x_t[60] = 11'b00000101111;
        x_t[61] = 11'b00000010110;
        x_t[62] = 11'b00000100010;
        x_t[63] = 11'b00000101011;
        
        h_t_prev[0] = 11'b00000000111;
        h_t_prev[1] = 11'b11111111011;
        h_t_prev[2] = 11'b11111100100;
        h_t_prev[3] = 11'b11111001111;
        h_t_prev[4] = 11'b11111000111;
        h_t_prev[5] = 11'b11110111101;
        h_t_prev[6] = 11'b11111001011;
        h_t_prev[7] = 11'b00000010111;
        h_t_prev[8] = 11'b11111110110;
        h_t_prev[9] = 11'b11111110001;
        h_t_prev[10] = 11'b11111100101;
        h_t_prev[11] = 11'b11111001100;
        h_t_prev[12] = 11'b11111000111;
        h_t_prev[13] = 11'b11111010000;
        h_t_prev[14] = 11'b00000010111;
        h_t_prev[15] = 11'b00000000011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 64 timeout!");
                $fdisplay(fd_cycles, "Test Vector  64: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  64: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 64");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 65
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111001010;
        x_t[1] = 11'b11111011110;
        x_t[2] = 11'b11111100001;
        x_t[3] = 11'b11111110101;
        x_t[4] = 11'b11111111001;
        x_t[5] = 11'b11111111000;
        x_t[6] = 11'b11111101000;
        x_t[7] = 11'b11111011011;
        x_t[8] = 11'b11111101100;
        x_t[9] = 11'b11111110011;
        x_t[10] = 11'b11111111011;
        x_t[11] = 11'b00000000000;
        x_t[12] = 11'b00000000011;
        x_t[13] = 11'b11111111001;
        x_t[14] = 11'b11111101100;
        x_t[15] = 11'b11111110100;
        x_t[16] = 11'b11111111000;
        x_t[17] = 11'b00000000100;
        x_t[18] = 11'b00000000101;
        x_t[19] = 11'b00000001001;
        x_t[20] = 11'b00000001100;
        x_t[21] = 11'b11111001100;
        x_t[22] = 11'b11111001001;
        x_t[23] = 11'b11111010010;
        x_t[24] = 11'b11111001000;
        x_t[25] = 11'b11111001001;
        x_t[26] = 11'b11111010110;
        x_t[27] = 11'b11111011001;
        x_t[28] = 11'b11111010110;
        x_t[29] = 11'b11111000101;
        x_t[30] = 11'b11111010011;
        x_t[31] = 11'b11111011011;
        x_t[32] = 11'b11111011101;
        x_t[33] = 11'b11111100011;
        x_t[34] = 11'b11111101010;
        x_t[35] = 11'b11111101001;
        x_t[36] = 11'b11111101000;
        x_t[37] = 11'b11111101010;
        x_t[38] = 11'b11111001010;
        x_t[39] = 11'b11111101011;
        x_t[40] = 11'b11111001110;
        x_t[41] = 11'b00000000000;
        x_t[42] = 11'b11110111110;
        x_t[43] = 11'b00000000110;
        x_t[44] = 11'b11111100001;
        x_t[45] = 11'b11111111100;
        x_t[46] = 11'b11111111101;
        x_t[47] = 11'b11111111100;
        x_t[48] = 11'b00000000011;
        x_t[49] = 11'b00000000101;
        x_t[50] = 11'b00000000110;
        x_t[51] = 11'b00000010010;
        x_t[52] = 11'b00000001011;
        x_t[53] = 11'b00000010001;
        x_t[54] = 11'b00000001011;
        x_t[55] = 11'b00000001101;
        x_t[56] = 11'b00000001101;
        x_t[57] = 11'b00000011100;
        x_t[58] = 11'b00000011100;
        x_t[59] = 11'b00000010110;
        x_t[60] = 11'b00000011101;
        x_t[61] = 11'b00000100111;
        x_t[62] = 11'b00000001011;
        x_t[63] = 11'b00000011010;
        
        h_t_prev[0] = 11'b11111001010;
        h_t_prev[1] = 11'b11111011110;
        h_t_prev[2] = 11'b11111100001;
        h_t_prev[3] = 11'b11111110101;
        h_t_prev[4] = 11'b11111111001;
        h_t_prev[5] = 11'b11111111000;
        h_t_prev[6] = 11'b11111101000;
        h_t_prev[7] = 11'b11111011011;
        h_t_prev[8] = 11'b11111101100;
        h_t_prev[9] = 11'b11111110011;
        h_t_prev[10] = 11'b11111111011;
        h_t_prev[11] = 11'b00000000000;
        h_t_prev[12] = 11'b00000000011;
        h_t_prev[13] = 11'b11111111001;
        h_t_prev[14] = 11'b11111101100;
        h_t_prev[15] = 11'b11111110100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 65 timeout!");
                $fdisplay(fd_cycles, "Test Vector  65: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  65: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 65");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 66
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111001110;
        x_t[1] = 11'b11111100100;
        x_t[2] = 11'b11111100111;
        x_t[3] = 11'b11111110101;
        x_t[4] = 11'b11111111011;
        x_t[5] = 11'b11111111110;
        x_t[6] = 11'b11111111000;
        x_t[7] = 11'b11111100010;
        x_t[8] = 11'b11111110001;
        x_t[9] = 11'b11111110100;
        x_t[10] = 11'b11111110110;
        x_t[11] = 11'b11111111111;
        x_t[12] = 11'b00000000101;
        x_t[13] = 11'b00000000101;
        x_t[14] = 11'b11111101011;
        x_t[15] = 11'b11111110011;
        x_t[16] = 11'b11111110110;
        x_t[17] = 11'b11111111100;
        x_t[18] = 11'b11111111000;
        x_t[19] = 11'b11111111111;
        x_t[20] = 11'b00000000101;
        x_t[21] = 11'b11111001001;
        x_t[22] = 11'b11111001100;
        x_t[23] = 11'b11111010111;
        x_t[24] = 11'b11111000111;
        x_t[25] = 11'b11111001000;
        x_t[26] = 11'b11111010111;
        x_t[27] = 11'b11111011111;
        x_t[28] = 11'b11111011101;
        x_t[29] = 11'b11111000111;
        x_t[30] = 11'b11111011001;
        x_t[31] = 11'b11111011111;
        x_t[32] = 11'b11111011101;
        x_t[33] = 11'b11111100100;
        x_t[34] = 11'b11111101100;
        x_t[35] = 11'b11111101011;
        x_t[36] = 11'b11111110010;
        x_t[37] = 11'b11111110000;
        x_t[38] = 11'b11111001100;
        x_t[39] = 11'b11111111100;
        x_t[40] = 11'b11111010000;
        x_t[41] = 11'b00000101001;
        x_t[42] = 11'b11110111111;
        x_t[43] = 11'b11111011111;
        x_t[44] = 11'b11111011000;
        x_t[45] = 11'b11111101011;
        x_t[46] = 11'b11111110011;
        x_t[47] = 11'b11111111001;
        x_t[48] = 11'b00000000011;
        x_t[49] = 11'b00000000001;
        x_t[50] = 11'b11111111110;
        x_t[51] = 11'b00000001000;
        x_t[52] = 11'b00000000010;
        x_t[53] = 11'b00000001011;
        x_t[54] = 11'b00000000110;
        x_t[55] = 11'b00000001100;
        x_t[56] = 11'b00000001011;
        x_t[57] = 11'b00000011001;
        x_t[58] = 11'b00000011000;
        x_t[59] = 11'b00000010101;
        x_t[60] = 11'b00000011001;
        x_t[61] = 11'b00000100011;
        x_t[62] = 11'b00000000101;
        x_t[63] = 11'b00000010111;
        
        h_t_prev[0] = 11'b11111001110;
        h_t_prev[1] = 11'b11111100100;
        h_t_prev[2] = 11'b11111100111;
        h_t_prev[3] = 11'b11111110101;
        h_t_prev[4] = 11'b11111111011;
        h_t_prev[5] = 11'b11111111110;
        h_t_prev[6] = 11'b11111111000;
        h_t_prev[7] = 11'b11111100010;
        h_t_prev[8] = 11'b11111110001;
        h_t_prev[9] = 11'b11111110100;
        h_t_prev[10] = 11'b11111110110;
        h_t_prev[11] = 11'b11111111111;
        h_t_prev[12] = 11'b00000000101;
        h_t_prev[13] = 11'b00000000101;
        h_t_prev[14] = 11'b11111101011;
        h_t_prev[15] = 11'b11111110011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 66 timeout!");
                $fdisplay(fd_cycles, "Test Vector  66: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  66: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 66");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 67
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111010101;
        x_t[1] = 11'b11111101011;
        x_t[2] = 11'b11111101011;
        x_t[3] = 11'b11111110100;
        x_t[4] = 11'b11111111001;
        x_t[5] = 11'b11111111110;
        x_t[6] = 11'b00000000000;
        x_t[7] = 11'b11111101011;
        x_t[8] = 11'b11111110111;
        x_t[9] = 11'b11111110010;
        x_t[10] = 11'b11111101111;
        x_t[11] = 11'b11111111000;
        x_t[12] = 11'b00000000010;
        x_t[13] = 11'b00000001010;
        x_t[14] = 11'b11111110000;
        x_t[15] = 11'b11111110111;
        x_t[16] = 11'b11111110100;
        x_t[17] = 11'b11111111000;
        x_t[18] = 11'b11111110000;
        x_t[19] = 11'b11111111000;
        x_t[20] = 11'b00000000110;
        x_t[21] = 11'b11111010001;
        x_t[22] = 11'b11111010001;
        x_t[23] = 11'b11111011010;
        x_t[24] = 11'b11111001111;
        x_t[25] = 11'b11111001111;
        x_t[26] = 11'b11111011011;
        x_t[27] = 11'b11111100001;
        x_t[28] = 11'b11111011101;
        x_t[29] = 11'b11111010001;
        x_t[30] = 11'b11111011010;
        x_t[31] = 11'b11111100011;
        x_t[32] = 11'b11111100011;
        x_t[33] = 11'b11111100111;
        x_t[34] = 11'b11111101110;
        x_t[35] = 11'b11111101110;
        x_t[36] = 11'b11111110010;
        x_t[37] = 11'b11111101110;
        x_t[38] = 11'b11111011011;
        x_t[39] = 11'b11111111000;
        x_t[40] = 11'b11111100000;
        x_t[41] = 11'b00000010011;
        x_t[42] = 11'b11110111100;
        x_t[43] = 11'b00000000110;
        x_t[44] = 11'b11111100100;
        x_t[45] = 11'b11111111000;
        x_t[46] = 11'b11111111111;
        x_t[47] = 11'b00000000001;
        x_t[48] = 11'b00000001001;
        x_t[49] = 11'b00000000100;
        x_t[50] = 11'b11111111111;
        x_t[51] = 11'b00000000101;
        x_t[52] = 11'b00000000000;
        x_t[53] = 11'b00000001110;
        x_t[54] = 11'b00000010000;
        x_t[55] = 11'b00000001110;
        x_t[56] = 11'b00000001101;
        x_t[57] = 11'b00000011001;
        x_t[58] = 11'b00000011011;
        x_t[59] = 11'b00000011001;
        x_t[60] = 11'b00000010111;
        x_t[61] = 11'b00000100001;
        x_t[62] = 11'b00000000101;
        x_t[63] = 11'b00000011000;
        
        h_t_prev[0] = 11'b11111010101;
        h_t_prev[1] = 11'b11111101011;
        h_t_prev[2] = 11'b11111101011;
        h_t_prev[3] = 11'b11111110100;
        h_t_prev[4] = 11'b11111111001;
        h_t_prev[5] = 11'b11111111110;
        h_t_prev[6] = 11'b00000000000;
        h_t_prev[7] = 11'b11111101011;
        h_t_prev[8] = 11'b11111110111;
        h_t_prev[9] = 11'b11111110010;
        h_t_prev[10] = 11'b11111101111;
        h_t_prev[11] = 11'b11111111000;
        h_t_prev[12] = 11'b00000000010;
        h_t_prev[13] = 11'b00000001010;
        h_t_prev[14] = 11'b11111110000;
        h_t_prev[15] = 11'b11111110111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 67 timeout!");
                $fdisplay(fd_cycles, "Test Vector  67: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  67: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 67");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 68
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111100010;
        x_t[1] = 11'b11111110010;
        x_t[2] = 11'b11111101111;
        x_t[3] = 11'b11111110101;
        x_t[4] = 11'b11111111000;
        x_t[5] = 11'b11111111010;
        x_t[6] = 11'b11111111000;
        x_t[7] = 11'b11111110101;
        x_t[8] = 11'b11111111011;
        x_t[9] = 11'b11111110101;
        x_t[10] = 11'b11111110100;
        x_t[11] = 11'b11111110100;
        x_t[12] = 11'b11111111000;
        x_t[13] = 11'b11111110011;
        x_t[14] = 11'b11111111001;
        x_t[15] = 11'b11111111010;
        x_t[16] = 11'b11111111000;
        x_t[17] = 11'b11111111000;
        x_t[18] = 11'b11111101011;
        x_t[19] = 11'b11111101111;
        x_t[20] = 11'b11111111000;
        x_t[21] = 11'b11111010001;
        x_t[22] = 11'b11111010000;
        x_t[23] = 11'b11111011001;
        x_t[24] = 11'b11111010000;
        x_t[25] = 11'b11111010001;
        x_t[26] = 11'b11111011100;
        x_t[27] = 11'b11111100001;
        x_t[28] = 11'b11111011101;
        x_t[29] = 11'b11111010100;
        x_t[30] = 11'b11111011111;
        x_t[31] = 11'b11111100010;
        x_t[32] = 11'b11111100100;
        x_t[33] = 11'b11111100111;
        x_t[34] = 11'b11111101111;
        x_t[35] = 11'b11111110000;
        x_t[36] = 11'b11111101100;
        x_t[37] = 11'b11111101101;
        x_t[38] = 11'b11111011000;
        x_t[39] = 11'b11111100101;
        x_t[40] = 11'b11111010111;
        x_t[41] = 11'b11111010000;
        x_t[42] = 11'b11111000100;
        x_t[43] = 11'b11111100111;
        x_t[44] = 11'b11111100001;
        x_t[45] = 11'b11111101100;
        x_t[46] = 11'b11111110110;
        x_t[47] = 11'b11111110110;
        x_t[48] = 11'b11111111101;
        x_t[49] = 11'b11111111011;
        x_t[50] = 11'b11111111100;
        x_t[51] = 11'b11111111110;
        x_t[52] = 11'b11111111001;
        x_t[53] = 11'b00000000010;
        x_t[54] = 11'b00000000011;
        x_t[55] = 11'b11111111001;
        x_t[56] = 11'b11111111011;
        x_t[57] = 11'b00000001110;
        x_t[58] = 11'b00000001110;
        x_t[59] = 11'b00000001101;
        x_t[60] = 11'b00000001100;
        x_t[61] = 11'b00000010111;
        x_t[62] = 11'b11111111110;
        x_t[63] = 11'b00000001100;
        
        h_t_prev[0] = 11'b11111100010;
        h_t_prev[1] = 11'b11111110010;
        h_t_prev[2] = 11'b11111101111;
        h_t_prev[3] = 11'b11111110101;
        h_t_prev[4] = 11'b11111111000;
        h_t_prev[5] = 11'b11111111010;
        h_t_prev[6] = 11'b11111111000;
        h_t_prev[7] = 11'b11111110101;
        h_t_prev[8] = 11'b11111111011;
        h_t_prev[9] = 11'b11111110101;
        h_t_prev[10] = 11'b11111110100;
        h_t_prev[11] = 11'b11111110100;
        h_t_prev[12] = 11'b11111111000;
        h_t_prev[13] = 11'b11111110011;
        h_t_prev[14] = 11'b11111111001;
        h_t_prev[15] = 11'b11111111010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 68 timeout!");
                $fdisplay(fd_cycles, "Test Vector  68: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  68: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 68");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 69
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111011111;
        x_t[1] = 11'b11111101111;
        x_t[2] = 11'b11111101110;
        x_t[3] = 11'b11111110101;
        x_t[4] = 11'b11111110111;
        x_t[5] = 11'b11111110111;
        x_t[6] = 11'b11111101110;
        x_t[7] = 11'b11111101100;
        x_t[8] = 11'b11111110111;
        x_t[9] = 11'b11111110111;
        x_t[10] = 11'b11111111001;
        x_t[11] = 11'b11111111100;
        x_t[12] = 11'b11111110110;
        x_t[13] = 11'b11111101111;
        x_t[14] = 11'b11111101010;
        x_t[15] = 11'b11111110011;
        x_t[16] = 11'b11111111001;
        x_t[17] = 11'b11111111100;
        x_t[18] = 11'b11111110101;
        x_t[19] = 11'b11111110110;
        x_t[20] = 11'b11111111100;
        x_t[21] = 11'b11111001011;
        x_t[22] = 11'b11111001001;
        x_t[23] = 11'b11111010001;
        x_t[24] = 11'b11111001001;
        x_t[25] = 11'b11111001011;
        x_t[26] = 11'b11111011001;
        x_t[27] = 11'b11111011011;
        x_t[28] = 11'b11111010111;
        x_t[29] = 11'b11111001110;
        x_t[30] = 11'b11111100110;
        x_t[31] = 11'b11111100100;
        x_t[32] = 11'b11111100011;
        x_t[33] = 11'b11111101000;
        x_t[34] = 11'b11111101111;
        x_t[35] = 11'b11111101110;
        x_t[36] = 11'b11111101000;
        x_t[37] = 11'b11111110000;
        x_t[38] = 11'b11111011010;
        x_t[39] = 11'b11111101110;
        x_t[40] = 11'b11111100101;
        x_t[41] = 11'b00000010001;
        x_t[42] = 11'b11111000011;
        x_t[43] = 11'b11111101000;
        x_t[44] = 11'b11111100010;
        x_t[45] = 11'b11111110011;
        x_t[46] = 11'b11111101101;
        x_t[47] = 11'b11111110001;
        x_t[48] = 11'b00000000000;
        x_t[49] = 11'b00000000001;
        x_t[50] = 11'b00000000110;
        x_t[51] = 11'b00000001101;
        x_t[52] = 11'b00000001010;
        x_t[53] = 11'b00000001110;
        x_t[54] = 11'b00000001110;
        x_t[55] = 11'b11111110100;
        x_t[56] = 11'b11111111010;
        x_t[57] = 11'b00000010001;
        x_t[58] = 11'b00000010111;
        x_t[59] = 11'b00000010101;
        x_t[60] = 11'b00000000000;
        x_t[61] = 11'b00000001100;
        x_t[62] = 11'b11111111001;
        x_t[63] = 11'b11111111110;
        
        h_t_prev[0] = 11'b11111011111;
        h_t_prev[1] = 11'b11111101111;
        h_t_prev[2] = 11'b11111101110;
        h_t_prev[3] = 11'b11111110101;
        h_t_prev[4] = 11'b11111110111;
        h_t_prev[5] = 11'b11111110111;
        h_t_prev[6] = 11'b11111101110;
        h_t_prev[7] = 11'b11111101100;
        h_t_prev[8] = 11'b11111110111;
        h_t_prev[9] = 11'b11111110111;
        h_t_prev[10] = 11'b11111111001;
        h_t_prev[11] = 11'b11111111100;
        h_t_prev[12] = 11'b11111110110;
        h_t_prev[13] = 11'b11111101111;
        h_t_prev[14] = 11'b11111101010;
        h_t_prev[15] = 11'b11111110011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 69 timeout!");
                $fdisplay(fd_cycles, "Test Vector  69: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  69: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 69");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 70
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111100000;
        x_t[1] = 11'b11111110000;
        x_t[2] = 11'b11111110100;
        x_t[3] = 11'b11111111110;
        x_t[4] = 11'b00000000010;
        x_t[5] = 11'b00000000100;
        x_t[6] = 11'b11111111101;
        x_t[7] = 11'b11111110010;
        x_t[8] = 11'b11111111100;
        x_t[9] = 11'b11111111110;
        x_t[10] = 11'b00000000000;
        x_t[11] = 11'b00000000100;
        x_t[12] = 11'b00000001000;
        x_t[13] = 11'b00000000101;
        x_t[14] = 11'b11111101000;
        x_t[15] = 11'b11111110110;
        x_t[16] = 11'b11111111101;
        x_t[17] = 11'b00000000100;
        x_t[18] = 11'b00000000101;
        x_t[19] = 11'b00000000110;
        x_t[20] = 11'b00000000110;
        x_t[21] = 11'b11111001110;
        x_t[22] = 11'b11111001111;
        x_t[23] = 11'b11111010110;
        x_t[24] = 11'b11111001011;
        x_t[25] = 11'b11111001100;
        x_t[26] = 11'b11111011100;
        x_t[27] = 11'b11111011111;
        x_t[28] = 11'b11111011010;
        x_t[29] = 11'b11111010101;
        x_t[30] = 11'b11111011111;
        x_t[31] = 11'b11111100011;
        x_t[32] = 11'b11111100100;
        x_t[33] = 11'b11111101000;
        x_t[34] = 11'b11111110010;
        x_t[35] = 11'b11111101110;
        x_t[36] = 11'b11111101011;
        x_t[37] = 11'b11111110011;
        x_t[38] = 11'b11111011000;
        x_t[39] = 11'b11111101101;
        x_t[40] = 11'b11111010000;
        x_t[41] = 11'b11111100110;
        x_t[42] = 11'b11110111101;
        x_t[43] = 11'b00000000100;
        x_t[44] = 11'b11111011011;
        x_t[45] = 11'b11111100111;
        x_t[46] = 11'b11111100110;
        x_t[47] = 11'b11111101000;
        x_t[48] = 11'b11111110111;
        x_t[49] = 11'b11111111000;
        x_t[50] = 11'b00000000000;
        x_t[51] = 11'b00000001100;
        x_t[52] = 11'b00000001000;
        x_t[53] = 11'b00000001001;
        x_t[54] = 11'b00000000110;
        x_t[55] = 11'b11111101110;
        x_t[56] = 11'b11111110011;
        x_t[57] = 11'b00000001011;
        x_t[58] = 11'b00000010000;
        x_t[59] = 11'b00000001101;
        x_t[60] = 11'b11111110111;
        x_t[61] = 11'b00000000101;
        x_t[62] = 11'b11111110101;
        x_t[63] = 11'b11111110010;
        
        h_t_prev[0] = 11'b11111100000;
        h_t_prev[1] = 11'b11111110000;
        h_t_prev[2] = 11'b11111110100;
        h_t_prev[3] = 11'b11111111110;
        h_t_prev[4] = 11'b00000000010;
        h_t_prev[5] = 11'b00000000100;
        h_t_prev[6] = 11'b11111111101;
        h_t_prev[7] = 11'b11111110010;
        h_t_prev[8] = 11'b11111111100;
        h_t_prev[9] = 11'b11111111110;
        h_t_prev[10] = 11'b00000000000;
        h_t_prev[11] = 11'b00000000100;
        h_t_prev[12] = 11'b00000001000;
        h_t_prev[13] = 11'b00000000101;
        h_t_prev[14] = 11'b11111101000;
        h_t_prev[15] = 11'b11111110110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 70 timeout!");
                $fdisplay(fd_cycles, "Test Vector  70: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  70: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 70");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 71
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111010001;
        x_t[1] = 11'b11111100100;
        x_t[2] = 11'b11111100111;
        x_t[3] = 11'b11111110111;
        x_t[4] = 11'b11111111011;
        x_t[5] = 11'b11111111100;
        x_t[6] = 11'b11111110010;
        x_t[7] = 11'b11111011111;
        x_t[8] = 11'b11111101110;
        x_t[9] = 11'b11111101111;
        x_t[10] = 11'b11111110100;
        x_t[11] = 11'b11111111111;
        x_t[12] = 11'b00000000101;
        x_t[13] = 11'b11111111001;
        x_t[14] = 11'b11111011111;
        x_t[15] = 11'b11111101000;
        x_t[16] = 11'b11111110001;
        x_t[17] = 11'b11111111100;
        x_t[18] = 11'b00000000010;
        x_t[19] = 11'b00000000110;
        x_t[20] = 11'b00000000010;
        x_t[21] = 11'b11111001010;
        x_t[22] = 11'b11111001100;
        x_t[23] = 11'b11111010110;
        x_t[24] = 11'b11111001000;
        x_t[25] = 11'b11111001001;
        x_t[26] = 11'b11111010111;
        x_t[27] = 11'b11111011111;
        x_t[28] = 11'b11111011011;
        x_t[29] = 11'b11111001110;
        x_t[30] = 11'b11111011110;
        x_t[31] = 11'b11111100000;
        x_t[32] = 11'b11111011110;
        x_t[33] = 11'b11111100011;
        x_t[34] = 11'b11111101111;
        x_t[35] = 11'b11111101110;
        x_t[36] = 11'b11111101110;
        x_t[37] = 11'b11111110010;
        x_t[38] = 11'b11111001100;
        x_t[39] = 11'b11111110011;
        x_t[40] = 11'b11111000101;
        x_t[41] = 11'b11111100111;
        x_t[42] = 11'b11111000010;
        x_t[43] = 11'b11111111011;
        x_t[44] = 11'b11111011100;
        x_t[45] = 11'b11111110001;
        x_t[46] = 11'b11111101101;
        x_t[47] = 11'b11111101101;
        x_t[48] = 11'b11111111000;
        x_t[49] = 11'b11111111010;
        x_t[50] = 11'b00000000110;
        x_t[51] = 11'b00000010101;
        x_t[52] = 11'b00000010001;
        x_t[53] = 11'b00000010011;
        x_t[54] = 11'b00000001111;
        x_t[55] = 11'b11111111001;
        x_t[56] = 11'b11111111100;
        x_t[57] = 11'b00000010110;
        x_t[58] = 11'b00000011000;
        x_t[59] = 11'b00000010100;
        x_t[60] = 11'b11111111000;
        x_t[61] = 11'b00000000101;
        x_t[62] = 11'b11111110111;
        x_t[63] = 11'b11111110001;
        
        h_t_prev[0] = 11'b11111010001;
        h_t_prev[1] = 11'b11111100100;
        h_t_prev[2] = 11'b11111100111;
        h_t_prev[3] = 11'b11111110111;
        h_t_prev[4] = 11'b11111111011;
        h_t_prev[5] = 11'b11111111100;
        h_t_prev[6] = 11'b11111110010;
        h_t_prev[7] = 11'b11111011111;
        h_t_prev[8] = 11'b11111101110;
        h_t_prev[9] = 11'b11111101111;
        h_t_prev[10] = 11'b11111110100;
        h_t_prev[11] = 11'b11111111111;
        h_t_prev[12] = 11'b00000000101;
        h_t_prev[13] = 11'b11111111001;
        h_t_prev[14] = 11'b11111011111;
        h_t_prev[15] = 11'b11111101000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 71 timeout!");
                $fdisplay(fd_cycles, "Test Vector  71: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  71: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 71");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 72
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111010101;
        x_t[1] = 11'b11111101010;
        x_t[2] = 11'b11111101010;
        x_t[3] = 11'b11111111011;
        x_t[4] = 11'b00000000100;
        x_t[5] = 11'b00000001001;
        x_t[6] = 11'b11111111010;
        x_t[7] = 11'b11111101011;
        x_t[8] = 11'b11111110010;
        x_t[9] = 11'b11111110100;
        x_t[10] = 11'b11111111100;
        x_t[11] = 11'b00000001011;
        x_t[12] = 11'b00000010011;
        x_t[13] = 11'b00000001001;
        x_t[14] = 11'b11111101000;
        x_t[15] = 11'b11111101011;
        x_t[16] = 11'b11111110101;
        x_t[17] = 11'b00000000100;
        x_t[18] = 11'b00000010001;
        x_t[19] = 11'b00000010101;
        x_t[20] = 11'b00000010011;
        x_t[21] = 11'b11111010001;
        x_t[22] = 11'b11111010100;
        x_t[23] = 11'b11111011010;
        x_t[24] = 11'b11111001110;
        x_t[25] = 11'b11111001111;
        x_t[26] = 11'b11111100000;
        x_t[27] = 11'b11111100111;
        x_t[28] = 11'b11111011111;
        x_t[29] = 11'b11111010100;
        x_t[30] = 11'b11111101010;
        x_t[31] = 11'b11111101011;
        x_t[32] = 11'b11111100100;
        x_t[33] = 11'b11111101010;
        x_t[34] = 11'b11111110111;
        x_t[35] = 11'b11111110111;
        x_t[36] = 11'b11111110111;
        x_t[37] = 11'b11111110010;
        x_t[38] = 11'b11111011101;
        x_t[39] = 11'b11111111011;
        x_t[40] = 11'b11111101000;
        x_t[41] = 11'b11111110101;
        x_t[42] = 11'b11111000111;
        x_t[43] = 11'b00000000101;
        x_t[44] = 11'b11111100101;
        x_t[45] = 11'b00000000001;
        x_t[46] = 11'b11111110110;
        x_t[47] = 11'b11111110011;
        x_t[48] = 11'b11111111010;
        x_t[49] = 11'b00000000010;
        x_t[50] = 11'b00000001110;
        x_t[51] = 11'b00000011110;
        x_t[52] = 11'b00000011000;
        x_t[53] = 11'b00000011010;
        x_t[54] = 11'b00000010110;
        x_t[55] = 11'b00000000001;
        x_t[56] = 11'b00000000011;
        x_t[57] = 11'b00000011011;
        x_t[58] = 11'b00000011110;
        x_t[59] = 11'b00000011001;
        x_t[60] = 11'b00000000010;
        x_t[61] = 11'b00000010001;
        x_t[62] = 11'b00000000010;
        x_t[63] = 11'b11111111110;
        
        h_t_prev[0] = 11'b11111010101;
        h_t_prev[1] = 11'b11111101010;
        h_t_prev[2] = 11'b11111101010;
        h_t_prev[3] = 11'b11111111011;
        h_t_prev[4] = 11'b00000000100;
        h_t_prev[5] = 11'b00000001001;
        h_t_prev[6] = 11'b11111111010;
        h_t_prev[7] = 11'b11111101011;
        h_t_prev[8] = 11'b11111110010;
        h_t_prev[9] = 11'b11111110100;
        h_t_prev[10] = 11'b11111111100;
        h_t_prev[11] = 11'b00000001011;
        h_t_prev[12] = 11'b00000010011;
        h_t_prev[13] = 11'b00000001001;
        h_t_prev[14] = 11'b11111101000;
        h_t_prev[15] = 11'b11111101011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 72 timeout!");
                $fdisplay(fd_cycles, "Test Vector  72: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  72: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 72");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 73
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111100100;
        x_t[1] = 11'b11111110010;
        x_t[2] = 11'b11111110000;
        x_t[3] = 11'b00000000000;
        x_t[4] = 11'b00000000110;
        x_t[5] = 11'b00000000111;
        x_t[6] = 11'b11111111100;
        x_t[7] = 11'b11111101110;
        x_t[8] = 11'b11111110010;
        x_t[9] = 11'b11111110111;
        x_t[10] = 11'b11111111111;
        x_t[11] = 11'b00000001001;
        x_t[12] = 11'b00000001110;
        x_t[13] = 11'b00000000001;
        x_t[14] = 11'b11111100001;
        x_t[15] = 11'b11111101010;
        x_t[16] = 11'b11111111000;
        x_t[17] = 11'b00000000101;
        x_t[18] = 11'b00000001101;
        x_t[19] = 11'b00000001110;
        x_t[20] = 11'b00000001010;
        x_t[21] = 11'b11111011000;
        x_t[22] = 11'b11111011001;
        x_t[23] = 11'b11111011101;
        x_t[24] = 11'b11111010101;
        x_t[25] = 11'b11111010110;
        x_t[26] = 11'b11111100110;
        x_t[27] = 11'b11111100111;
        x_t[28] = 11'b11111011101;
        x_t[29] = 11'b11111011011;
        x_t[30] = 11'b11111110011;
        x_t[31] = 11'b11111101011;
        x_t[32] = 11'b11111101011;
        x_t[33] = 11'b11111101110;
        x_t[34] = 11'b11111110111;
        x_t[35] = 11'b11111111000;
        x_t[36] = 11'b11111110001;
        x_t[37] = 11'b11111110010;
        x_t[38] = 11'b11111100101;
        x_t[39] = 11'b11111110011;
        x_t[40] = 11'b11111011110;
        x_t[41] = 11'b00000001011;
        x_t[42] = 11'b11111000110;
        x_t[43] = 11'b11111101110;
        x_t[44] = 11'b11111100111;
        x_t[45] = 11'b11111101001;
        x_t[46] = 11'b11111111000;
        x_t[47] = 11'b11111110001;
        x_t[48] = 11'b11111111010;
        x_t[49] = 11'b11111111101;
        x_t[50] = 11'b00000000111;
        x_t[51] = 11'b00000001100;
        x_t[52] = 11'b00000000101;
        x_t[53] = 11'b00000000101;
        x_t[54] = 11'b11111111100;
        x_t[55] = 11'b11111111101;
        x_t[56] = 11'b11111111110;
        x_t[57] = 11'b00000001110;
        x_t[58] = 11'b00000001001;
        x_t[59] = 11'b00000000010;
        x_t[60] = 11'b00000000111;
        x_t[61] = 11'b00000010000;
        x_t[62] = 11'b11111111111;
        x_t[63] = 11'b11111111011;
        
        h_t_prev[0] = 11'b11111100100;
        h_t_prev[1] = 11'b11111110010;
        h_t_prev[2] = 11'b11111110000;
        h_t_prev[3] = 11'b00000000000;
        h_t_prev[4] = 11'b00000000110;
        h_t_prev[5] = 11'b00000000111;
        h_t_prev[6] = 11'b11111111100;
        h_t_prev[7] = 11'b11111101110;
        h_t_prev[8] = 11'b11111110010;
        h_t_prev[9] = 11'b11111110111;
        h_t_prev[10] = 11'b11111111111;
        h_t_prev[11] = 11'b00000001001;
        h_t_prev[12] = 11'b00000001110;
        h_t_prev[13] = 11'b00000000001;
        h_t_prev[14] = 11'b11111100001;
        h_t_prev[15] = 11'b11111101010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 73 timeout!");
                $fdisplay(fd_cycles, "Test Vector  73: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  73: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 73");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 74
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111100111;
        x_t[1] = 11'b11111111000;
        x_t[2] = 11'b11111110011;
        x_t[3] = 11'b00000000010;
        x_t[4] = 11'b00000000010;
        x_t[5] = 11'b00000000001;
        x_t[6] = 11'b11111111000;
        x_t[7] = 11'b11111110011;
        x_t[8] = 11'b11111110111;
        x_t[9] = 11'b11111111100;
        x_t[10] = 11'b00000000010;
        x_t[11] = 11'b00000001001;
        x_t[12] = 11'b00000001001;
        x_t[13] = 11'b11111111111;
        x_t[14] = 11'b11111101100;
        x_t[15] = 11'b11111110100;
        x_t[16] = 11'b11111111110;
        x_t[17] = 11'b00000001001;
        x_t[18] = 11'b00000000110;
        x_t[19] = 11'b00000000110;
        x_t[20] = 11'b00000000101;
        x_t[21] = 11'b11111011010;
        x_t[22] = 11'b11111011010;
        x_t[23] = 11'b11111100000;
        x_t[24] = 11'b11111011000;
        x_t[25] = 11'b11111011000;
        x_t[26] = 11'b11111101010;
        x_t[27] = 11'b11111101010;
        x_t[28] = 11'b11111100010;
        x_t[29] = 11'b11111011010;
        x_t[30] = 11'b11111110100;
        x_t[31] = 11'b11111101111;
        x_t[32] = 11'b11111101111;
        x_t[33] = 11'b11111110010;
        x_t[34] = 11'b11111111010;
        x_t[35] = 11'b11111111010;
        x_t[36] = 11'b11111110100;
        x_t[37] = 11'b11111111100;
        x_t[38] = 11'b11111011011;
        x_t[39] = 11'b11111111011;
        x_t[40] = 11'b11111011001;
        x_t[41] = 11'b00000011000;
        x_t[42] = 11'b11111001111;
        x_t[43] = 11'b11111100111;
        x_t[44] = 11'b11111101100;
        x_t[45] = 11'b11111110010;
        x_t[46] = 11'b11111111110;
        x_t[47] = 11'b11111111111;
        x_t[48] = 11'b00000001001;
        x_t[49] = 11'b00000001000;
        x_t[50] = 11'b00000001100;
        x_t[51] = 11'b00000001101;
        x_t[52] = 11'b00000000111;
        x_t[53] = 11'b00000000111;
        x_t[54] = 11'b00000000101;
        x_t[55] = 11'b00000001101;
        x_t[56] = 11'b00000001011;
        x_t[57] = 11'b00000010101;
        x_t[58] = 11'b00000001001;
        x_t[59] = 11'b00000000101;
        x_t[60] = 11'b00000001100;
        x_t[61] = 11'b00000001100;
        x_t[62] = 11'b11111111001;
        x_t[63] = 11'b11111111010;
        
        h_t_prev[0] = 11'b11111100111;
        h_t_prev[1] = 11'b11111111000;
        h_t_prev[2] = 11'b11111110011;
        h_t_prev[3] = 11'b00000000010;
        h_t_prev[4] = 11'b00000000010;
        h_t_prev[5] = 11'b00000000001;
        h_t_prev[6] = 11'b11111111000;
        h_t_prev[7] = 11'b11111110011;
        h_t_prev[8] = 11'b11111110111;
        h_t_prev[9] = 11'b11111111100;
        h_t_prev[10] = 11'b00000000010;
        h_t_prev[11] = 11'b00000001001;
        h_t_prev[12] = 11'b00000001001;
        h_t_prev[13] = 11'b11111111111;
        h_t_prev[14] = 11'b11111101100;
        h_t_prev[15] = 11'b11111110100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 74 timeout!");
                $fdisplay(fd_cycles, "Test Vector  74: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  74: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 74");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 75
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111100100;
        x_t[1] = 11'b11111111010;
        x_t[2] = 11'b11111110100;
        x_t[3] = 11'b00000000010;
        x_t[4] = 11'b00000000001;
        x_t[5] = 11'b00000000100;
        x_t[6] = 11'b11111111010;
        x_t[7] = 11'b11111111100;
        x_t[8] = 11'b00000000000;
        x_t[9] = 11'b11111111110;
        x_t[10] = 11'b11111111111;
        x_t[11] = 11'b00000001001;
        x_t[12] = 11'b00000000110;
        x_t[13] = 11'b00000000001;
        x_t[14] = 11'b11111110111;
        x_t[15] = 11'b11111111101;
        x_t[16] = 11'b00000000000;
        x_t[17] = 11'b00000000100;
        x_t[18] = 11'b00000000000;
        x_t[19] = 11'b11111111111;
        x_t[20] = 11'b00000000010;
        x_t[21] = 11'b11111011011;
        x_t[22] = 11'b11111011101;
        x_t[23] = 11'b11111100010;
        x_t[24] = 11'b11111010101;
        x_t[25] = 11'b11111010110;
        x_t[26] = 11'b11111101010;
        x_t[27] = 11'b11111101011;
        x_t[28] = 11'b11111100101;
        x_t[29] = 11'b11111010110;
        x_t[30] = 11'b11111101100;
        x_t[31] = 11'b11111101010;
        x_t[32] = 11'b11111101001;
        x_t[33] = 11'b11111101100;
        x_t[34] = 11'b11111110101;
        x_t[35] = 11'b11111110011;
        x_t[36] = 11'b11111110001;
        x_t[37] = 11'b11111110101;
        x_t[38] = 11'b11111011111;
        x_t[39] = 11'b11111101111;
        x_t[40] = 11'b11111100111;
        x_t[41] = 11'b11111101100;
        x_t[42] = 11'b11111010111;
        x_t[43] = 11'b11111011011;
        x_t[44] = 11'b11111101110;
        x_t[45] = 11'b11111100100;
        x_t[46] = 11'b11111111110;
        x_t[47] = 11'b11111111100;
        x_t[48] = 11'b00000000011;
        x_t[49] = 11'b11111111101;
        x_t[50] = 11'b11111111010;
        x_t[51] = 11'b11111111010;
        x_t[52] = 11'b11111110001;
        x_t[53] = 11'b11111110111;
        x_t[54] = 11'b11111110110;
        x_t[55] = 11'b00000000111;
        x_t[56] = 11'b00000000011;
        x_t[57] = 11'b00000000101;
        x_t[58] = 11'b11111110111;
        x_t[59] = 11'b11111111100;
        x_t[60] = 11'b00000001101;
        x_t[61] = 11'b00000000111;
        x_t[62] = 11'b11111110101;
        x_t[63] = 11'b11111111101;
        
        h_t_prev[0] = 11'b11111100100;
        h_t_prev[1] = 11'b11111111010;
        h_t_prev[2] = 11'b11111110100;
        h_t_prev[3] = 11'b00000000010;
        h_t_prev[4] = 11'b00000000001;
        h_t_prev[5] = 11'b00000000100;
        h_t_prev[6] = 11'b11111111010;
        h_t_prev[7] = 11'b11111111100;
        h_t_prev[8] = 11'b00000000000;
        h_t_prev[9] = 11'b11111111110;
        h_t_prev[10] = 11'b11111111111;
        h_t_prev[11] = 11'b00000001001;
        h_t_prev[12] = 11'b00000000110;
        h_t_prev[13] = 11'b00000000001;
        h_t_prev[14] = 11'b11111110111;
        h_t_prev[15] = 11'b11111111101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 75 timeout!");
                $fdisplay(fd_cycles, "Test Vector  75: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  75: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 75");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 76
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111011101;
        x_t[1] = 11'b11111101000;
        x_t[2] = 11'b11111100111;
        x_t[3] = 11'b11111110111;
        x_t[4] = 11'b11111110110;
        x_t[5] = 11'b11111110011;
        x_t[6] = 11'b11111101011;
        x_t[7] = 11'b11111101100;
        x_t[8] = 11'b11111110001;
        x_t[9] = 11'b11111101110;
        x_t[10] = 11'b11111101111;
        x_t[11] = 11'b11111111010;
        x_t[12] = 11'b11111110011;
        x_t[13] = 11'b11111101001;
        x_t[14] = 11'b11111101110;
        x_t[15] = 11'b11111110000;
        x_t[16] = 11'b11111110001;
        x_t[17] = 11'b11111110001;
        x_t[18] = 11'b11111101101;
        x_t[19] = 11'b11111101110;
        x_t[20] = 11'b11111110000;
        x_t[21] = 11'b11111011011;
        x_t[22] = 11'b11111011100;
        x_t[23] = 11'b11111100001;
        x_t[24] = 11'b11111010110;
        x_t[25] = 11'b11111010110;
        x_t[26] = 11'b11111101010;
        x_t[27] = 11'b11111101000;
        x_t[28] = 11'b11111100010;
        x_t[29] = 11'b11111011001;
        x_t[30] = 11'b11111101100;
        x_t[31] = 11'b11111100110;
        x_t[32] = 11'b11111101010;
        x_t[33] = 11'b11111101111;
        x_t[34] = 11'b11111110110;
        x_t[35] = 11'b11111110011;
        x_t[36] = 11'b11111101100;
        x_t[37] = 11'b11111110001;
        x_t[38] = 11'b11111101101;
        x_t[39] = 11'b11111101010;
        x_t[40] = 11'b11111110100;
        x_t[41] = 11'b11111100010;
        x_t[42] = 11'b11111101010;
        x_t[43] = 11'b11111100111;
        x_t[44] = 11'b11111110000;
        x_t[45] = 11'b11111101100;
        x_t[46] = 11'b00000000001;
        x_t[47] = 11'b11111111110;
        x_t[48] = 11'b00000000010;
        x_t[49] = 11'b11111111010;
        x_t[50] = 11'b11111110110;
        x_t[51] = 11'b11111110110;
        x_t[52] = 11'b11111110010;
        x_t[53] = 11'b11111111101;
        x_t[54] = 11'b00000000000;
        x_t[55] = 11'b00000001100;
        x_t[56] = 11'b00000001000;
        x_t[57] = 11'b00000000100;
        x_t[58] = 11'b11111111010;
        x_t[59] = 11'b00000000110;
        x_t[60] = 11'b00000001100;
        x_t[61] = 11'b00000000110;
        x_t[62] = 11'b11111110111;
        x_t[63] = 11'b00000000111;
        
        h_t_prev[0] = 11'b11111011101;
        h_t_prev[1] = 11'b11111101000;
        h_t_prev[2] = 11'b11111100111;
        h_t_prev[3] = 11'b11111110111;
        h_t_prev[4] = 11'b11111110110;
        h_t_prev[5] = 11'b11111110011;
        h_t_prev[6] = 11'b11111101011;
        h_t_prev[7] = 11'b11111101100;
        h_t_prev[8] = 11'b11111110001;
        h_t_prev[9] = 11'b11111101110;
        h_t_prev[10] = 11'b11111101111;
        h_t_prev[11] = 11'b11111111010;
        h_t_prev[12] = 11'b11111110011;
        h_t_prev[13] = 11'b11111101001;
        h_t_prev[14] = 11'b11111101110;
        h_t_prev[15] = 11'b11111110000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 76 timeout!");
                $fdisplay(fd_cycles, "Test Vector  76: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  76: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 76");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 77
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111110001;
        x_t[1] = 11'b11111111011;
        x_t[2] = 11'b11111111000;
        x_t[3] = 11'b00000000111;
        x_t[4] = 11'b00000000110;
        x_t[5] = 11'b00000000001;
        x_t[6] = 11'b11111110101;
        x_t[7] = 11'b00000001011;
        x_t[8] = 11'b00000000110;
        x_t[9] = 11'b00000000000;
        x_t[10] = 11'b00000000001;
        x_t[11] = 11'b00000001101;
        x_t[12] = 11'b00000000100;
        x_t[13] = 11'b11111111001;
        x_t[14] = 11'b00000000011;
        x_t[15] = 11'b00000000101;
        x_t[16] = 11'b00000000010;
        x_t[17] = 11'b00000000010;
        x_t[18] = 11'b11111111100;
        x_t[19] = 11'b11111111111;
        x_t[20] = 11'b00000000100;
        x_t[21] = 11'b11111100011;
        x_t[22] = 11'b11111100101;
        x_t[23] = 11'b11111100111;
        x_t[24] = 11'b11111100010;
        x_t[25] = 11'b11111100010;
        x_t[26] = 11'b11111110101;
        x_t[27] = 11'b11111110010;
        x_t[28] = 11'b11111100111;
        x_t[29] = 11'b11111101001;
        x_t[30] = 11'b00000000000;
        x_t[31] = 11'b11111110110;
        x_t[32] = 11'b11111110111;
        x_t[33] = 11'b11111111010;
        x_t[34] = 11'b00000000011;
        x_t[35] = 11'b11111111111;
        x_t[36] = 11'b11111110111;
        x_t[37] = 11'b11111111001;
        x_t[38] = 11'b11111111100;
        x_t[39] = 11'b11111101101;
        x_t[40] = 11'b00000000010;
        x_t[41] = 11'b11111110000;
        x_t[42] = 11'b11111101000;
        x_t[43] = 11'b11111111101;
        x_t[44] = 11'b00000000000;
        x_t[45] = 11'b11111110010;
        x_t[46] = 11'b00000001011;
        x_t[47] = 11'b00000001000;
        x_t[48] = 11'b00000001100;
        x_t[49] = 11'b00000000001;
        x_t[50] = 11'b11111111010;
        x_t[51] = 11'b11111111000;
        x_t[52] = 11'b11111110010;
        x_t[53] = 11'b11111111011;
        x_t[54] = 11'b11111111101;
        x_t[55] = 11'b00000001110;
        x_t[56] = 11'b00000001010;
        x_t[57] = 11'b00000000010;
        x_t[58] = 11'b11111110110;
        x_t[59] = 11'b11111111010;
        x_t[60] = 11'b00000001110;
        x_t[61] = 11'b00000001010;
        x_t[62] = 11'b11111110111;
        x_t[63] = 11'b00000010010;
        
        h_t_prev[0] = 11'b11111110001;
        h_t_prev[1] = 11'b11111111011;
        h_t_prev[2] = 11'b11111111000;
        h_t_prev[3] = 11'b00000000111;
        h_t_prev[4] = 11'b00000000110;
        h_t_prev[5] = 11'b00000000001;
        h_t_prev[6] = 11'b11111110101;
        h_t_prev[7] = 11'b00000001011;
        h_t_prev[8] = 11'b00000000110;
        h_t_prev[9] = 11'b00000000000;
        h_t_prev[10] = 11'b00000000001;
        h_t_prev[11] = 11'b00000001101;
        h_t_prev[12] = 11'b00000000100;
        h_t_prev[13] = 11'b11111111001;
        h_t_prev[14] = 11'b00000000011;
        h_t_prev[15] = 11'b00000000101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 77 timeout!");
                $fdisplay(fd_cycles, "Test Vector  77: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  77: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 77");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 78
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111110101;
        x_t[1] = 11'b11111111011;
        x_t[2] = 11'b11111110100;
        x_t[3] = 11'b11111111111;
        x_t[4] = 11'b11111111101;
        x_t[5] = 11'b11111111001;
        x_t[6] = 11'b11111101110;
        x_t[7] = 11'b00000000100;
        x_t[8] = 11'b11111111111;
        x_t[9] = 11'b11111111001;
        x_t[10] = 11'b11111110111;
        x_t[11] = 11'b11111111101;
        x_t[12] = 11'b11111110001;
        x_t[13] = 11'b11111101001;
        x_t[14] = 11'b11111110100;
        x_t[15] = 11'b11111111000;
        x_t[16] = 11'b11111110101;
        x_t[17] = 11'b11111110101;
        x_t[18] = 11'b11111101011;
        x_t[19] = 11'b11111101001;
        x_t[20] = 11'b11111101010;
        x_t[21] = 11'b11111011110;
        x_t[22] = 11'b11111011111;
        x_t[23] = 11'b11111100000;
        x_t[24] = 11'b11111011011;
        x_t[25] = 11'b11111011100;
        x_t[26] = 11'b11111101010;
        x_t[27] = 11'b11111101001;
        x_t[28] = 11'b11111100000;
        x_t[29] = 11'b11111011001;
        x_t[30] = 11'b11111111101;
        x_t[31] = 11'b11111101000;
        x_t[32] = 11'b11111101000;
        x_t[33] = 11'b11111101001;
        x_t[34] = 11'b11111110011;
        x_t[35] = 11'b11111110000;
        x_t[36] = 11'b11111101001;
        x_t[37] = 11'b11111101011;
        x_t[38] = 11'b11111100100;
        x_t[39] = 11'b11111011110;
        x_t[40] = 11'b11111100100;
        x_t[41] = 11'b11111101100;
        x_t[42] = 11'b11111001011;
        x_t[43] = 11'b11111011101;
        x_t[44] = 11'b11111101001;
        x_t[45] = 11'b11111001100;
        x_t[46] = 11'b11111110010;
        x_t[47] = 11'b11111101110;
        x_t[48] = 11'b11111110000;
        x_t[49] = 11'b11111100111;
        x_t[50] = 11'b11111100011;
        x_t[51] = 11'b11111100000;
        x_t[52] = 11'b11111011001;
        x_t[53] = 11'b11111011111;
        x_t[54] = 11'b11111011100;
        x_t[55] = 11'b11111111001;
        x_t[56] = 11'b11111110110;
        x_t[57] = 11'b11111101110;
        x_t[58] = 11'b11111100011;
        x_t[59] = 11'b11111100101;
        x_t[60] = 11'b00000000111;
        x_t[61] = 11'b11111111111;
        x_t[62] = 11'b11111100110;
        x_t[63] = 11'b00000000110;
        
        h_t_prev[0] = 11'b11111110101;
        h_t_prev[1] = 11'b11111111011;
        h_t_prev[2] = 11'b11111110100;
        h_t_prev[3] = 11'b11111111111;
        h_t_prev[4] = 11'b11111111101;
        h_t_prev[5] = 11'b11111111001;
        h_t_prev[6] = 11'b11111101110;
        h_t_prev[7] = 11'b00000000100;
        h_t_prev[8] = 11'b11111111111;
        h_t_prev[9] = 11'b11111111001;
        h_t_prev[10] = 11'b11111110111;
        h_t_prev[11] = 11'b11111111101;
        h_t_prev[12] = 11'b11111110001;
        h_t_prev[13] = 11'b11111101001;
        h_t_prev[14] = 11'b11111110100;
        h_t_prev[15] = 11'b11111111000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 78 timeout!");
                $fdisplay(fd_cycles, "Test Vector  78: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  78: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 78");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 79
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111101001;
        x_t[1] = 11'b11111110010;
        x_t[2] = 11'b11111101101;
        x_t[3] = 11'b11111110100;
        x_t[4] = 11'b11111110101;
        x_t[5] = 11'b11111110011;
        x_t[6] = 11'b11111101110;
        x_t[7] = 11'b11111110000;
        x_t[8] = 11'b11111110001;
        x_t[9] = 11'b11111101111;
        x_t[10] = 11'b11111101101;
        x_t[11] = 11'b11111110111;
        x_t[12] = 11'b11111101100;
        x_t[13] = 11'b11111101001;
        x_t[14] = 11'b11111100111;
        x_t[15] = 11'b11111101001;
        x_t[16] = 11'b11111101010;
        x_t[17] = 11'b11111101011;
        x_t[18] = 11'b11111100111;
        x_t[19] = 11'b11111100111;
        x_t[20] = 11'b11111101001;
        x_t[21] = 11'b11111011111;
        x_t[22] = 11'b11111100000;
        x_t[23] = 11'b11111100001;
        x_t[24] = 11'b11111011110;
        x_t[25] = 11'b11111011101;
        x_t[26] = 11'b11111101111;
        x_t[27] = 11'b11111101100;
        x_t[28] = 11'b11111100000;
        x_t[29] = 11'b11111100000;
        x_t[30] = 11'b11111111010;
        x_t[31] = 11'b11111101011;
        x_t[32] = 11'b11111110000;
        x_t[33] = 11'b11111110010;
        x_t[34] = 11'b11111111001;
        x_t[35] = 11'b11111110110;
        x_t[36] = 11'b11111101111;
        x_t[37] = 11'b11111110001;
        x_t[38] = 11'b11111101011;
        x_t[39] = 11'b11111110100;
        x_t[40] = 11'b11111110011;
        x_t[41] = 11'b00000001100;
        x_t[42] = 11'b11111010010;
        x_t[43] = 11'b11111010000;
        x_t[44] = 11'b11111101011;
        x_t[45] = 11'b11111011001;
        x_t[46] = 11'b11111110101;
        x_t[47] = 11'b11111101110;
        x_t[48] = 11'b11111110001;
        x_t[49] = 11'b11111101100;
        x_t[50] = 11'b11111101011;
        x_t[51] = 11'b11111110000;
        x_t[52] = 11'b11111101001;
        x_t[53] = 11'b11111101110;
        x_t[54] = 11'b11111101011;
        x_t[55] = 11'b11111111100;
        x_t[56] = 11'b11111111001;
        x_t[57] = 11'b11111111001;
        x_t[58] = 11'b11111110110;
        x_t[59] = 11'b11111110110;
        x_t[60] = 11'b11111111111;
        x_t[61] = 11'b11111110111;
        x_t[62] = 11'b11111011111;
        x_t[63] = 11'b11111111011;
        
        h_t_prev[0] = 11'b11111101001;
        h_t_prev[1] = 11'b11111110010;
        h_t_prev[2] = 11'b11111101101;
        h_t_prev[3] = 11'b11111110100;
        h_t_prev[4] = 11'b11111110101;
        h_t_prev[5] = 11'b11111110011;
        h_t_prev[6] = 11'b11111101110;
        h_t_prev[7] = 11'b11111110000;
        h_t_prev[8] = 11'b11111110001;
        h_t_prev[9] = 11'b11111101111;
        h_t_prev[10] = 11'b11111101101;
        h_t_prev[11] = 11'b11111110111;
        h_t_prev[12] = 11'b11111101100;
        h_t_prev[13] = 11'b11111101001;
        h_t_prev[14] = 11'b11111100111;
        h_t_prev[15] = 11'b11111101001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 79 timeout!");
                $fdisplay(fd_cycles, "Test Vector  79: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  79: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 79");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 80
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111101011;
        x_t[1] = 11'b11111110110;
        x_t[2] = 11'b11111110100;
        x_t[3] = 11'b11111111101;
        x_t[4] = 11'b11111111111;
        x_t[5] = 11'b00000000000;
        x_t[6] = 11'b11111110101;
        x_t[7] = 11'b11111111000;
        x_t[8] = 11'b11111110101;
        x_t[9] = 11'b11111110100;
        x_t[10] = 11'b11111110101;
        x_t[11] = 11'b00000000001;
        x_t[12] = 11'b11111111011;
        x_t[13] = 11'b11111111000;
        x_t[14] = 11'b11111101011;
        x_t[15] = 11'b11111101101;
        x_t[16] = 11'b11111110010;
        x_t[17] = 11'b11111110010;
        x_t[18] = 11'b11111110101;
        x_t[19] = 11'b11111111000;
        x_t[20] = 11'b11111111000;
        x_t[21] = 11'b11111100000;
        x_t[22] = 11'b11111011110;
        x_t[23] = 11'b11111100000;
        x_t[24] = 11'b11111011110;
        x_t[25] = 11'b11111011111;
        x_t[26] = 11'b11111101101;
        x_t[27] = 11'b11111101010;
        x_t[28] = 11'b11111011111;
        x_t[29] = 11'b11111100011;
        x_t[30] = 11'b11111110101;
        x_t[31] = 11'b11111101110;
        x_t[32] = 11'b11111101111;
        x_t[33] = 11'b11111110011;
        x_t[34] = 11'b11111111001;
        x_t[35] = 11'b11111110100;
        x_t[36] = 11'b11111101110;
        x_t[37] = 11'b11111110001;
        x_t[38] = 11'b11111101100;
        x_t[39] = 11'b11111110111;
        x_t[40] = 11'b11111011010;
        x_t[41] = 11'b11111111010;
        x_t[42] = 11'b11111001111;
        x_t[43] = 11'b11111110111;
        x_t[44] = 11'b11111101001;
        x_t[45] = 11'b11111101101;
        x_t[46] = 11'b11111110001;
        x_t[47] = 11'b11111101110;
        x_t[48] = 11'b11111110001;
        x_t[49] = 11'b11111110011;
        x_t[50] = 11'b11111110101;
        x_t[51] = 11'b11111111110;
        x_t[52] = 11'b11111111010;
        x_t[53] = 11'b11111111110;
        x_t[54] = 11'b11111111011;
        x_t[55] = 11'b11111111000;
        x_t[56] = 11'b11111110101;
        x_t[57] = 11'b00000000001;
        x_t[58] = 11'b00000000100;
        x_t[59] = 11'b00000000100;
        x_t[60] = 11'b11111111100;
        x_t[61] = 11'b11111111010;
        x_t[62] = 11'b11111101011;
        x_t[63] = 11'b11111111110;
        
        h_t_prev[0] = 11'b11111101011;
        h_t_prev[1] = 11'b11111110110;
        h_t_prev[2] = 11'b11111110100;
        h_t_prev[3] = 11'b11111111101;
        h_t_prev[4] = 11'b11111111111;
        h_t_prev[5] = 11'b00000000000;
        h_t_prev[6] = 11'b11111110101;
        h_t_prev[7] = 11'b11111111000;
        h_t_prev[8] = 11'b11111110101;
        h_t_prev[9] = 11'b11111110100;
        h_t_prev[10] = 11'b11111110101;
        h_t_prev[11] = 11'b00000000001;
        h_t_prev[12] = 11'b11111111011;
        h_t_prev[13] = 11'b11111111000;
        h_t_prev[14] = 11'b11111101011;
        h_t_prev[15] = 11'b11111101101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 80 timeout!");
                $fdisplay(fd_cycles, "Test Vector  80: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  80: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 80");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 81
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000001110;
        x_t[1] = 11'b00000001110;
        x_t[2] = 11'b00000000110;
        x_t[3] = 11'b00000001100;
        x_t[4] = 11'b00000010000;
        x_t[5] = 11'b00000000111;
        x_t[6] = 11'b00000000111;
        x_t[7] = 11'b00000000011;
        x_t[8] = 11'b00000001010;
        x_t[9] = 11'b00000001100;
        x_t[10] = 11'b00000010001;
        x_t[11] = 11'b00000000010;
        x_t[12] = 11'b00000001011;
        x_t[13] = 11'b00000010000;
        x_t[14] = 11'b00000001011;
        x_t[15] = 11'b00000001100;
        x_t[16] = 11'b00000001101;
        x_t[17] = 11'b00000001011;
        x_t[18] = 11'b00000001011;
        x_t[19] = 11'b00000010000;
        x_t[20] = 11'b00000001000;
        x_t[21] = 11'b00000000100;
        x_t[22] = 11'b00000000110;
        x_t[23] = 11'b11111111100;
        x_t[24] = 11'b11111111011;
        x_t[25] = 11'b11111111100;
        x_t[26] = 11'b11111111100;
        x_t[27] = 11'b11111111101;
        x_t[28] = 11'b00000000100;
        x_t[29] = 11'b00000000110;
        x_t[30] = 11'b11111111100;
        x_t[31] = 11'b11111110110;
        x_t[32] = 11'b11111111101;
        x_t[33] = 11'b11111111011;
        x_t[34] = 11'b11111111000;
        x_t[35] = 11'b11111111011;
        x_t[36] = 11'b11111111011;
        x_t[37] = 11'b00000001000;
        x_t[38] = 11'b11111111100;
        x_t[39] = 11'b00000001100;
        x_t[40] = 11'b11111111111;
        x_t[41] = 11'b11111110000;
        x_t[42] = 11'b11111111011;
        x_t[43] = 11'b00000011110;
        x_t[44] = 11'b11111110001;
        x_t[45] = 11'b00000010101;
        x_t[46] = 11'b00000001000;
        x_t[47] = 11'b00000000111;
        x_t[48] = 11'b00000001001;
        x_t[49] = 11'b00000001000;
        x_t[50] = 11'b00000001101;
        x_t[51] = 11'b00000001111;
        x_t[52] = 11'b00000001101;
        x_t[53] = 11'b00000001011;
        x_t[54] = 11'b00000000111;
        x_t[55] = 11'b00000001010;
        x_t[56] = 11'b00000000111;
        x_t[57] = 11'b00000010010;
        x_t[58] = 11'b00000010101;
        x_t[59] = 11'b00000010111;
        x_t[60] = 11'b00000010111;
        x_t[61] = 11'b00000100101;
        x_t[62] = 11'b00000010010;
        x_t[63] = 11'b00000001111;
        
        h_t_prev[0] = 11'b00000001110;
        h_t_prev[1] = 11'b00000001110;
        h_t_prev[2] = 11'b00000000110;
        h_t_prev[3] = 11'b00000001100;
        h_t_prev[4] = 11'b00000010000;
        h_t_prev[5] = 11'b00000000111;
        h_t_prev[6] = 11'b00000000111;
        h_t_prev[7] = 11'b00000000011;
        h_t_prev[8] = 11'b00000001010;
        h_t_prev[9] = 11'b00000001100;
        h_t_prev[10] = 11'b00000010001;
        h_t_prev[11] = 11'b00000000010;
        h_t_prev[12] = 11'b00000001011;
        h_t_prev[13] = 11'b00000010000;
        h_t_prev[14] = 11'b00000001011;
        h_t_prev[15] = 11'b00000001100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 81 timeout!");
                $fdisplay(fd_cycles, "Test Vector  81: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  81: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 81");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 82
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000000101;
        x_t[1] = 11'b00000000110;
        x_t[2] = 11'b00000000001;
        x_t[3] = 11'b00000001010;
        x_t[4] = 11'b00000001101;
        x_t[5] = 11'b00000000000;
        x_t[6] = 11'b11111111110;
        x_t[7] = 11'b11111111011;
        x_t[8] = 11'b00000000011;
        x_t[9] = 11'b00000001001;
        x_t[10] = 11'b00000001101;
        x_t[11] = 11'b00000000011;
        x_t[12] = 11'b00000000110;
        x_t[13] = 11'b00000000111;
        x_t[14] = 11'b00000000110;
        x_t[15] = 11'b00000000100;
        x_t[16] = 11'b00000000110;
        x_t[17] = 11'b00000000110;
        x_t[18] = 11'b00000001000;
        x_t[19] = 11'b00000001011;
        x_t[20] = 11'b00000000010;
        x_t[21] = 11'b00000000111;
        x_t[22] = 11'b00000001001;
        x_t[23] = 11'b00000000000;
        x_t[24] = 11'b11111111100;
        x_t[25] = 11'b11111111101;
        x_t[26] = 11'b00000000000;
        x_t[27] = 11'b00000000001;
        x_t[28] = 11'b00000000110;
        x_t[29] = 11'b00000000011;
        x_t[30] = 11'b11111111100;
        x_t[31] = 11'b11111111000;
        x_t[32] = 11'b00000000001;
        x_t[33] = 11'b00000000001;
        x_t[34] = 11'b11111111101;
        x_t[35] = 11'b11111111101;
        x_t[36] = 11'b11111111000;
        x_t[37] = 11'b00000000110;
        x_t[38] = 11'b11111111001;
        x_t[39] = 11'b00000000000;
        x_t[40] = 11'b00000000000;
        x_t[41] = 11'b11111011010;
        x_t[42] = 11'b11111101101;
        x_t[43] = 11'b00000010000;
        x_t[44] = 11'b11111101100;
        x_t[45] = 11'b00000100001;
        x_t[46] = 11'b00000000011;
        x_t[47] = 11'b00000000011;
        x_t[48] = 11'b00000000111;
        x_t[49] = 11'b00000001000;
        x_t[50] = 11'b00000001011;
        x_t[51] = 11'b00000001111;
        x_t[52] = 11'b00000001100;
        x_t[53] = 11'b00000001100;
        x_t[54] = 11'b00000001101;
        x_t[55] = 11'b00000001001;
        x_t[56] = 11'b00000000110;
        x_t[57] = 11'b00000010001;
        x_t[58] = 11'b00000010010;
        x_t[59] = 11'b00000011000;
        x_t[60] = 11'b00000010111;
        x_t[61] = 11'b00000100000;
        x_t[62] = 11'b00000001010;
        x_t[63] = 11'b00000010010;
        
        h_t_prev[0] = 11'b00000000101;
        h_t_prev[1] = 11'b00000000110;
        h_t_prev[2] = 11'b00000000001;
        h_t_prev[3] = 11'b00000001010;
        h_t_prev[4] = 11'b00000001101;
        h_t_prev[5] = 11'b00000000000;
        h_t_prev[6] = 11'b11111111110;
        h_t_prev[7] = 11'b11111111011;
        h_t_prev[8] = 11'b00000000011;
        h_t_prev[9] = 11'b00000001001;
        h_t_prev[10] = 11'b00000001101;
        h_t_prev[11] = 11'b00000000011;
        h_t_prev[12] = 11'b00000000110;
        h_t_prev[13] = 11'b00000000111;
        h_t_prev[14] = 11'b00000000110;
        h_t_prev[15] = 11'b00000000100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 82 timeout!");
                $fdisplay(fd_cycles, "Test Vector  82: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  82: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 82");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 83
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111111011;
        x_t[1] = 11'b00000000000;
        x_t[2] = 11'b00000000000;
        x_t[3] = 11'b00000001100;
        x_t[4] = 11'b00000001110;
        x_t[5] = 11'b00000000000;
        x_t[6] = 11'b11111111010;
        x_t[7] = 11'b11111101111;
        x_t[8] = 11'b11111111010;
        x_t[9] = 11'b00000000101;
        x_t[10] = 11'b00000001111;
        x_t[11] = 11'b00000000000;
        x_t[12] = 11'b00000000011;
        x_t[13] = 11'b00000000110;
        x_t[14] = 11'b11111110111;
        x_t[15] = 11'b11111111110;
        x_t[16] = 11'b00000000010;
        x_t[17] = 11'b00000000100;
        x_t[18] = 11'b00000000100;
        x_t[19] = 11'b00000000101;
        x_t[20] = 11'b11111111111;
        x_t[21] = 11'b11111111101;
        x_t[22] = 11'b11111111110;
        x_t[23] = 11'b11111111000;
        x_t[24] = 11'b11111101101;
        x_t[25] = 11'b11111101110;
        x_t[26] = 11'b11111110100;
        x_t[27] = 11'b11111110101;
        x_t[28] = 11'b11111111110;
        x_t[29] = 11'b11111110010;
        x_t[30] = 11'b11111101001;
        x_t[31] = 11'b11111101110;
        x_t[32] = 11'b11111110011;
        x_t[33] = 11'b11111110101;
        x_t[34] = 11'b11111110000;
        x_t[35] = 11'b11111101110;
        x_t[36] = 11'b11111101000;
        x_t[37] = 11'b11111111000;
        x_t[38] = 11'b11111100111;
        x_t[39] = 11'b11111111010;
        x_t[40] = 11'b11111100101;
        x_t[41] = 11'b11111100100;
        x_t[42] = 11'b11111100010;
        x_t[43] = 11'b11111111110;
        x_t[44] = 11'b11111100000;
        x_t[45] = 11'b00000011111;
        x_t[46] = 11'b11111111000;
        x_t[47] = 11'b11111111100;
        x_t[48] = 11'b00000000000;
        x_t[49] = 11'b00000000010;
        x_t[50] = 11'b00000000011;
        x_t[51] = 11'b00000000101;
        x_t[52] = 11'b00000000010;
        x_t[53] = 11'b00000000101;
        x_t[54] = 11'b00000001101;
        x_t[55] = 11'b00000001010;
        x_t[56] = 11'b00000000011;
        x_t[57] = 11'b00000001001;
        x_t[58] = 11'b00000001011;
        x_t[59] = 11'b00000011000;
        x_t[60] = 11'b00000010101;
        x_t[61] = 11'b00000011100;
        x_t[62] = 11'b00000000010;
        x_t[63] = 11'b00000010001;
        
        h_t_prev[0] = 11'b11111111011;
        h_t_prev[1] = 11'b00000000000;
        h_t_prev[2] = 11'b00000000000;
        h_t_prev[3] = 11'b00000001100;
        h_t_prev[4] = 11'b00000001110;
        h_t_prev[5] = 11'b00000000000;
        h_t_prev[6] = 11'b11111111010;
        h_t_prev[7] = 11'b11111101111;
        h_t_prev[8] = 11'b11111111010;
        h_t_prev[9] = 11'b00000000101;
        h_t_prev[10] = 11'b00000001111;
        h_t_prev[11] = 11'b00000000000;
        h_t_prev[12] = 11'b00000000011;
        h_t_prev[13] = 11'b00000000110;
        h_t_prev[14] = 11'b11111110111;
        h_t_prev[15] = 11'b11111111110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 83 timeout!");
                $fdisplay(fd_cycles, "Test Vector  83: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  83: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 83");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 84
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111101101;
        x_t[1] = 11'b11111110011;
        x_t[2] = 11'b11111110010;
        x_t[3] = 11'b11111111100;
        x_t[4] = 11'b11111111110;
        x_t[5] = 11'b11111110000;
        x_t[6] = 11'b11111101001;
        x_t[7] = 11'b11111100001;
        x_t[8] = 11'b11111110000;
        x_t[9] = 11'b11111111010;
        x_t[10] = 11'b00000000100;
        x_t[11] = 11'b11111101110;
        x_t[12] = 11'b11111110101;
        x_t[13] = 11'b11111111110;
        x_t[14] = 11'b11111110111;
        x_t[15] = 11'b11111111101;
        x_t[16] = 11'b11111111011;
        x_t[17] = 11'b11111111010;
        x_t[18] = 11'b11111110110;
        x_t[19] = 11'b11111111000;
        x_t[20] = 11'b11111110011;
        x_t[21] = 11'b11111111010;
        x_t[22] = 11'b11111111000;
        x_t[23] = 11'b11111110001;
        x_t[24] = 11'b11111101100;
        x_t[25] = 11'b11111101100;
        x_t[26] = 11'b11111101111;
        x_t[27] = 11'b11111101101;
        x_t[28] = 11'b11111110101;
        x_t[29] = 11'b11111110100;
        x_t[30] = 11'b11111101011;
        x_t[31] = 11'b11111100101;
        x_t[32] = 11'b11111110000;
        x_t[33] = 11'b11111101110;
        x_t[34] = 11'b11111101001;
        x_t[35] = 11'b11111101011;
        x_t[36] = 11'b11111100010;
        x_t[37] = 11'b11111110010;
        x_t[38] = 11'b11111110000;
        x_t[39] = 11'b00000000011;
        x_t[40] = 11'b11111111011;
        x_t[41] = 11'b11111111101;
        x_t[42] = 11'b11111110010;
        x_t[43] = 11'b11111101100;
        x_t[44] = 11'b11111101010;
        x_t[45] = 11'b00000001110;
        x_t[46] = 11'b00000000010;
        x_t[47] = 11'b00000000001;
        x_t[48] = 11'b11111111100;
        x_t[49] = 11'b11111111111;
        x_t[50] = 11'b11111111001;
        x_t[51] = 11'b11111111000;
        x_t[52] = 11'b11111110100;
        x_t[53] = 11'b11111110111;
        x_t[54] = 11'b00000000111;
        x_t[55] = 11'b00000001110;
        x_t[56] = 11'b00000000010;
        x_t[57] = 11'b11111111111;
        x_t[58] = 11'b00000000011;
        x_t[59] = 11'b00000011000;
        x_t[60] = 11'b00000010101;
        x_t[61] = 11'b00000011010;
        x_t[62] = 11'b00000000000;
        x_t[63] = 11'b00000010001;
        
        h_t_prev[0] = 11'b11111101101;
        h_t_prev[1] = 11'b11111110011;
        h_t_prev[2] = 11'b11111110010;
        h_t_prev[3] = 11'b11111111100;
        h_t_prev[4] = 11'b11111111110;
        h_t_prev[5] = 11'b11111110000;
        h_t_prev[6] = 11'b11111101001;
        h_t_prev[7] = 11'b11111100001;
        h_t_prev[8] = 11'b11111110000;
        h_t_prev[9] = 11'b11111111010;
        h_t_prev[10] = 11'b00000000100;
        h_t_prev[11] = 11'b11111101110;
        h_t_prev[12] = 11'b11111110101;
        h_t_prev[13] = 11'b11111111110;
        h_t_prev[14] = 11'b11111110111;
        h_t_prev[15] = 11'b11111111101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 84 timeout!");
                $fdisplay(fd_cycles, "Test Vector  84: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  84: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 84");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 85
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111110101;
        x_t[1] = 11'b11111111010;
        x_t[2] = 11'b11111110000;
        x_t[3] = 11'b11111110110;
        x_t[4] = 11'b11111110110;
        x_t[5] = 11'b11111101011;
        x_t[6] = 11'b11111101011;
        x_t[7] = 11'b11111101100;
        x_t[8] = 11'b11111110101;
        x_t[9] = 11'b11111110111;
        x_t[10] = 11'b11111111100;
        x_t[11] = 11'b11111101000;
        x_t[12] = 11'b11111101011;
        x_t[13] = 11'b11111111001;
        x_t[14] = 11'b11111111011;
        x_t[15] = 11'b11111111101;
        x_t[16] = 11'b11111110111;
        x_t[17] = 11'b11111110001;
        x_t[18] = 11'b11111101001;
        x_t[19] = 11'b11111101010;
        x_t[20] = 11'b11111100101;
        x_t[21] = 11'b11111110110;
        x_t[22] = 11'b11111110011;
        x_t[23] = 11'b11111101101;
        x_t[24] = 11'b11111101000;
        x_t[25] = 11'b11111101000;
        x_t[26] = 11'b11111101000;
        x_t[27] = 11'b11111101001;
        x_t[28] = 11'b11111110011;
        x_t[29] = 11'b11111101011;
        x_t[30] = 11'b11111100110;
        x_t[31] = 11'b11111100100;
        x_t[32] = 11'b11111101101;
        x_t[33] = 11'b11111101000;
        x_t[34] = 11'b11111100011;
        x_t[35] = 11'b11111100101;
        x_t[36] = 11'b11111100000;
        x_t[37] = 11'b11111101110;
        x_t[38] = 11'b11111101010;
        x_t[39] = 11'b11111110111;
        x_t[40] = 11'b11111101101;
        x_t[41] = 11'b11111100100;
        x_t[42] = 11'b11111100111;
        x_t[43] = 11'b00000010000;
        x_t[44] = 11'b11111101011;
        x_t[45] = 11'b00000001001;
        x_t[46] = 11'b00000000010;
        x_t[47] = 11'b00000000000;
        x_t[48] = 11'b11111111000;
        x_t[49] = 11'b11111111011;
        x_t[50] = 11'b11111110001;
        x_t[51] = 11'b11111110000;
        x_t[52] = 11'b11111101100;
        x_t[53] = 11'b11111110100;
        x_t[54] = 11'b00000000101;
        x_t[55] = 11'b00000000111;
        x_t[56] = 11'b11111111101;
        x_t[57] = 11'b11111110110;
        x_t[58] = 11'b11111111110;
        x_t[59] = 11'b00000011010;
        x_t[60] = 11'b00000010011;
        x_t[61] = 11'b00000010111;
        x_t[62] = 11'b00000000100;
        x_t[63] = 11'b00000010001;
        
        h_t_prev[0] = 11'b11111110101;
        h_t_prev[1] = 11'b11111111010;
        h_t_prev[2] = 11'b11111110000;
        h_t_prev[3] = 11'b11111110110;
        h_t_prev[4] = 11'b11111110110;
        h_t_prev[5] = 11'b11111101011;
        h_t_prev[6] = 11'b11111101011;
        h_t_prev[7] = 11'b11111101100;
        h_t_prev[8] = 11'b11111110101;
        h_t_prev[9] = 11'b11111110111;
        h_t_prev[10] = 11'b11111111100;
        h_t_prev[11] = 11'b11111101000;
        h_t_prev[12] = 11'b11111101011;
        h_t_prev[13] = 11'b11111111001;
        h_t_prev[14] = 11'b11111111011;
        h_t_prev[15] = 11'b11111111101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 85 timeout!");
                $fdisplay(fd_cycles, "Test Vector  85: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  85: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 85");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 86
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111110101;
        x_t[1] = 11'b11111111010;
        x_t[2] = 11'b11111110011;
        x_t[3] = 11'b11111110101;
        x_t[4] = 11'b11111111010;
        x_t[5] = 11'b11111110000;
        x_t[6] = 11'b11111101101;
        x_t[7] = 11'b11111110011;
        x_t[8] = 11'b11111111010;
        x_t[9] = 11'b11111111100;
        x_t[10] = 11'b11111111110;
        x_t[11] = 11'b11111101101;
        x_t[12] = 11'b11111110000;
        x_t[13] = 11'b11111111001;
        x_t[14] = 11'b00000000010;
        x_t[15] = 11'b00000000100;
        x_t[16] = 11'b11111111011;
        x_t[17] = 11'b11111110100;
        x_t[18] = 11'b11111101100;
        x_t[19] = 11'b11111101101;
        x_t[20] = 11'b11111101000;
        x_t[21] = 11'b11111111100;
        x_t[22] = 11'b11111110110;
        x_t[23] = 11'b11111101110;
        x_t[24] = 11'b11111101110;
        x_t[25] = 11'b11111101110;
        x_t[26] = 11'b11111101111;
        x_t[27] = 11'b11111101110;
        x_t[28] = 11'b11111110011;
        x_t[29] = 11'b11111110110;
        x_t[30] = 11'b11111101111;
        x_t[31] = 11'b11111101110;
        x_t[32] = 11'b11111110110;
        x_t[33] = 11'b11111110010;
        x_t[34] = 11'b11111101101;
        x_t[35] = 11'b11111110000;
        x_t[36] = 11'b11111101011;
        x_t[37] = 11'b11111110100;
        x_t[38] = 11'b11111110101;
        x_t[39] = 11'b00000000000;
        x_t[40] = 11'b11111111110;
        x_t[41] = 11'b11111011111;
        x_t[42] = 11'b11111111110;
        x_t[43] = 11'b00000010000;
        x_t[44] = 11'b11111111010;
        x_t[45] = 11'b00000010010;
        x_t[46] = 11'b00000001001;
        x_t[47] = 11'b00000000101;
        x_t[48] = 11'b11111111101;
        x_t[49] = 11'b11111111101;
        x_t[50] = 11'b11111110010;
        x_t[51] = 11'b11111110001;
        x_t[52] = 11'b11111101110;
        x_t[53] = 11'b11111110111;
        x_t[54] = 11'b00000000010;
        x_t[55] = 11'b00000000110;
        x_t[56] = 11'b11111111100;
        x_t[57] = 11'b11111110011;
        x_t[58] = 11'b11111111100;
        x_t[59] = 11'b00000010011;
        x_t[60] = 11'b00000010000;
        x_t[61] = 11'b00000010010;
        x_t[62] = 11'b00000000101;
        x_t[63] = 11'b00000001101;
        
        h_t_prev[0] = 11'b11111110101;
        h_t_prev[1] = 11'b11111111010;
        h_t_prev[2] = 11'b11111110011;
        h_t_prev[3] = 11'b11111110101;
        h_t_prev[4] = 11'b11111111010;
        h_t_prev[5] = 11'b11111110000;
        h_t_prev[6] = 11'b11111101101;
        h_t_prev[7] = 11'b11111110011;
        h_t_prev[8] = 11'b11111111010;
        h_t_prev[9] = 11'b11111111100;
        h_t_prev[10] = 11'b11111111110;
        h_t_prev[11] = 11'b11111101101;
        h_t_prev[12] = 11'b11111110000;
        h_t_prev[13] = 11'b11111111001;
        h_t_prev[14] = 11'b00000000010;
        h_t_prev[15] = 11'b00000000100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 86 timeout!");
                $fdisplay(fd_cycles, "Test Vector  86: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  86: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 86");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 87
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000000001;
        x_t[1] = 11'b00000000011;
        x_t[2] = 11'b11111111010;
        x_t[3] = 11'b11111111011;
        x_t[4] = 11'b00000000010;
        x_t[5] = 11'b11111111110;
        x_t[6] = 11'b11111111111;
        x_t[7] = 11'b11111111011;
        x_t[8] = 11'b00000000000;
        x_t[9] = 11'b00000000010;
        x_t[10] = 11'b00000000100;
        x_t[11] = 11'b11111110100;
        x_t[12] = 11'b11111111111;
        x_t[13] = 11'b00000001001;
        x_t[14] = 11'b00000001001;
        x_t[15] = 11'b00000000111;
        x_t[16] = 11'b00000000000;
        x_t[17] = 11'b11111111001;
        x_t[18] = 11'b11111110110;
        x_t[19] = 11'b11111111001;
        x_t[20] = 11'b11111110101;
        x_t[21] = 11'b00000000111;
        x_t[22] = 11'b00000000011;
        x_t[23] = 11'b11111111010;
        x_t[24] = 11'b11111111010;
        x_t[25] = 11'b11111111001;
        x_t[26] = 11'b11111110110;
        x_t[27] = 11'b11111111011;
        x_t[28] = 11'b11111111111;
        x_t[29] = 11'b00000000101;
        x_t[30] = 11'b11111111011;
        x_t[31] = 11'b11111110011;
        x_t[32] = 11'b11111111010;
        x_t[33] = 11'b11111110101;
        x_t[34] = 11'b11111110011;
        x_t[35] = 11'b11111111000;
        x_t[36] = 11'b11111111000;
        x_t[37] = 11'b11111111111;
        x_t[38] = 11'b00000000001;
        x_t[39] = 11'b00000010110;
        x_t[40] = 11'b00000010000;
        x_t[41] = 11'b00000000101;
        x_t[42] = 11'b00000000111;
        x_t[43] = 11'b00000010001;
        x_t[44] = 11'b11111111110;
        x_t[45] = 11'b00000011001;
        x_t[46] = 11'b00000001101;
        x_t[47] = 11'b00000001011;
        x_t[48] = 11'b00000000010;
        x_t[49] = 11'b11111111111;
        x_t[50] = 11'b11111110111;
        x_t[51] = 11'b11111110010;
        x_t[52] = 11'b11111110010;
        x_t[53] = 11'b11111111010;
        x_t[54] = 11'b11111111111;
        x_t[55] = 11'b00000001001;
        x_t[56] = 11'b00000000010;
        x_t[57] = 11'b11111110101;
        x_t[58] = 11'b11111110110;
        x_t[59] = 11'b00000000110;
        x_t[60] = 11'b00000001001;
        x_t[61] = 11'b00000000101;
        x_t[62] = 11'b11111111001;
        x_t[63] = 11'b11111111111;
        
        h_t_prev[0] = 11'b00000000001;
        h_t_prev[1] = 11'b00000000011;
        h_t_prev[2] = 11'b11111111010;
        h_t_prev[3] = 11'b11111111011;
        h_t_prev[4] = 11'b00000000010;
        h_t_prev[5] = 11'b11111111110;
        h_t_prev[6] = 11'b11111111111;
        h_t_prev[7] = 11'b11111111011;
        h_t_prev[8] = 11'b00000000000;
        h_t_prev[9] = 11'b00000000010;
        h_t_prev[10] = 11'b00000000100;
        h_t_prev[11] = 11'b11111110100;
        h_t_prev[12] = 11'b11111111111;
        h_t_prev[13] = 11'b00000001001;
        h_t_prev[14] = 11'b00000001001;
        h_t_prev[15] = 11'b00000000111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 87 timeout!");
                $fdisplay(fd_cycles, "Test Vector  87: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  87: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 87");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 88
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000001000;
        x_t[1] = 11'b00000001000;
        x_t[2] = 11'b11111111111;
        x_t[3] = 11'b00000000000;
        x_t[4] = 11'b00000000100;
        x_t[5] = 11'b00000000000;
        x_t[6] = 11'b00000000000;
        x_t[7] = 11'b00000000100;
        x_t[8] = 11'b00000000111;
        x_t[9] = 11'b00000001010;
        x_t[10] = 11'b00000010001;
        x_t[11] = 11'b11111111011;
        x_t[12] = 11'b00000000111;
        x_t[13] = 11'b00000001110;
        x_t[14] = 11'b00000010101;
        x_t[15] = 11'b00000010000;
        x_t[16] = 11'b00000001000;
        x_t[17] = 11'b00000000010;
        x_t[18] = 11'b11111111110;
        x_t[19] = 11'b00000000010;
        x_t[20] = 11'b11111111110;
        x_t[21] = 11'b11111111111;
        x_t[22] = 11'b00000000000;
        x_t[23] = 11'b11111111000;
        x_t[24] = 11'b11111110110;
        x_t[25] = 11'b11111110101;
        x_t[26] = 11'b11111110001;
        x_t[27] = 11'b11111111000;
        x_t[28] = 11'b00000000000;
        x_t[29] = 11'b00000000000;
        x_t[30] = 11'b11111110101;
        x_t[31] = 11'b11111110001;
        x_t[32] = 11'b11111111000;
        x_t[33] = 11'b11111110010;
        x_t[34] = 11'b11111101101;
        x_t[35] = 11'b11111110001;
        x_t[36] = 11'b11111110000;
        x_t[37] = 11'b11111110010;
        x_t[38] = 11'b00000000000;
        x_t[39] = 11'b00000001011;
        x_t[40] = 11'b00000011000;
        x_t[41] = 11'b11111101110;
        x_t[42] = 11'b11111110001;
        x_t[43] = 11'b00000011110;
        x_t[44] = 11'b00000000101;
        x_t[45] = 11'b00000011011;
        x_t[46] = 11'b00000011101;
        x_t[47] = 11'b00000011010;
        x_t[48] = 11'b00000001101;
        x_t[49] = 11'b00000001101;
        x_t[50] = 11'b00000000010;
        x_t[51] = 11'b11111110101;
        x_t[52] = 11'b11111110100;
        x_t[53] = 11'b11111111010;
        x_t[54] = 11'b11111111011;
        x_t[55] = 11'b00000010010;
        x_t[56] = 11'b00000010000;
        x_t[57] = 11'b11111111010;
        x_t[58] = 11'b11111101101;
        x_t[59] = 11'b11111111000;
        x_t[60] = 11'b00000001001;
        x_t[61] = 11'b11111111001;
        x_t[62] = 11'b11111100101;
        x_t[63] = 11'b11111110110;
        
        h_t_prev[0] = 11'b00000001000;
        h_t_prev[1] = 11'b00000001000;
        h_t_prev[2] = 11'b11111111111;
        h_t_prev[3] = 11'b00000000000;
        h_t_prev[4] = 11'b00000000100;
        h_t_prev[5] = 11'b00000000000;
        h_t_prev[6] = 11'b00000000000;
        h_t_prev[7] = 11'b00000000100;
        h_t_prev[8] = 11'b00000000111;
        h_t_prev[9] = 11'b00000001010;
        h_t_prev[10] = 11'b00000010001;
        h_t_prev[11] = 11'b11111111011;
        h_t_prev[12] = 11'b00000000111;
        h_t_prev[13] = 11'b00000001110;
        h_t_prev[14] = 11'b00000010101;
        h_t_prev[15] = 11'b00000010000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 88 timeout!");
                $fdisplay(fd_cycles, "Test Vector  88: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  88: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 88");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 89
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000001011;
        x_t[1] = 11'b00000001001;
        x_t[2] = 11'b00000000001;
        x_t[3] = 11'b00000000110;
        x_t[4] = 11'b00000001001;
        x_t[5] = 11'b00000000000;
        x_t[6] = 11'b11111110101;
        x_t[7] = 11'b00000001000;
        x_t[8] = 11'b00000000111;
        x_t[9] = 11'b00000001100;
        x_t[10] = 11'b00000010101;
        x_t[11] = 11'b00000000000;
        x_t[12] = 11'b00000001011;
        x_t[13] = 11'b00000001111;
        x_t[14] = 11'b00000010110;
        x_t[15] = 11'b00000001111;
        x_t[16] = 11'b00000001100;
        x_t[17] = 11'b00000001001;
        x_t[18] = 11'b00000000010;
        x_t[19] = 11'b00000000011;
        x_t[20] = 11'b11111111111;
        x_t[21] = 11'b11111111011;
        x_t[22] = 11'b11111111101;
        x_t[23] = 11'b11111110101;
        x_t[24] = 11'b11111110101;
        x_t[25] = 11'b11111110100;
        x_t[26] = 11'b11111110011;
        x_t[27] = 11'b11111110100;
        x_t[28] = 11'b11111111010;
        x_t[29] = 11'b00000000000;
        x_t[30] = 11'b11111110011;
        x_t[31] = 11'b11111110010;
        x_t[32] = 11'b11111111110;
        x_t[33] = 11'b11111111000;
        x_t[34] = 11'b11111110001;
        x_t[35] = 11'b11111110111;
        x_t[36] = 11'b11111101110;
        x_t[37] = 11'b11111101100;
        x_t[38] = 11'b00000000100;
        x_t[39] = 11'b00000000001;
        x_t[40] = 11'b00000001010;
        x_t[41] = 11'b11111011010;
        x_t[42] = 11'b11111110011;
        x_t[43] = 11'b00000010000;
        x_t[44] = 11'b11111110111;
        x_t[45] = 11'b00000001101;
        x_t[46] = 11'b00000001010;
        x_t[47] = 11'b00000001110;
        x_t[48] = 11'b00000000110;
        x_t[49] = 11'b00000001001;
        x_t[50] = 11'b11111111110;
        x_t[51] = 11'b11111101011;
        x_t[52] = 11'b11111101010;
        x_t[53] = 11'b11111100111;
        x_t[54] = 11'b11111100101;
        x_t[55] = 11'b00000000011;
        x_t[56] = 11'b00000000110;
        x_t[57] = 11'b11111101110;
        x_t[58] = 11'b11111010100;
        x_t[59] = 11'b11111010011;
        x_t[60] = 11'b00000000000;
        x_t[61] = 11'b11111100111;
        x_t[62] = 11'b11111000110;
        x_t[63] = 11'b11111100011;
        
        h_t_prev[0] = 11'b00000001011;
        h_t_prev[1] = 11'b00000001001;
        h_t_prev[2] = 11'b00000000001;
        h_t_prev[3] = 11'b00000000110;
        h_t_prev[4] = 11'b00000001001;
        h_t_prev[5] = 11'b00000000000;
        h_t_prev[6] = 11'b11111110101;
        h_t_prev[7] = 11'b00000001000;
        h_t_prev[8] = 11'b00000000111;
        h_t_prev[9] = 11'b00000001100;
        h_t_prev[10] = 11'b00000010101;
        h_t_prev[11] = 11'b00000000000;
        h_t_prev[12] = 11'b00000001011;
        h_t_prev[13] = 11'b00000001111;
        h_t_prev[14] = 11'b00000010110;
        h_t_prev[15] = 11'b00000001111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 89 timeout!");
                $fdisplay(fd_cycles, "Test Vector  89: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  89: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 89");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 90
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000001110;
        x_t[1] = 11'b00000001110;
        x_t[2] = 11'b00000001001;
        x_t[3] = 11'b00000001111;
        x_t[4] = 11'b00000010101;
        x_t[5] = 11'b00000001011;
        x_t[6] = 11'b00000000000;
        x_t[7] = 11'b00000000000;
        x_t[8] = 11'b00000000101;
        x_t[9] = 11'b00000001111;
        x_t[10] = 11'b00000011100;
        x_t[11] = 11'b00000001101;
        x_t[12] = 11'b00000001110;
        x_t[13] = 11'b00000001110;
        x_t[14] = 11'b00000000100;
        x_t[15] = 11'b00000000111;
        x_t[16] = 11'b00000001010;
        x_t[17] = 11'b00000001010;
        x_t[18] = 11'b00000000011;
        x_t[19] = 11'b11111111111;
        x_t[20] = 11'b11111111000;
        x_t[21] = 11'b00000000011;
        x_t[22] = 11'b00000000101;
        x_t[23] = 11'b11111111110;
        x_t[24] = 11'b11111111001;
        x_t[25] = 11'b11111111000;
        x_t[26] = 11'b00000000000;
        x_t[27] = 11'b00000000010;
        x_t[28] = 11'b00000000110;
        x_t[29] = 11'b11111111011;
        x_t[30] = 11'b11111111010;
        x_t[31] = 11'b11111111111;
        x_t[32] = 11'b00000001000;
        x_t[33] = 11'b00000001000;
        x_t[34] = 11'b00000000000;
        x_t[35] = 11'b00000000011;
        x_t[36] = 11'b00000000010;
        x_t[37] = 11'b00000000100;
        x_t[38] = 11'b11111111110;
        x_t[39] = 11'b00000011000;
        x_t[40] = 11'b11111111110;
        x_t[41] = 11'b11111100011;
        x_t[42] = 11'b11111100111;
        x_t[43] = 11'b00000000001;
        x_t[44] = 11'b11111100111;
        x_t[45] = 11'b00000000101;
        x_t[46] = 11'b11111110011;
        x_t[47] = 11'b11111111010;
        x_t[48] = 11'b11111110111;
        x_t[49] = 11'b11111111111;
        x_t[50] = 11'b11111111001;
        x_t[51] = 11'b11111100001;
        x_t[52] = 11'b11111011111;
        x_t[53] = 11'b11111010110;
        x_t[54] = 11'b11111010000;
        x_t[55] = 11'b11111101111;
        x_t[56] = 11'b11111110010;
        x_t[57] = 11'b11111100001;
        x_t[58] = 11'b11111000011;
        x_t[59] = 11'b11110110100;
        x_t[60] = 11'b11111101011;
        x_t[61] = 11'b11111001100;
        x_t[62] = 11'b11110100011;
        x_t[63] = 11'b11111000110;
        
        h_t_prev[0] = 11'b00000001110;
        h_t_prev[1] = 11'b00000001110;
        h_t_prev[2] = 11'b00000001001;
        h_t_prev[3] = 11'b00000001111;
        h_t_prev[4] = 11'b00000010101;
        h_t_prev[5] = 11'b00000001011;
        h_t_prev[6] = 11'b00000000000;
        h_t_prev[7] = 11'b00000000000;
        h_t_prev[8] = 11'b00000000101;
        h_t_prev[9] = 11'b00000001111;
        h_t_prev[10] = 11'b00000011100;
        h_t_prev[11] = 11'b00000001101;
        h_t_prev[12] = 11'b00000001110;
        h_t_prev[13] = 11'b00000001110;
        h_t_prev[14] = 11'b00000000100;
        h_t_prev[15] = 11'b00000000111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 90 timeout!");
                $fdisplay(fd_cycles, "Test Vector  90: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  90: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 90");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 91
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000001001;
        x_t[1] = 11'b00000010010;
        x_t[2] = 11'b00000010101;
        x_t[3] = 11'b00000011101;
        x_t[4] = 11'b00000011101;
        x_t[5] = 11'b00000010001;
        x_t[6] = 11'b00000001011;
        x_t[7] = 11'b00000000000;
        x_t[8] = 11'b00000001000;
        x_t[9] = 11'b00000011000;
        x_t[10] = 11'b00000100110;
        x_t[11] = 11'b00000001111;
        x_t[12] = 11'b00000001100;
        x_t[13] = 11'b00000001010;
        x_t[14] = 11'b11111111011;
        x_t[15] = 11'b00000001000;
        x_t[16] = 11'b00000001100;
        x_t[17] = 11'b00000001100;
        x_t[18] = 11'b00000000100;
        x_t[19] = 11'b11111111101;
        x_t[20] = 11'b11111110001;
        x_t[21] = 11'b00000000111;
        x_t[22] = 11'b00000001000;
        x_t[23] = 11'b00000000010;
        x_t[24] = 11'b11111111011;
        x_t[25] = 11'b11111111011;
        x_t[26] = 11'b00000000111;
        x_t[27] = 11'b00000000110;
        x_t[28] = 11'b00000001010;
        x_t[29] = 11'b11111111011;
        x_t[30] = 11'b11111111111;
        x_t[31] = 11'b00000000101;
        x_t[32] = 11'b00000010000;
        x_t[33] = 11'b00000010001;
        x_t[34] = 11'b00000001010;
        x_t[35] = 11'b00000001010;
        x_t[36] = 11'b00000000101;
        x_t[37] = 11'b00000000001;
        x_t[38] = 11'b11111111010;
        x_t[39] = 11'b00000011001;
        x_t[40] = 11'b11111110110;
        x_t[41] = 11'b11111111110;
        x_t[42] = 11'b11111110111;
        x_t[43] = 11'b00000011110;
        x_t[44] = 11'b11111110101;
        x_t[45] = 11'b00000000011;
        x_t[46] = 11'b11111110111;
        x_t[47] = 11'b11111111100;
        x_t[48] = 11'b11111111010;
        x_t[49] = 11'b00000000111;
        x_t[50] = 11'b00000000100;
        x_t[51] = 11'b11111101110;
        x_t[52] = 11'b11111101011;
        x_t[53] = 11'b11111100011;
        x_t[54] = 11'b11111011010;
        x_t[55] = 11'b11111110010;
        x_t[56] = 11'b11111110110;
        x_t[57] = 11'b11111101111;
        x_t[58] = 11'b11111010011;
        x_t[59] = 11'b11111000111;
        x_t[60] = 11'b11111011110;
        x_t[61] = 11'b11111000000;
        x_t[62] = 11'b11110010111;
        x_t[63] = 11'b11110111110;
        
        h_t_prev[0] = 11'b00000001001;
        h_t_prev[1] = 11'b00000010010;
        h_t_prev[2] = 11'b00000010101;
        h_t_prev[3] = 11'b00000011101;
        h_t_prev[4] = 11'b00000011101;
        h_t_prev[5] = 11'b00000010001;
        h_t_prev[6] = 11'b00000001011;
        h_t_prev[7] = 11'b00000000000;
        h_t_prev[8] = 11'b00000001000;
        h_t_prev[9] = 11'b00000011000;
        h_t_prev[10] = 11'b00000100110;
        h_t_prev[11] = 11'b00000001111;
        h_t_prev[12] = 11'b00000001100;
        h_t_prev[13] = 11'b00000001010;
        h_t_prev[14] = 11'b11111111011;
        h_t_prev[15] = 11'b00000001000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 91 timeout!");
                $fdisplay(fd_cycles, "Test Vector  91: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  91: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 91");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 92
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000001110;
        x_t[1] = 11'b00000011011;
        x_t[2] = 11'b00000011111;
        x_t[3] = 11'b00000100101;
        x_t[4] = 11'b00000100001;
        x_t[5] = 11'b00000010100;
        x_t[6] = 11'b00000001011;
        x_t[7] = 11'b00000000001;
        x_t[8] = 11'b00000010101;
        x_t[9] = 11'b00000100110;
        x_t[10] = 11'b00000110010;
        x_t[11] = 11'b00000010011;
        x_t[12] = 11'b00000010001;
        x_t[13] = 11'b00000010110;
        x_t[14] = 11'b00000000111;
        x_t[15] = 11'b00000010110;
        x_t[16] = 11'b00000011101;
        x_t[17] = 11'b00000011100;
        x_t[18] = 11'b00000010000;
        x_t[19] = 11'b00000000111;
        x_t[20] = 11'b11111111011;
        x_t[21] = 11'b00000001011;
        x_t[22] = 11'b00000001001;
        x_t[23] = 11'b11111111110;
        x_t[24] = 11'b00000000101;
        x_t[25] = 11'b00000000100;
        x_t[26] = 11'b00000000110;
        x_t[27] = 11'b00000000011;
        x_t[28] = 11'b00000000110;
        x_t[29] = 11'b00000010010;
        x_t[30] = 11'b11111111101;
        x_t[31] = 11'b00000000100;
        x_t[32] = 11'b00000010001;
        x_t[33] = 11'b00000001111;
        x_t[34] = 11'b00000001011;
        x_t[35] = 11'b00000001011;
        x_t[36] = 11'b00000000010;
        x_t[37] = 11'b11111110101;
        x_t[38] = 11'b00000001110;
        x_t[39] = 11'b00000011001;
        x_t[40] = 11'b00000010101;
        x_t[41] = 11'b11111111100;
        x_t[42] = 11'b00000010001;
        x_t[43] = 11'b00000001000;
        x_t[44] = 11'b00000000110;
        x_t[45] = 11'b00000000011;
        x_t[46] = 11'b00000000101;
        x_t[47] = 11'b00000001010;
        x_t[48] = 11'b00000000101;
        x_t[49] = 11'b00000010100;
        x_t[50] = 11'b00000010101;
        x_t[51] = 11'b00000000000;
        x_t[52] = 11'b11111111011;
        x_t[53] = 11'b11111110000;
        x_t[54] = 11'b11111100011;
        x_t[55] = 11'b11111111001;
        x_t[56] = 11'b00000000000;
        x_t[57] = 11'b00000000001;
        x_t[58] = 11'b11111101001;
        x_t[59] = 11'b11111011100;
        x_t[60] = 11'b11111100001;
        x_t[61] = 11'b11111001101;
        x_t[62] = 11'b11110100111;
        x_t[63] = 11'b11110111111;
        
        h_t_prev[0] = 11'b00000001110;
        h_t_prev[1] = 11'b00000011011;
        h_t_prev[2] = 11'b00000011111;
        h_t_prev[3] = 11'b00000100101;
        h_t_prev[4] = 11'b00000100001;
        h_t_prev[5] = 11'b00000010100;
        h_t_prev[6] = 11'b00000001011;
        h_t_prev[7] = 11'b00000000001;
        h_t_prev[8] = 11'b00000010101;
        h_t_prev[9] = 11'b00000100110;
        h_t_prev[10] = 11'b00000110010;
        h_t_prev[11] = 11'b00000010011;
        h_t_prev[12] = 11'b00000010001;
        h_t_prev[13] = 11'b00000010110;
        h_t_prev[14] = 11'b00000000111;
        h_t_prev[15] = 11'b00000010110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 92 timeout!");
                $fdisplay(fd_cycles, "Test Vector  92: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  92: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 92");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 93
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000011010;
        x_t[1] = 11'b00000100110;
        x_t[2] = 11'b00000100111;
        x_t[3] = 11'b00000101011;
        x_t[4] = 11'b00000100111;
        x_t[5] = 11'b00000011011;
        x_t[6] = 11'b00000010010;
        x_t[7] = 11'b00000010110;
        x_t[8] = 11'b00000100111;
        x_t[9] = 11'b00000110101;
        x_t[10] = 11'b00001000010;
        x_t[11] = 11'b00000100110;
        x_t[12] = 11'b00000011101;
        x_t[13] = 11'b00000011100;
        x_t[14] = 11'b00000100000;
        x_t[15] = 11'b00000101101;
        x_t[16] = 11'b00000110011;
        x_t[17] = 11'b00000110001;
        x_t[18] = 11'b00000100111;
        x_t[19] = 11'b00000011110;
        x_t[20] = 11'b00000001100;
        x_t[21] = 11'b00000010011;
        x_t[22] = 11'b00000010000;
        x_t[23] = 11'b00000000110;
        x_t[24] = 11'b00000001100;
        x_t[25] = 11'b00000001011;
        x_t[26] = 11'b00000001111;
        x_t[27] = 11'b00000001111;
        x_t[28] = 11'b00000001111;
        x_t[29] = 11'b00000011001;
        x_t[30] = 11'b00000000101;
        x_t[31] = 11'b00000010001;
        x_t[32] = 11'b00000011100;
        x_t[33] = 11'b00000011010;
        x_t[34] = 11'b00000010101;
        x_t[35] = 11'b00000010111;
        x_t[36] = 11'b00000010001;
        x_t[37] = 11'b00000000001;
        x_t[38] = 11'b00000011101;
        x_t[39] = 11'b00000100001;
        x_t[40] = 11'b00000101110;
        x_t[41] = 11'b00000000011;
        x_t[42] = 11'b00000010010;
        x_t[43] = 11'b11111111001;
        x_t[44] = 11'b00000011111;
        x_t[45] = 11'b00000011001;
        x_t[46] = 11'b00000011100;
        x_t[47] = 11'b00000100011;
        x_t[48] = 11'b00000011101;
        x_t[49] = 11'b00000101010;
        x_t[50] = 11'b00000101100;
        x_t[51] = 11'b00000100000;
        x_t[52] = 11'b00000011011;
        x_t[53] = 11'b00000001110;
        x_t[54] = 11'b00000000011;
        x_t[55] = 11'b00000001110;
        x_t[56] = 11'b00000010101;
        x_t[57] = 11'b00000011001;
        x_t[58] = 11'b00000001010;
        x_t[59] = 11'b11111111101;
        x_t[60] = 11'b11111110111;
        x_t[61] = 11'b11111101011;
        x_t[62] = 11'b11111001110;
        x_t[63] = 11'b11111001111;
        
        h_t_prev[0] = 11'b00000011010;
        h_t_prev[1] = 11'b00000100110;
        h_t_prev[2] = 11'b00000100111;
        h_t_prev[3] = 11'b00000101011;
        h_t_prev[4] = 11'b00000100111;
        h_t_prev[5] = 11'b00000011011;
        h_t_prev[6] = 11'b00000010010;
        h_t_prev[7] = 11'b00000010110;
        h_t_prev[8] = 11'b00000100111;
        h_t_prev[9] = 11'b00000110101;
        h_t_prev[10] = 11'b00001000010;
        h_t_prev[11] = 11'b00000100110;
        h_t_prev[12] = 11'b00000011101;
        h_t_prev[13] = 11'b00000011100;
        h_t_prev[14] = 11'b00000100000;
        h_t_prev[15] = 11'b00000101101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 93 timeout!");
                $fdisplay(fd_cycles, "Test Vector  93: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  93: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 93");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 94
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000100100;
        x_t[1] = 11'b00000101111;
        x_t[2] = 11'b00000101111;
        x_t[3] = 11'b00000110001;
        x_t[4] = 11'b00000101110;
        x_t[5] = 11'b00000100010;
        x_t[6] = 11'b00000011000;
        x_t[7] = 11'b00000100001;
        x_t[8] = 11'b00000110000;
        x_t[9] = 11'b00000111001;
        x_t[10] = 11'b00001000001;
        x_t[11] = 11'b00000101110;
        x_t[12] = 11'b00000101000;
        x_t[13] = 11'b00000100111;
        x_t[14] = 11'b00000101000;
        x_t[15] = 11'b00000110001;
        x_t[16] = 11'b00000110101;
        x_t[17] = 11'b00000110000;
        x_t[18] = 11'b00000101101;
        x_t[19] = 11'b00000101011;
        x_t[20] = 11'b00000011010;
        x_t[21] = 11'b00000001101;
        x_t[22] = 11'b00000001010;
        x_t[23] = 11'b11111111101;
        x_t[24] = 11'b00000000010;
        x_t[25] = 11'b00000000010;
        x_t[26] = 11'b00000000111;
        x_t[27] = 11'b00000000100;
        x_t[28] = 11'b11111111110;
        x_t[29] = 11'b00000001100;
        x_t[30] = 11'b00000000000;
        x_t[31] = 11'b00000000111;
        x_t[32] = 11'b00000010010;
        x_t[33] = 11'b00000001111;
        x_t[34] = 11'b00000001000;
        x_t[35] = 11'b00000001001;
        x_t[36] = 11'b11111111101;
        x_t[37] = 11'b11111110100;
        x_t[38] = 11'b00000010010;
        x_t[39] = 11'b00000010101;
        x_t[40] = 11'b00000011101;
        x_t[41] = 11'b11111111000;
        x_t[42] = 11'b00000000001;
        x_t[43] = 11'b11111011111;
        x_t[44] = 11'b00000001110;
        x_t[45] = 11'b00000010010;
        x_t[46] = 11'b00000010110;
        x_t[47] = 11'b00000011100;
        x_t[48] = 11'b00000010100;
        x_t[49] = 11'b00000100000;
        x_t[50] = 11'b00000011111;
        x_t[51] = 11'b00000011110;
        x_t[52] = 11'b00000011010;
        x_t[53] = 11'b00000010001;
        x_t[54] = 11'b00000000100;
        x_t[55] = 11'b00000001100;
        x_t[56] = 11'b00000001111;
        x_t[57] = 11'b00000011000;
        x_t[58] = 11'b00000010010;
        x_t[59] = 11'b00000001010;
        x_t[60] = 11'b00000001010;
        x_t[61] = 11'b00000000101;
        x_t[62] = 11'b11111110010;
        x_t[63] = 11'b11111100011;
        
        h_t_prev[0] = 11'b00000100100;
        h_t_prev[1] = 11'b00000101111;
        h_t_prev[2] = 11'b00000101111;
        h_t_prev[3] = 11'b00000110001;
        h_t_prev[4] = 11'b00000101110;
        h_t_prev[5] = 11'b00000100010;
        h_t_prev[6] = 11'b00000011000;
        h_t_prev[7] = 11'b00000100001;
        h_t_prev[8] = 11'b00000110000;
        h_t_prev[9] = 11'b00000111001;
        h_t_prev[10] = 11'b00001000001;
        h_t_prev[11] = 11'b00000101110;
        h_t_prev[12] = 11'b00000101000;
        h_t_prev[13] = 11'b00000100111;
        h_t_prev[14] = 11'b00000101000;
        h_t_prev[15] = 11'b00000110001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 94 timeout!");
                $fdisplay(fd_cycles, "Test Vector  94: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  94: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 94");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 95
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000010010;
        x_t[1] = 11'b00000011010;
        x_t[2] = 11'b00000010110;
        x_t[3] = 11'b00000010101;
        x_t[4] = 11'b00000010001;
        x_t[5] = 11'b00000000011;
        x_t[6] = 11'b11111110100;
        x_t[7] = 11'b00000001111;
        x_t[8] = 11'b00000011101;
        x_t[9] = 11'b00000100000;
        x_t[10] = 11'b00000100111;
        x_t[11] = 11'b00000010110;
        x_t[12] = 11'b00000010100;
        x_t[13] = 11'b00000001101;
        x_t[14] = 11'b00000011000;
        x_t[15] = 11'b00000100001;
        x_t[16] = 11'b00000100011;
        x_t[17] = 11'b00000011110;
        x_t[18] = 11'b00000011111;
        x_t[19] = 11'b00000011111;
        x_t[20] = 11'b00000010001;
        x_t[21] = 11'b11111111011;
        x_t[22] = 11'b11111111010;
        x_t[23] = 11'b11111110001;
        x_t[24] = 11'b11111110010;
        x_t[25] = 11'b11111110010;
        x_t[26] = 11'b11111110010;
        x_t[27] = 11'b11111110001;
        x_t[28] = 11'b11111111100;
        x_t[29] = 11'b11111111100;
        x_t[30] = 11'b11111110010;
        x_t[31] = 11'b11111101111;
        x_t[32] = 11'b11111111111;
        x_t[33] = 11'b11111110111;
        x_t[34] = 11'b11111101111;
        x_t[35] = 11'b11111110011;
        x_t[36] = 11'b11111100111;
        x_t[37] = 11'b11111101010;
        x_t[38] = 11'b00000000000;
        x_t[39] = 11'b00000000000;
        x_t[40] = 11'b00000000111;
        x_t[41] = 11'b11111010111;
        x_t[42] = 11'b00000000001;
        x_t[43] = 11'b00000010110;
        x_t[44] = 11'b00000000111;
        x_t[45] = 11'b00000011010;
        x_t[46] = 11'b00000011011;
        x_t[47] = 11'b00000011100;
        x_t[48] = 11'b00000011000;
        x_t[49] = 11'b00000100101;
        x_t[50] = 11'b00000100011;
        x_t[51] = 11'b00000101000;
        x_t[52] = 11'b00000100101;
        x_t[53] = 11'b00000100000;
        x_t[54] = 11'b00000011001;
        x_t[55] = 11'b00000011001;
        x_t[56] = 11'b00000011101;
        x_t[57] = 11'b00000101000;
        x_t[58] = 11'b00000100111;
        x_t[59] = 11'b00000100101;
        x_t[60] = 11'b00000011011;
        x_t[61] = 11'b00000011110;
        x_t[62] = 11'b00000001101;
        x_t[63] = 11'b11111111110;
        
        h_t_prev[0] = 11'b00000010010;
        h_t_prev[1] = 11'b00000011010;
        h_t_prev[2] = 11'b00000010110;
        h_t_prev[3] = 11'b00000010101;
        h_t_prev[4] = 11'b00000010001;
        h_t_prev[5] = 11'b00000000011;
        h_t_prev[6] = 11'b11111110100;
        h_t_prev[7] = 11'b00000001111;
        h_t_prev[8] = 11'b00000011101;
        h_t_prev[9] = 11'b00000100000;
        h_t_prev[10] = 11'b00000100111;
        h_t_prev[11] = 11'b00000010110;
        h_t_prev[12] = 11'b00000010100;
        h_t_prev[13] = 11'b00000001101;
        h_t_prev[14] = 11'b00000011000;
        h_t_prev[15] = 11'b00000100001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 95 timeout!");
                $fdisplay(fd_cycles, "Test Vector  95: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  95: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 95");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 96
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000001001;
        x_t[1] = 11'b00000010000;
        x_t[2] = 11'b00000001011;
        x_t[3] = 11'b00000001011;
        x_t[4] = 11'b00000000110;
        x_t[5] = 11'b11111111001;
        x_t[6] = 11'b11111101110;
        x_t[7] = 11'b00000001001;
        x_t[8] = 11'b00000010100;
        x_t[9] = 11'b00000011010;
        x_t[10] = 11'b00000100100;
        x_t[11] = 11'b00000010011;
        x_t[12] = 11'b00000010010;
        x_t[13] = 11'b00000001010;
        x_t[14] = 11'b00000010101;
        x_t[15] = 11'b00000011110;
        x_t[16] = 11'b00000100000;
        x_t[17] = 11'b00000100001;
        x_t[18] = 11'b00000100011;
        x_t[19] = 11'b00000100100;
        x_t[20] = 11'b00000010111;
        x_t[21] = 11'b11111110111;
        x_t[22] = 11'b11111110100;
        x_t[23] = 11'b11111101100;
        x_t[24] = 11'b11111101111;
        x_t[25] = 11'b11111110000;
        x_t[26] = 11'b11111101011;
        x_t[27] = 11'b11111101100;
        x_t[28] = 11'b11111111011;
        x_t[29] = 11'b11111111101;
        x_t[30] = 11'b11111110001;
        x_t[31] = 11'b11111101110;
        x_t[32] = 11'b11111111010;
        x_t[33] = 11'b11111110100;
        x_t[34] = 11'b11111101011;
        x_t[35] = 11'b11111101101;
        x_t[36] = 11'b11111100110;
        x_t[37] = 11'b11111100111;
        x_t[38] = 11'b11111111111;
        x_t[39] = 11'b11111110111;
        x_t[40] = 11'b00000001000;
        x_t[41] = 11'b11111001111;
        x_t[42] = 11'b00000001000;
        x_t[43] = 11'b00000011110;
        x_t[44] = 11'b11111111101;
        x_t[45] = 11'b00000101001;
        x_t[46] = 11'b00000010010;
        x_t[47] = 11'b00000011001;
        x_t[48] = 11'b00000010110;
        x_t[49] = 11'b00000100110;
        x_t[50] = 11'b00000101000;
        x_t[51] = 11'b00000101101;
        x_t[52] = 11'b00000101001;
        x_t[53] = 11'b00000100111;
        x_t[54] = 11'b00000100110;
        x_t[55] = 11'b00000011101;
        x_t[56] = 11'b00000011110;
        x_t[57] = 11'b00000110000;
        x_t[58] = 11'b00000101110;
        x_t[59] = 11'b00000110000;
        x_t[60] = 11'b00000101001;
        x_t[61] = 11'b00000110011;
        x_t[62] = 11'b00000011111;
        x_t[63] = 11'b00000011001;
        
        h_t_prev[0] = 11'b00000001001;
        h_t_prev[1] = 11'b00000010000;
        h_t_prev[2] = 11'b00000001011;
        h_t_prev[3] = 11'b00000001011;
        h_t_prev[4] = 11'b00000000110;
        h_t_prev[5] = 11'b11111111001;
        h_t_prev[6] = 11'b11111101110;
        h_t_prev[7] = 11'b00000001001;
        h_t_prev[8] = 11'b00000010100;
        h_t_prev[9] = 11'b00000011010;
        h_t_prev[10] = 11'b00000100100;
        h_t_prev[11] = 11'b00000010011;
        h_t_prev[12] = 11'b00000010010;
        h_t_prev[13] = 11'b00000001010;
        h_t_prev[14] = 11'b00000010101;
        h_t_prev[15] = 11'b00000011110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 96 timeout!");
                $fdisplay(fd_cycles, "Test Vector  96: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  96: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 96");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 97
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111111001;
        x_t[1] = 11'b11111111001;
        x_t[2] = 11'b11111101111;
        x_t[3] = 11'b11111110101;
        x_t[4] = 11'b11111111000;
        x_t[5] = 11'b11111110100;
        x_t[6] = 11'b11111111001;
        x_t[7] = 11'b11111111111;
        x_t[8] = 11'b11111110010;
        x_t[9] = 11'b11111101011;
        x_t[10] = 11'b11111101110;
        x_t[11] = 11'b11111101101;
        x_t[12] = 11'b11111111000;
        x_t[13] = 11'b00000000101;
        x_t[14] = 11'b11111110010;
        x_t[15] = 11'b11111110011;
        x_t[16] = 11'b11111101110;
        x_t[17] = 11'b11111101100;
        x_t[18] = 11'b11111110101;
        x_t[19] = 11'b11111110001;
        x_t[20] = 11'b00000000110;
        x_t[21] = 11'b00000001100;
        x_t[22] = 11'b00000001100;
        x_t[23] = 11'b00000000111;
        x_t[24] = 11'b00000000111;
        x_t[25] = 11'b00000000111;
        x_t[26] = 11'b00000000011;
        x_t[27] = 11'b11111111011;
        x_t[28] = 11'b11111110111;
        x_t[29] = 11'b00000000010;
        x_t[30] = 11'b00000001000;
        x_t[31] = 11'b11111111101;
        x_t[32] = 11'b00000000010;
        x_t[33] = 11'b11111111010;
        x_t[34] = 11'b11111111010;
        x_t[35] = 11'b11111111100;
        x_t[36] = 11'b11111111000;
        x_t[37] = 11'b11111111001;
        x_t[38] = 11'b00000000000;
        x_t[39] = 11'b00000010010;
        x_t[40] = 11'b11111111110;
        x_t[41] = 11'b00000110001;
        x_t[42] = 11'b11111111010;
        x_t[43] = 11'b00000010000;
        x_t[44] = 11'b11111110000;
        x_t[45] = 11'b00000010101;
        x_t[46] = 11'b11111101000;
        x_t[47] = 11'b11111110011;
        x_t[48] = 11'b11111110011;
        x_t[49] = 11'b11111110101;
        x_t[50] = 11'b11111110011;
        x_t[51] = 11'b11111110111;
        x_t[52] = 11'b11111110111;
        x_t[53] = 11'b11111111110;
        x_t[54] = 11'b00000000110;
        x_t[55] = 11'b11111101010;
        x_t[56] = 11'b11111110101;
        x_t[57] = 11'b11111111000;
        x_t[58] = 11'b11111111010;
        x_t[59] = 11'b11111111001;
        x_t[60] = 11'b11111111001;
        x_t[61] = 11'b11111110100;
        x_t[62] = 11'b11111110101;
        x_t[63] = 11'b00000000010;
        
        h_t_prev[0] = 11'b11111111001;
        h_t_prev[1] = 11'b11111111001;
        h_t_prev[2] = 11'b11111101111;
        h_t_prev[3] = 11'b11111110101;
        h_t_prev[4] = 11'b11111111000;
        h_t_prev[5] = 11'b11111110100;
        h_t_prev[6] = 11'b11111111001;
        h_t_prev[7] = 11'b11111111111;
        h_t_prev[8] = 11'b11111110010;
        h_t_prev[9] = 11'b11111101011;
        h_t_prev[10] = 11'b11111101110;
        h_t_prev[11] = 11'b11111101101;
        h_t_prev[12] = 11'b11111111000;
        h_t_prev[13] = 11'b00000000101;
        h_t_prev[14] = 11'b11111110010;
        h_t_prev[15] = 11'b11111110011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 97 timeout!");
                $fdisplay(fd_cycles, "Test Vector  97: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  97: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 97");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 98
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b00000000001;
        x_t[1] = 11'b00000000000;
        x_t[2] = 11'b11111110101;
        x_t[3] = 11'b11111111101;
        x_t[4] = 11'b11111111100;
        x_t[5] = 11'b11111110111;
        x_t[6] = 11'b11111111010;
        x_t[7] = 11'b00000000011;
        x_t[8] = 11'b11111110100;
        x_t[9] = 11'b11111101110;
        x_t[10] = 11'b11111110011;
        x_t[11] = 11'b11111110011;
        x_t[12] = 11'b11111111010;
        x_t[13] = 11'b00000001011;
        x_t[14] = 11'b11111110011;
        x_t[15] = 11'b11111110000;
        x_t[16] = 11'b11111101110;
        x_t[17] = 11'b11111101110;
        x_t[18] = 11'b11111110101;
        x_t[19] = 11'b11111101111;
        x_t[20] = 11'b00000000011;
        x_t[21] = 11'b00000001101;
        x_t[22] = 11'b00000001011;
        x_t[23] = 11'b00000000110;
        x_t[24] = 11'b00000001000;
        x_t[25] = 11'b00000000111;
        x_t[26] = 11'b00000000010;
        x_t[27] = 11'b11111111100;
        x_t[28] = 11'b11111110101;
        x_t[29] = 11'b00000000010;
        x_t[30] = 11'b00000001000;
        x_t[31] = 11'b11111111110;
        x_t[32] = 11'b00000000010;
        x_t[33] = 11'b11111111001;
        x_t[34] = 11'b11111111001;
        x_t[35] = 11'b11111111001;
        x_t[36] = 11'b11111110111;
        x_t[37] = 11'b11111110100;
        x_t[38] = 11'b11111111111;
        x_t[39] = 11'b00000001001;
        x_t[40] = 11'b11111110111;
        x_t[41] = 11'b00000000101;
        x_t[42] = 11'b11111110011;
        x_t[43] = 11'b00000001001;
        x_t[44] = 11'b11111101000;
        x_t[45] = 11'b00000001010;
        x_t[46] = 11'b11111100001;
        x_t[47] = 11'b11111101010;
        x_t[48] = 11'b11111101011;
        x_t[49] = 11'b11111101110;
        x_t[50] = 11'b11111101101;
        x_t[51] = 11'b11111110000;
        x_t[52] = 11'b11111110000;
        x_t[53] = 11'b11111110100;
        x_t[54] = 11'b11111110111;
        x_t[55] = 11'b11111011111;
        x_t[56] = 11'b11111101010;
        x_t[57] = 11'b11111101111;
        x_t[58] = 11'b11111110011;
        x_t[59] = 11'b11111110100;
        x_t[60] = 11'b11111110010;
        x_t[61] = 11'b11111110000;
        x_t[62] = 11'b11111110100;
        x_t[63] = 11'b11111111101;
        
        h_t_prev[0] = 11'b00000000001;
        h_t_prev[1] = 11'b00000000000;
        h_t_prev[2] = 11'b11111110101;
        h_t_prev[3] = 11'b11111111101;
        h_t_prev[4] = 11'b11111111100;
        h_t_prev[5] = 11'b11111110111;
        h_t_prev[6] = 11'b11111111010;
        h_t_prev[7] = 11'b00000000011;
        h_t_prev[8] = 11'b11111110100;
        h_t_prev[9] = 11'b11111101110;
        h_t_prev[10] = 11'b11111110011;
        h_t_prev[11] = 11'b11111110011;
        h_t_prev[12] = 11'b11111111010;
        h_t_prev[13] = 11'b00000001011;
        h_t_prev[14] = 11'b11111110011;
        h_t_prev[15] = 11'b11111110000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 98 timeout!");
                $fdisplay(fd_cycles, "Test Vector  98: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  98: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 98");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 99
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111110111;
        x_t[1] = 11'b11111110101;
        x_t[2] = 11'b11111101100;
        x_t[3] = 11'b11111110100;
        x_t[4] = 11'b11111110011;
        x_t[5] = 11'b11111101110;
        x_t[6] = 11'b11111101110;
        x_t[7] = 11'b11111110101;
        x_t[8] = 11'b11111100101;
        x_t[9] = 11'b11111100000;
        x_t[10] = 11'b11111100110;
        x_t[11] = 11'b11111100100;
        x_t[12] = 11'b11111101000;
        x_t[13] = 11'b11111110010;
        x_t[14] = 11'b11111100110;
        x_t[15] = 11'b11111011111;
        x_t[16] = 11'b11111011100;
        x_t[17] = 11'b11111011111;
        x_t[18] = 11'b11111100011;
        x_t[19] = 11'b11111011010;
        x_t[20] = 11'b11111100110;
        x_t[21] = 11'b00000001001;
        x_t[22] = 11'b00000000111;
        x_t[23] = 11'b00000000011;
        x_t[24] = 11'b00000000001;
        x_t[25] = 11'b00000000001;
        x_t[26] = 11'b11111111010;
        x_t[27] = 11'b11111110101;
        x_t[28] = 11'b11111110000;
        x_t[29] = 11'b11111111011;
        x_t[30] = 11'b00000000001;
        x_t[31] = 11'b11111110101;
        x_t[32] = 11'b11111110111;
        x_t[33] = 11'b11111101111;
        x_t[34] = 11'b11111110000;
        x_t[35] = 11'b11111110001;
        x_t[36] = 11'b11111101100;
        x_t[37] = 11'b11111101100;
        x_t[38] = 11'b11111111000;
        x_t[39] = 11'b11111110010;
        x_t[40] = 11'b11111110001;
        x_t[41] = 11'b11111100011;
        x_t[42] = 11'b11111101110;
        x_t[43] = 11'b11111110110;
        x_t[44] = 11'b11111100010;
        x_t[45] = 11'b11111100001;
        x_t[46] = 11'b11111011001;
        x_t[47] = 11'b11111011100;
        x_t[48] = 11'b11111011010;
        x_t[49] = 11'b11111011001;
        x_t[50] = 11'b11111011001;
        x_t[51] = 11'b11111011000;
        x_t[52] = 11'b11111010101;
        x_t[53] = 11'b11111010011;
        x_t[54] = 11'b11111001110;
        x_t[55] = 11'b11111010011;
        x_t[56] = 11'b11111011010;
        x_t[57] = 11'b11111011100;
        x_t[58] = 11'b11111011100;
        x_t[59] = 11'b11111011001;
        x_t[60] = 11'b11111100111;
        x_t[61] = 11'b11111100011;
        x_t[62] = 11'b11111101001;
        x_t[63] = 11'b11111110000;
        
        h_t_prev[0] = 11'b11111110111;
        h_t_prev[1] = 11'b11111110101;
        h_t_prev[2] = 11'b11111101100;
        h_t_prev[3] = 11'b11111110100;
        h_t_prev[4] = 11'b11111110011;
        h_t_prev[5] = 11'b11111101110;
        h_t_prev[6] = 11'b11111101110;
        h_t_prev[7] = 11'b11111110101;
        h_t_prev[8] = 11'b11111100101;
        h_t_prev[9] = 11'b11111100000;
        h_t_prev[10] = 11'b11111100110;
        h_t_prev[11] = 11'b11111100100;
        h_t_prev[12] = 11'b11111101000;
        h_t_prev[13] = 11'b11111110010;
        h_t_prev[14] = 11'b11111100110;
        h_t_prev[15] = 11'b11111011111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 99 timeout!");
                $fdisplay(fd_cycles, "Test Vector  99: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  99: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 99");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 100
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 11'b11111110111;
        x_t[1] = 11'b11111110010;
        x_t[2] = 11'b11111100101;
        x_t[3] = 11'b11111101111;
        x_t[4] = 11'b11111101111;
        x_t[5] = 11'b11111101001;
        x_t[6] = 11'b11111101100;
        x_t[7] = 11'b11111111001;
        x_t[8] = 11'b11111011111;
        x_t[9] = 11'b11111011000;
        x_t[10] = 11'b11111011011;
        x_t[11] = 11'b11111011000;
        x_t[12] = 11'b11111011001;
        x_t[13] = 11'b11111100010;
        x_t[14] = 11'b11111100111;
        x_t[15] = 11'b11111011011;
        x_t[16] = 11'b11111010010;
        x_t[17] = 11'b11111010011;
        x_t[18] = 11'b11111011000;
        x_t[19] = 11'b11111001001;
        x_t[20] = 11'b11111010010;
        x_t[21] = 11'b00000010001;
        x_t[22] = 11'b00000010010;
        x_t[23] = 11'b00000001101;
        x_t[24] = 11'b00000001011;
        x_t[25] = 11'b00000001010;
        x_t[26] = 11'b00000000110;
        x_t[27] = 11'b00000000001;
        x_t[28] = 11'b11111111001;
        x_t[29] = 11'b00000001001;
        x_t[30] = 11'b00000001001;
        x_t[31] = 11'b11111111110;
        x_t[32] = 11'b11111111110;
        x_t[33] = 11'b11111111011;
        x_t[34] = 11'b11111111101;
        x_t[35] = 11'b11111111101;
        x_t[36] = 11'b11111111011;
        x_t[37] = 11'b11111111010;
        x_t[38] = 11'b00000000110;
        x_t[39] = 11'b11111111101;
        x_t[40] = 11'b00000000011;
        x_t[41] = 11'b11111111000;
        x_t[42] = 11'b00000000100;
        x_t[43] = 11'b11111011011;
        x_t[44] = 11'b11111101001;
        x_t[45] = 11'b11111000100;
        x_t[46] = 11'b11111011101;
        x_t[47] = 11'b11111011100;
        x_t[48] = 11'b11111010111;
        x_t[49] = 11'b11111010010;
        x_t[50] = 11'b11111010000;
        x_t[51] = 11'b11111001111;
        x_t[52] = 11'b11111001110;
        x_t[53] = 11'b11111001000;
        x_t[54] = 11'b11111000010;
        x_t[55] = 11'b11111001111;
        x_t[56] = 11'b11111010010;
        x_t[57] = 11'b11111010100;
        x_t[58] = 11'b11111010011;
        x_t[59] = 11'b11111010000;
        x_t[60] = 11'b11111011110;
        x_t[61] = 11'b11111011000;
        x_t[62] = 11'b11111011110;
        x_t[63] = 11'b11111101011;
        
        h_t_prev[0] = 11'b11111110111;
        h_t_prev[1] = 11'b11111110010;
        h_t_prev[2] = 11'b11111100101;
        h_t_prev[3] = 11'b11111101111;
        h_t_prev[4] = 11'b11111101111;
        h_t_prev[5] = 11'b11111101001;
        h_t_prev[6] = 11'b11111101100;
        h_t_prev[7] = 11'b11111111001;
        h_t_prev[8] = 11'b11111011111;
        h_t_prev[9] = 11'b11111011000;
        h_t_prev[10] = 11'b11111011011;
        h_t_prev[11] = 11'b11111011000;
        h_t_prev[12] = 11'b11111011001;
        h_t_prev[13] = 11'b11111100010;
        h_t_prev[14] = 11'b11111100111;
        h_t_prev[15] = 11'b11111011011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 100 timeout!");
                $fdisplay(fd_cycles, "Test Vector 100: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector 100: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b %011b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 100");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Write summary to cycles file
    $fdisplay(fd_cycles, "");
    $fdisplay(fd_cycles, "==========================================================");
    $fdisplay(fd_cycles, "SUMMARY");
    $fdisplay(fd_cycles, "==========================================================");
    $fdisplay(fd_cycles, "Total Test Vectors: %0d", 100);
    $fdisplay(fd_cycles, "Total Cycles:       %0d", total_cycles);
    $fdisplay(fd_cycles, "Average Cycles:     %.2f", real'(total_cycles) / 100);
    $fdisplay(fd_cycles, "Total Time:         %.2f us @ 100MHz", total_cycles * 0.01);
    $fdisplay(fd_cycles, "Average Time:       %.2f us @ 100MHz", (total_cycles * 0.01) / 100);
    $fdisplay(fd_cycles, "Throughput:         %.2f computations/ms @ 100MHz", 100000.0 / (real'(total_cycles) / 100));
    $fdisplay(fd_cycles, "==========================================================");
    
    $fclose(fd_output);
    $fclose(fd_cycles);
    
    $display("");
    $display("==========================================================");
    $display("Simulation Complete");
    $display("==========================================================");
    $display("Test Vectors:   %0d", 100);
    $display("Total Cycles:   %0d", total_cycles);
    $display("Average Cycles: %.2f", real'(total_cycles) / 100);
    $display("==========================================================");
    $display("Output file:    output_d64_h16_dw11_fb5_np1.txt");
    $display("Cycles file:    cycles_d64_h16_dw11_fb5_np1.txt");
    $display("==========================================================");
    
    $finish;
end

endmodule