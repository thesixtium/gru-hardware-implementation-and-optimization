`timescale 1ns / 1ps

module gru_tb;

// Parameters
parameter int INT_WIDTH  = 5;
parameter int FRAC_WIDTH = 5;
parameter int WIDTH      = INT_WIDTH + FRAC_WIDTH + 1;
parameter real CLK_PERIOD = 10.0;

// Clock and reset
logic clk;
logic reset;

// Inputs
logic signed [WIDTH-1:0] x_0 = 0;
logic signed [WIDTH-1:0] x_1 = 0;
logic signed [WIDTH-1:0] x_2 = 0;
logic signed [WIDTH-1:0] x_3 = 0;
logic signed [WIDTH-1:0] x_4 = 0;

logic signed [WIDTH-1:0] h_0 = 0;
logic signed [WIDTH-1:0] h_1 = 0;
logic signed [WIDTH-1:0] h_2 = 0;
logic signed [WIDTH-1:0] h_3 = 0;

// Input weights (h×d for each gate)
logic signed [WIDTH-1:0] w_ir_0_0 = 'b0000000011;
logic signed [WIDTH-1:0] w_ir_0_1 = 'b0000000101;
logic signed [WIDTH-1:0] w_ir_0_2 = 'b0000000100;
logic signed [WIDTH-1:0] w_ir_0_3 = 'b0000000100;
logic signed [WIDTH-1:0] w_ir_0_4 = 'b1111111110;
logic signed [WIDTH-1:0] w_ir_1_0 = 'b1111111011;
logic signed [WIDTH-1:0] w_ir_1_1 = 'b0000000100;
logic signed [WIDTH-1:0] w_ir_1_2 = 'b0000000010;
logic signed [WIDTH-1:0] w_ir_1_3 = 'b1111111001;
logic signed [WIDTH-1:0] w_ir_1_4 = 'b0000000001;
logic signed [WIDTH-1:0] w_ir_2_0 = 'b0000001000;
logic signed [WIDTH-1:0] w_ir_2_1 = 'b0000000000;
logic signed [WIDTH-1:0] w_ir_2_2 = 'b0000000101;
logic signed [WIDTH-1:0] w_ir_2_3 = 'b0000000001;
logic signed [WIDTH-1:0] w_ir_2_4 = 'b0000000001;
logic signed [WIDTH-1:0] w_ir_3_0 = 'b0000000110;
logic signed [WIDTH-1:0] w_ir_3_1 = 'b1111111111;
logic signed [WIDTH-1:0] w_ir_3_2 = 'b0000000111;
logic signed [WIDTH-1:0] w_ir_3_3 = 'b1111111111;
logic signed [WIDTH-1:0] w_ir_3_4 = 'b0000000101;

logic signed [WIDTH-1:0] w_iz_0_0 = 'b1111111111;
logic signed [WIDTH-1:0] w_iz_0_1 = 'b0000000100;
logic signed [WIDTH-1:0] w_iz_0_2 = 'b0000000011;
logic signed [WIDTH-1:0] w_iz_0_3 = 'b0000000011;
logic signed [WIDTH-1:0] w_iz_0_4 = 'b1111111011;
logic signed [WIDTH-1:0] w_iz_1_0 = 'b0000000100;
logic signed [WIDTH-1:0] w_iz_1_1 = 'b0000000100;
logic signed [WIDTH-1:0] w_iz_1_2 = 'b0000000011;
logic signed [WIDTH-1:0] w_iz_1_3 = 'b0000000111;
logic signed [WIDTH-1:0] w_iz_1_4 = 'b1111111001;
logic signed [WIDTH-1:0] w_iz_2_0 = 'b1111111110;
logic signed [WIDTH-1:0] w_iz_2_1 = 'b0000000011;
logic signed [WIDTH-1:0] w_iz_2_2 = 'b0000000010;
logic signed [WIDTH-1:0] w_iz_2_3 = 'b0000000100;
logic signed [WIDTH-1:0] w_iz_2_4 = 'b0000000100;
logic signed [WIDTH-1:0] w_iz_3_0 = 'b0000000001;
logic signed [WIDTH-1:0] w_iz_3_1 = 'b0000001000;
logic signed [WIDTH-1:0] w_iz_3_2 = 'b0000000011;
logic signed [WIDTH-1:0] w_iz_3_3 = 'b1111111110;
logic signed [WIDTH-1:0] w_iz_3_4 = 'b0000000010;

logic signed [WIDTH-1:0] w_in_0_0 = 'b0000000101;
logic signed [WIDTH-1:0] w_in_0_1 = 'b1111111010;
logic signed [WIDTH-1:0] w_in_0_2 = 'b0000000010;
logic signed [WIDTH-1:0] w_in_0_3 = 'b1111111101;
logic signed [WIDTH-1:0] w_in_0_4 = 'b0000000000;
logic signed [WIDTH-1:0] w_in_1_0 = 'b1111111100;
logic signed [WIDTH-1:0] w_in_1_1 = 'b1111111010;
logic signed [WIDTH-1:0] w_in_1_2 = 'b0000000111;
logic signed [WIDTH-1:0] w_in_1_3 = 'b1111111110;
logic signed [WIDTH-1:0] w_in_1_4 = 'b1111111101;
logic signed [WIDTH-1:0] w_in_2_0 = 'b1111111111;
logic signed [WIDTH-1:0] w_in_2_1 = 'b0000000000;
logic signed [WIDTH-1:0] w_in_2_2 = 'b1111111001;
logic signed [WIDTH-1:0] w_in_2_3 = 'b1111111101;
logic signed [WIDTH-1:0] w_in_2_4 = 'b0000000010;
logic signed [WIDTH-1:0] w_in_3_0 = 'b1111111101;
logic signed [WIDTH-1:0] w_in_3_1 = 'b0000000101;
logic signed [WIDTH-1:0] w_in_3_2 = 'b1111111101;
logic signed [WIDTH-1:0] w_in_3_3 = 'b1111111101;
logic signed [WIDTH-1:0] w_in_3_4 = 'b0000000100;

// Recurrent weights (h×h for each gate)
logic signed [WIDTH-1:0] w_hr_0_0 = 'b0000000000;
logic signed [WIDTH-1:0] w_hr_0_1 = 'b0000000001;
logic signed [WIDTH-1:0] w_hr_0_2 = 'b0000000010;
logic signed [WIDTH-1:0] w_hr_0_3 = 'b1111111011;
logic signed [WIDTH-1:0] w_hr_1_0 = 'b0000001001;
logic signed [WIDTH-1:0] w_hr_1_1 = 'b0000001001;
logic signed [WIDTH-1:0] w_hr_1_2 = 'b0000001001;
logic signed [WIDTH-1:0] w_hr_1_3 = 'b1111110111;
logic signed [WIDTH-1:0] w_hr_2_0 = 'b0000001000;
logic signed [WIDTH-1:0] w_hr_2_1 = 'b0000001001;
logic signed [WIDTH-1:0] w_hr_2_2 = 'b1111111100;
logic signed [WIDTH-1:0] w_hr_2_3 = 'b1111111011;
logic signed [WIDTH-1:0] w_hr_3_0 = 'b0000000100;
logic signed [WIDTH-1:0] w_hr_3_1 = 'b0000000101;
logic signed [WIDTH-1:0] w_hr_3_2 = 'b0000001011;
logic signed [WIDTH-1:0] w_hr_3_3 = 'b1111111000;

logic signed [WIDTH-1:0] w_hz_0_0 = 'b0000000111;
logic signed [WIDTH-1:0] w_hz_0_1 = 'b0000000100;
logic signed [WIDTH-1:0] w_hz_0_2 = 'b1111111101;
logic signed [WIDTH-1:0] w_hz_0_3 = 'b0000000100;
logic signed [WIDTH-1:0] w_hz_1_0 = 'b0000001101;
logic signed [WIDTH-1:0] w_hz_1_1 = 'b1111110100;
logic signed [WIDTH-1:0] w_hz_1_2 = 'b0000000000;
logic signed [WIDTH-1:0] w_hz_1_3 = 'b0000001001;
logic signed [WIDTH-1:0] w_hz_2_0 = 'b0000000111;
logic signed [WIDTH-1:0] w_hz_2_1 = 'b0000000000;
logic signed [WIDTH-1:0] w_hz_2_2 = 'b1111110000;
logic signed [WIDTH-1:0] w_hz_2_3 = 'b0000001110;
logic signed [WIDTH-1:0] w_hz_3_0 = 'b0000001100;
logic signed [WIDTH-1:0] w_hz_3_1 = 'b0000000100;
logic signed [WIDTH-1:0] w_hz_3_2 = 'b1111110111;
logic signed [WIDTH-1:0] w_hz_3_3 = 'b0000010101;

logic signed [WIDTH-1:0] w_hn_0_0 = 'b1111111111;
logic signed [WIDTH-1:0] w_hn_0_1 = 'b1111111110;
logic signed [WIDTH-1:0] w_hn_0_2 = 'b0000000101;
logic signed [WIDTH-1:0] w_hn_0_3 = 'b1111111010;
logic signed [WIDTH-1:0] w_hn_1_0 = 'b1111111010;
logic signed [WIDTH-1:0] w_hn_1_1 = 'b1111111111;
logic signed [WIDTH-1:0] w_hn_1_2 = 'b0000010111;
logic signed [WIDTH-1:0] w_hn_1_3 = 'b1111110100;
logic signed [WIDTH-1:0] w_hn_2_0 = 'b1111111111;
logic signed [WIDTH-1:0] w_hn_2_1 = 'b0000001110;
logic signed [WIDTH-1:0] w_hn_2_2 = 'b0000010100;
logic signed [WIDTH-1:0] w_hn_2_3 = 'b1111110010;
logic signed [WIDTH-1:0] w_hn_3_0 = 'b1111111011;
logic signed [WIDTH-1:0] w_hn_3_1 = 'b1111110110;
logic signed [WIDTH-1:0] w_hn_3_2 = 'b1111111001;
logic signed [WIDTH-1:0] w_hn_3_3 = 'b0000001010;

// Biases (h for each gate type)
logic signed [WIDTH-1:0] b_ir_0 = 'b0000000001;
logic signed [WIDTH-1:0] b_ir_1 = 'b0000001000;
logic signed [WIDTH-1:0] b_ir_2 = 'b0000001111;
logic signed [WIDTH-1:0] b_ir_3 = 'b0000000101;

logic signed [WIDTH-1:0] b_iz_0 = 'b0000000110;
logic signed [WIDTH-1:0] b_iz_1 = 'b0000000100;
logic signed [WIDTH-1:0] b_iz_2 = 'b0000010000;
logic signed [WIDTH-1:0] b_iz_3 = 'b0000000000;

logic signed [WIDTH-1:0] b_in_0 = 'b0000001011;
logic signed [WIDTH-1:0] b_in_1 = 'b0000000010;
logic signed [WIDTH-1:0] b_in_2 = 'b0000001110;
logic signed [WIDTH-1:0] b_in_3 = 'b0000000010;

logic signed [WIDTH-1:0] b_hr_0 = 'b0000000010;
logic signed [WIDTH-1:0] b_hr_1 = 'b0000001010;
logic signed [WIDTH-1:0] b_hr_2 = 'b0000000111;
logic signed [WIDTH-1:0] b_hr_3 = 'b0000001101;

logic signed [WIDTH-1:0] b_hz_0 = 'b0000000111;
logic signed [WIDTH-1:0] b_hz_1 = 'b0000001001;
logic signed [WIDTH-1:0] b_hz_2 = 'b0000000101;
logic signed [WIDTH-1:0] b_hz_3 = 'b0000011010;

logic signed [WIDTH-1:0] b_hn_0 = 'b0000000011;
logic signed [WIDTH-1:0] b_hn_1 = 'b0000010011;
logic signed [WIDTH-1:0] b_hn_2 = 'b0000000111;
logic signed [WIDTH-1:0] b_hn_3 = 'b1111110001;

// Outputs (h=4)
logic signed [WIDTH-1:0]  y_0 = 0;
logic signed [WIDTH-1:0]  y_1 = 0;
logic signed [WIDTH-1:0]  y_2 = 0;
logic signed [WIDTH-1:0]  y_3 = 0;

gru #(
        .INT_WIDTH(INT_WIDTH),
        .FRAC_WIDTH(FRAC_WIDTH)
    ) gru_inst (
        .clk(clk),
        .reset(reset),
        // Input features (d=64)
        	
.x_0(x_0), .x_1(x_1), .x_2(x_2), .x_3(x_3), .x_4(x_4), 	
.h_0(h_0), .h_1(h_1), .h_2(h_2), .h_3(h_3), 	
.w_ir_0_0(w_ir_0_0), .w_ir_0_1(w_ir_0_1), .w_ir_0_2(w_ir_0_2), .w_ir_0_3(w_ir_0_3), .w_ir_0_4(w_ir_0_4), .w_ir_1_0(w_ir_1_0), .w_ir_1_1(w_ir_1_1), .w_ir_1_2(w_ir_1_2), .w_ir_1_3(w_ir_1_3), .w_ir_1_4(w_ir_1_4), .w_ir_2_0(w_ir_2_0), .w_ir_2_1(w_ir_2_1), .w_ir_2_2(w_ir_2_2), .w_ir_2_3(w_ir_2_3), .w_ir_2_4(w_ir_2_4), .w_ir_3_0(w_ir_3_0), .w_ir_3_1(w_ir_3_1), .w_ir_3_2(w_ir_3_2), .w_ir_3_3(w_ir_3_3), .w_ir_3_4(w_ir_3_4), 	
.w_iz_0_0(w_iz_0_0), .w_iz_0_1(w_iz_0_1), .w_iz_0_2(w_iz_0_2), .w_iz_0_3(w_iz_0_3), .w_iz_0_4(w_iz_0_4), .w_iz_1_0(w_iz_1_0), .w_iz_1_1(w_iz_1_1), .w_iz_1_2(w_iz_1_2), .w_iz_1_3(w_iz_1_3), .w_iz_1_4(w_iz_1_4), .w_iz_2_0(w_iz_2_0), .w_iz_2_1(w_iz_2_1), .w_iz_2_2(w_iz_2_2), .w_iz_2_3(w_iz_2_3), .w_iz_2_4(w_iz_2_4), .w_iz_3_0(w_iz_3_0), .w_iz_3_1(w_iz_3_1), .w_iz_3_2(w_iz_3_2), .w_iz_3_3(w_iz_3_3), .w_iz_3_4(w_iz_3_4), 
.w_in_0_0(w_in_0_0), .w_in_0_1(w_in_0_1), .w_in_0_2(w_in_0_2), .w_in_0_3(w_in_0_3), .w_in_0_4(w_in_0_4), .w_in_1_0(w_in_1_0), .w_in_1_1(w_in_1_1), .w_in_1_2(w_in_1_2), .w_in_1_3(w_in_1_3), .w_in_1_4(w_in_1_4), .w_in_2_0(w_in_2_0), .w_in_2_1(w_in_2_1), .w_in_2_2(w_in_2_2), .w_in_2_3(w_in_2_3), .w_in_2_4(w_in_2_4), .w_in_3_0(w_in_3_0), .w_in_3_1(w_in_3_1), .w_in_3_2(w_in_3_2), .w_in_3_3(w_in_3_3), .w_in_3_4(w_in_3_4), 
.w_hr_0_0(w_hr_0_0), .w_hr_0_1(w_hr_0_1), .w_hr_0_2(w_hr_0_2), .w_hr_0_3(w_hr_0_3), .w_hr_1_0(w_hr_1_0), .w_hr_1_1(w_hr_1_1), .w_hr_1_2(w_hr_1_2), .w_hr_1_3(w_hr_1_3), .w_hr_2_0(w_hr_2_0), .w_hr_2_1(w_hr_2_1), .w_hr_2_2(w_hr_2_2), .w_hr_2_3(w_hr_2_3), .w_hr_3_0(w_hr_3_0), .w_hr_3_1(w_hr_3_1), .w_hr_3_2(w_hr_3_2), .w_hr_3_3(w_hr_3_3), 
.w_hz_0_0(w_hz_0_0), .w_hz_0_1(w_hz_0_1), .w_hz_0_2(w_hz_0_2), .w_hz_0_3(w_hz_0_3), .w_hz_1_0(w_hz_1_0), .w_hz_1_1(w_hz_1_1), .w_hz_1_2(w_hz_1_2), .w_hz_1_3(w_hz_1_3), .w_hz_2_0(w_hz_2_0), .w_hz_2_1(w_hz_2_1), .w_hz_2_2(w_hz_2_2), .w_hz_2_3(w_hz_2_3), .w_hz_3_0(w_hz_3_0), .w_hz_3_1(w_hz_3_1), .w_hz_3_2(w_hz_3_2), .w_hz_3_3(w_hz_3_3), 
.w_hn_0_0(w_hn_0_0), .w_hn_0_1(w_hn_0_1), .w_hn_0_2(w_hn_0_2), .w_hn_0_3(w_hn_0_3), .w_hn_1_0(w_hn_1_0), .w_hn_1_1(w_hn_1_1), .w_hn_1_2(w_hn_1_2), .w_hn_1_3(w_hn_1_3), .w_hn_2_0(w_hn_2_0), .w_hn_2_1(w_hn_2_1), .w_hn_2_2(w_hn_2_2), .w_hn_2_3(w_hn_2_3), .w_hn_3_0(w_hn_3_0), .w_hn_3_1(w_hn_3_1), .w_hn_3_2(w_hn_3_2), .w_hn_3_3(w_hn_3_3), 
.b_ir_0(b_ir_0), .b_ir_1(b_ir_1), .b_ir_2(b_ir_2), .b_ir_3(b_ir_3), 
.b_iz_0(b_iz_0), .b_iz_1(b_iz_1), .b_iz_2(b_iz_2), .b_iz_3(b_iz_3), 
.b_in_0(b_in_0), .b_in_1(b_in_1), .b_in_2(b_in_2), .b_in_3(b_in_3), 
.b_hr_0(b_hr_0), .b_hr_1(b_hr_1), .b_hr_2(b_hr_2), .b_hr_3(b_hr_3), 
.b_hz_0(b_hz_0), .b_hz_1(b_hz_1), .b_hz_2(b_hz_2), .b_hz_3(b_hz_3), 
.b_hn_0(b_hn_0), .b_hn_1(b_hn_1), .b_hn_2(b_hn_2), .b_hn_3(b_hn_3), 
.y_0(y_0), .y_1(y_1), .y_2(y_2), .y_3(y_3)
);

    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end
    
    initial begin
        // Open file for writing (overwrite existing)
        integer fd;
        fd = $fopen("../../../../../output_d5_h4_int5_frac5.txt", "w+");
        if (fd == 0) begin
            $display("ERROR: Failed to open file!");
            $finish;
        end
        x_0 = 'b0000011101;
    x_1 = 'b1111101000;
    x_2 = 'b1111110111;
    x_3 = 'b0000100000;
    x_4 = 'b1111101111;

    h_0 = 'b0000001111;
    h_1 = 'b0000100000;
    h_2 = 'b0000010011;
    h_3 = 'b1111110101;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000000101;
    x_1 = 'b1111110111;
    x_2 = 'b0000001101;
    x_3 = 'b1111101111;
    x_4 = 'b0000010101;

    h_0 = 'b0000011011;
    h_1 = 'b0000000101;
    h_2 = 'b1111100001;
    h_3 = 'b0000010101;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111101000;
    x_1 = 'b0000100000;
    x_2 = 'b1111101111;
    x_3 = 'b1111110111;
    x_4 = 'b0000011101;

    h_0 = 'b0000100000;
    h_1 = 'b1111100001;
    h_2 = 'b0000011110;
    h_3 = 'b1111100100;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100001;
    x_1 = 'b1111101111;
    x_2 = 'b0000010101;
    x_3 = 'b0000011101;
    x_4 = 'b1111111100;

    h_0 = 'b0000011101;
    h_1 = 'b1111110111;
    h_2 = 'b1111101111;
    h_3 = 'b0000100000;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111110111;
    x_1 = 'b1111101111;
    x_2 = 'b1111101000;
    x_3 = 'b1111100011;
    x_4 = 'b1111100000;

    h_0 = 'b0000010011;
    h_1 = 'b0000011110;
    h_2 = 'b1111111110;
    h_3 = 'b1111100001;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000010101;
    x_1 = 'b0000100000;
    x_2 = 'b0000011011;
    x_3 = 'b0000001001;
    x_4 = 'b1111110010;

    h_0 = 'b0000000101;
    h_1 = 'b0000001101;
    h_2 = 'b0000010101;
    h_3 = 'b0000011011;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000100000;
    x_1 = 'b1111110111;
    x_2 = 'b1111100011;
    x_3 = 'b0000010010;
    x_4 = 'b0000011000;

    h_0 = 'b1111110101;
    h_1 = 'b1111100100;
    h_2 = 'b1111100001;
    h_3 = 'b1111101101;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000001101;
    x_1 = 'b1111101000;
    x_2 = 'b0000011111;
    x_3 = 'b1111100000;
    x_4 = 'b0000011011;

    h_0 = 'b1111101000;
    h_1 = 'b1111101111;
    h_2 = 'b0000011101;
    h_3 = 'b0000001001;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111101111;
    x_1 = 'b0000011101;
    x_2 = 'b1111100000;
    x_3 = 'b0000011000;
    x_4 = 'b1111111000;

    h_0 = 'b1111100001;
    h_1 = 'b0000011010;
    h_2 = 'b1111110000;
    h_3 = 'b0000000011;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100000;
    x_1 = 'b0000000000;
    x_2 = 'b0000100000;
    x_3 = 'b0000000001;
    x_4 = 'b1111100000;

    h_0 = 'b1111100001;
    h_1 = 'b0000010101;
    h_2 = 'b1111111100;
    h_3 = 'b1111110010;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111101111;
    x_1 = 'b1111100011;
    x_2 = 'b1111100000;
    x_3 = 'b1111100111;
    x_4 = 'b1111110110;

    h_0 = 'b1111101001;
    h_1 = 'b1111101001;
    h_2 = 'b0000010110;
    h_3 = 'b0000010111;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000001101;
    x_1 = 'b0000011000;
    x_2 = 'b0000011111;
    x_3 = 'b0000100000;
    x_4 = 'b0000011010;

    h_0 = 'b1111110111;
    h_1 = 'b1111101000;
    h_2 = 'b1111100000;
    h_3 = 'b1111100011;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000100000;
    x_1 = 'b0000001001;
    x_2 = 'b1111100011;
    x_3 = 'b1111101111;
    x_4 = 'b0000011001;

    h_0 = 'b0000000111;
    h_1 = 'b0000010011;
    h_2 = 'b0000011100;
    h_3 = 'b0000100000;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000010101;
    x_1 = 'b1111100000;
    x_2 = 'b0000011011;
    x_3 = 'b1111110110;
    x_4 = 'b1111110100;

    h_0 = 'b0000010101;
    h_1 = 'b0000011011;
    h_2 = 'b1111110010;
    h_3 = 'b1111100001;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111110111;
    x_1 = 'b0000010010;
    x_2 = 'b1111100111;
    x_3 = 'b0000011101;
    x_4 = 'b1111100000;

    h_0 = 'b0000011110;
    h_1 = 'b1111110000;
    h_2 = 'b1111111010;
    h_3 = 'b0000011001;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100001;
    x_1 = 'b0000010001;
    x_2 = 'b0000010101;
    x_3 = 'b1111100011;
    x_4 = 'b1111111010;

    h_0 = 'b0000100000;
    h_1 = 'b1111100011;
    h_2 = 'b0000011000;
    h_3 = 'b1111101111;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111101000;
    x_1 = 'b1111100000;
    x_2 = 'b1111101110;
    x_3 = 'b0000001000;
    x_4 = 'b0000011101;

    h_0 = 'b0000011010;
    h_1 = 'b0000001011;
    h_2 = 'b1111100000;
    h_3 = 'b0000000110;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000000101;
    x_1 = 'b0000001001;
    x_2 = 'b0000001110;
    x_3 = 'b0000010010;
    x_4 = 'b0000010110;

    h_0 = 'b0000001101;
    h_1 = 'b0000011111;
    h_2 = 'b0000011011;
    h_3 = 'b0000000101;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000011101;
    x_1 = 'b0000011000;
    x_2 = 'b1111110110;
    x_3 = 'b1111100000;
    x_4 = 'b1111110000;

    h_0 = 'b1111111110;
    h_1 = 'b1111111001;
    h_2 = 'b1111110100;
    h_3 = 'b1111110000;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000011011;
    x_1 = 'b1111100011;
    x_2 = 'b0000000101;
    x_3 = 'b0000010111;
    x_4 = 'b1111100001;

    h_0 = 'b1111101111;
    h_1 = 'b1111100000;
    h_2 = 'b1111111000;
    h_3 = 'b0000011001;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000000000;
    x_1 = 'b0000000001;
    x_2 = 'b1111111111;
    x_3 = 'b0000000001;
    x_4 = 'b1111111111;

    h_0 = 'b1111100100;
    h_1 = 'b0000000011;
    h_2 = 'b0000011001;
    h_3 = 'b1111100010;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100101;
    x_1 = 'b0000011101;
    x_2 = 'b1111111100;
    x_3 = 'b1111100111;
    x_4 = 'b0000011110;

    h_0 = 'b1111100000;
    h_1 = 'b0000100000;
    h_2 = 'b1111100000;
    h_3 = 'b0000100000;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100011;
    x_1 = 'b1111100111;
    x_2 = 'b0000001000;
    x_3 = 'b0000011111;
    x_4 = 'b0000010011;

    h_0 = 'b1111100100;
    h_1 = 'b0000000010;
    h_2 = 'b0000011010;
    h_3 = 'b1111100010;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111111100;
    x_1 = 'b1111111000;
    x_2 = 'b1111110100;
    x_3 = 'b1111110000;
    x_4 = 'b1111101100;

    h_0 = 'b1111101111;
    h_1 = 'b1111100000;
    h_2 = 'b1111110110;
    h_3 = 'b0000010111;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000011000;
    x_1 = 'b0000100000;
    x_2 = 'b0000010000;
    x_3 = 'b1111110110;
    x_4 = 'b1111100010;

    h_0 = 'b1111111110;
    h_1 = 'b1111111010;
    h_2 = 'b1111110110;
    h_3 = 'b1111110010;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000011111;
    x_1 = 'b1111101110;
    x_2 = 'b1111101100;
    x_3 = 'b0000011110;
    x_4 = 'b0000000011;

    h_0 = 'b0000001101;
    h_1 = 'b0000011111;
    h_2 = 'b0000011010;
    h_3 = 'b0000000011;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000001001;
    x_1 = 'b1111101111;
    x_2 = 'b0000010111;
    x_3 = 'b1111100100;
    x_4 = 'b0000011111;

    h_0 = 'b0000011010;
    h_1 = 'b0000001011;
    h_2 = 'b1111100000;
    h_3 = 'b0000001000;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111101011;
    x_1 = 'b0000100000;
    x_2 = 'b1111100110;
    x_3 = 'b0000001000;
    x_4 = 'b0000001111;

    h_0 = 'b0000100000;
    h_1 = 'b1111100011;
    h_2 = 'b0000011001;
    h_3 = 'b1111101110;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100000;
    x_1 = 'b1111110110;
    x_2 = 'b0000011101;
    x_3 = 'b0000010011;
    x_4 = 'b1111101001;

    h_0 = 'b0000011110;
    h_1 = 'b1111110001;
    h_2 = 'b1111111000;
    h_3 = 'b0000011010;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111110011;
    x_1 = 'b1111101000;
    x_2 = 'b1111100010;
    x_3 = 'b1111100000;
    x_4 = 'b1111100100;

    h_0 = 'b0000010101;
    h_1 = 'b0000011011;
    h_2 = 'b1111110100;
    h_3 = 'b1111100001;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000010010;
    x_1 = 'b0000011101;
    x_2 = 'b0000011111;
    x_3 = 'b0000010111;
    x_4 = 'b0000000111;

    h_0 = 'b0000000111;
    h_1 = 'b0000010011;
    h_2 = 'b0000011100;
    h_3 = 'b0000100000;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000100000;
    x_1 = 'b1111111111;
    x_2 = 'b1111100000;
    x_3 = 'b0000000010;
    x_4 = 'b0000100000;

    h_0 = 'b1111110111;
    h_1 = 'b1111100111;
    h_2 = 'b1111100000;
    h_3 = 'b1111100100;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000010001;
    x_1 = 'b1111100011;
    x_2 = 'b0000100000;
    x_3 = 'b1111100111;
    x_4 = 'b0000001011;

    h_0 = 'b1111101001;
    h_1 = 'b1111101010;
    h_2 = 'b0000010111;
    h_3 = 'b0000010110;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111110010;
    x_1 = 'b0000011001;
    x_2 = 'b1111100001;
    x_3 = 'b0000011111;
    x_4 = 'b1111100110;

    h_0 = 'b1111100001;
    h_1 = 'b0000010101;
    h_2 = 'b1111111010;
    h_3 = 'b1111110100;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100000;
    x_1 = 'b0000001000;
    x_2 = 'b0000011110;
    x_3 = 'b1111110000;
    x_4 = 'b1111100110;

    h_0 = 'b1111100001;
    h_1 = 'b0000011001;
    h_2 = 'b1111110010;
    h_3 = 'b0000000001;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111101011;
    x_1 = 'b1111100000;
    x_2 = 'b1111100100;
    x_3 = 'b1111110101;
    x_4 = 'b0000001011;

    h_0 = 'b1111101000;
    h_1 = 'b1111101110;
    h_2 = 'b0000011101;
    h_3 = 'b0000001011;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000001001;
    x_1 = 'b0000010010;
    x_2 = 'b0000011001;
    x_3 = 'b0000011110;
    x_4 = 'b0000100000;

    h_0 = 'b1111110101;
    h_1 = 'b1111100100;
    h_2 = 'b1111100000;
    h_3 = 'b1111101100;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000011111;
    x_1 = 'b0000010000;
    x_2 = 'b1111101010;
    x_3 = 'b1111100100;
    x_4 = 'b0000000111;

    h_0 = 'b0000000101;
    h_1 = 'b0000001110;
    h_2 = 'b0000010110;
    h_3 = 'b0000011100;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000011000;
    x_1 = 'b1111100000;
    x_2 = 'b0000010011;
    x_3 = 'b0000000111;
    x_4 = 'b1111100100;

    h_0 = 'b0000010011;
    h_1 = 'b0000011110;
    h_2 = 'b1111111100;
    h_3 = 'b1111100000;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111111011;
    x_1 = 'b0000001010;
    x_2 = 'b1111110001;
    x_3 = 'b0000010011;
    x_4 = 'b1111101001;

    h_0 = 'b0000011101;
    h_1 = 'b1111110110;
    h_2 = 'b1111110000;
    h_3 = 'b0000011111;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100011;
    x_1 = 'b0000010111;
    x_2 = 'b0000001011;
    x_3 = 'b1111100000;
    x_4 = 'b0000001111;

    h_0 = 'b0000100000;
    h_1 = 'b1111100001;
    h_2 = 'b0000011101;
    h_3 = 'b1111100101;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100101;
    x_1 = 'b1111100010;
    x_2 = 'b1111111010;
    x_3 = 'b0000010111;
    x_4 = 'b0000011111;

    h_0 = 'b0000011011;
    h_1 = 'b0000000101;
    h_2 = 'b1111100001;
    h_3 = 'b0000010011;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000000001;
    x_1 = 'b0000000001;
    x_2 = 'b0000000010;
    x_3 = 'b0000000010;
    x_4 = 'b0000000011;

    h_0 = 'b0000001111;
    h_1 = 'b0000100000;
    h_2 = 'b0000010100;
    h_3 = 'b1111110111;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000011011;
    x_1 = 'b0000011101;
    x_2 = 'b0000000011;
    x_3 = 'b1111100110;
    x_4 = 'b1111100010;

    h_0 = 'b0000000000;
    h_1 = 'b1111111111;
    h_2 = 'b1111111111;
    h_3 = 'b1111111110;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000011101;
    x_1 = 'b1111100111;
    x_2 = 'b1111111001;
    x_3 = 'b0000011111;
    x_4 = 'b1111101100;

    h_0 = 'b1111110000;
    h_1 = 'b1111100000;
    h_2 = 'b1111101110;
    h_3 = 'b0000001101;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000000100;
    x_1 = 'b1111111000;
    x_2 = 'b0000001100;
    x_3 = 'b1111110001;
    x_4 = 'b0000010011;

    h_0 = 'b1111100101;
    h_1 = 'b1111111100;
    h_2 = 'b0000011110;
    h_3 = 'b1111101010;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100111;
    x_1 = 'b0000011111;
    x_2 = 'b1111110000;
    x_3 = 'b1111110101;
    x_4 = 'b0000011110;

    h_0 = 'b1111100000;
    h_1 = 'b0000011111;
    h_2 = 'b1111100010;
    h_3 = 'b0000011101;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100001;
    x_1 = 'b1111101110;
    x_2 = 'b0000010011;
    x_3 = 'b0000011110;
    x_4 = 'b1111111111;

    h_0 = 'b1111100011;
    h_1 = 'b0000001000;
    h_2 = 'b0000010011;
    h_3 = 'b1111100000;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111111000;
    x_1 = 'b1111110000;
    x_2 = 'b1111101001;
    x_3 = 'b1111100100;
    x_4 = 'b1111100001;

    h_0 = 'b1111101101;
    h_1 = 'b1111100010;
    h_2 = 'b0000000001;
    h_3 = 'b0000011111;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000010101;
    x_1 = 'b0000100000;
    x_2 = 'b0000011010;
    x_3 = 'b0000000110;
    x_4 = 'b1111110000;

    h_0 = 'b1111111100;
    h_1 = 'b1111110100;
    h_2 = 'b1111101100;
    h_3 = 'b1111100110;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000100000;
    x_1 = 'b1111110110;
    x_2 = 'b1111100100;
    x_3 = 'b0000010011;
    x_4 = 'b0000010110;

    h_0 = 'b0000001011;
    h_1 = 'b0000011101;
    h_2 = 'b0000011111;
    h_3 = 'b0000010001;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000001101;
    x_1 = 'b1111101001;
    x_2 = 'b0000011110;
    x_3 = 'b1111100000;
    x_4 = 'b0000011101;

    h_0 = 'b0000011000;
    h_1 = 'b0000010000;
    h_2 = 'b1111100010;
    h_3 = 'b1111111001;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111101110;
    x_1 = 'b0000011110;
    x_2 = 'b1111100001;
    x_3 = 'b0000010110;
    x_4 = 'b1111111010;

    h_0 = 'b0000011111;
    h_1 = 'b1111100110;
    h_2 = 'b0000010001;
    h_3 = 'b1111111011;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100000;
    x_1 = 'b1111111111;
    x_2 = 'b0000100000;
    x_3 = 'b0000000011;
    x_4 = 'b1111100000;

    h_0 = 'b0000011111;
    h_1 = 'b1111101100;
    h_2 = 'b0000000011;
    h_3 = 'b0000001111;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111101111;
    x_1 = 'b1111100100;
    x_2 = 'b1111100000;
    x_3 = 'b1111100110;
    x_4 = 'b1111110100;

    h_0 = 'b0000010110;
    h_1 = 'b0000010111;
    h_2 = 'b1111101011;
    h_3 = 'b1111101000;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000001110;
    x_1 = 'b0000011001;
    x_2 = 'b0000011111;
    x_3 = 'b0000011111;
    x_4 = 'b0000011001;

    h_0 = 'b0000001001;
    h_1 = 'b0000010111;
    h_2 = 'b0000011111;
    h_3 = 'b0000011110;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000100000;
    x_1 = 'b0000001000;
    x_2 = 'b1111100010;
    x_3 = 'b1111110001;
    x_4 = 'b0000011010;

    h_0 = 'b1111111001;
    h_1 = 'b1111101100;
    h_2 = 'b1111100011;
    h_3 = 'b1111100000;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000010100;
    x_1 = 'b1111100001;
    x_2 = 'b0000011100;
    x_3 = 'b1111110100;
    x_4 = 'b1111110110;

    h_0 = 'b1111101011;
    h_1 = 'b1111100110;
    h_2 = 'b0000001111;
    h_3 = 'b0000011110;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111110110;
    x_1 = 'b0000010011;
    x_2 = 'b1111100110;
    x_3 = 'b0000011110;
    x_4 = 'b1111100000;

    h_0 = 'b1111100010;
    h_1 = 'b0000010000;
    h_2 = 'b0000000101;
    h_3 = 'b1111101000;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100001;
    x_1 = 'b0000010000;
    x_2 = 'b0000010111;
    x_3 = 'b1111100100;
    x_4 = 'b1111111000;

    h_0 = 'b1111100000;
    h_1 = 'b0000011101;
    h_2 = 'b1111101001;
    h_3 = 'b0000001111;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111101000;
    x_1 = 'b1111100000;
    x_2 = 'b1111101101;
    x_3 = 'b0000000110;
    x_4 = 'b0000011011;

    h_0 = 'b1111100111;
    h_1 = 'b1111110100;
    h_2 = 'b0000100000;
    h_3 = 'b1111111100;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000000101;
    x_1 = 'b0000001011;
    x_2 = 'b0000001111;
    x_3 = 'b0000010100;
    x_4 = 'b0000011000;

    h_0 = 'b1111110011;
    h_1 = 'b1111100010;
    h_2 = 'b1111100100;
    h_3 = 'b1111111001;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000011101;
    x_1 = 'b0000010111;
    x_2 = 'b1111110101;
    x_3 = 'b1111100000;
    x_4 = 'b1111110010;

    h_0 = 'b0000000011;
    h_1 = 'b0000001000;
    h_2 = 'b0000001101;
    h_3 = 'b0000010010;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000011010;
    x_1 = 'b1111100010;
    x_2 = 'b0000000111;
    x_3 = 'b0000010110;
    x_4 = 'b1111100000;

    h_0 = 'b0000010010;
    h_1 = 'b0000011111;
    h_2 = 'b0000000111;
    h_3 = 'b1111100110;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111111111;
    x_1 = 'b0000000010;
    x_2 = 'b1111111101;
    x_3 = 'b0000000011;
    x_4 = 'b1111111100;

    h_0 = 'b0000011100;
    h_1 = 'b1111111100;
    h_2 = 'b1111101000;
    h_3 = 'b0000011111;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100101;
    x_1 = 'b0000011100;
    x_2 = 'b1111111110;
    x_3 = 'b1111100110;
    x_4 = 'b0000011101;

    h_0 = 'b0000100000;
    h_1 = 'b1111100000;
    h_2 = 'b0000100000;
    h_3 = 'b1111100000;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100011;
    x_1 = 'b1111100111;
    x_2 = 'b0000000110;
    x_3 = 'b0000011111;
    x_4 = 'b0000010101;

    h_0 = 'b0000011100;
    h_1 = 'b1111111111;
    h_2 = 'b1111100101;
    h_3 = 'b0000011101;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111111100;
    x_1 = 'b1111111001;
    x_2 = 'b1111110101;
    x_3 = 'b1111110010;
    x_4 = 'b1111101111;

    h_0 = 'b0000010001;
    h_1 = 'b0000100000;
    h_2 = 'b0000001011;
    h_3 = 'b1111101010;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000011001;
    x_1 = 'b0000011111;
    x_2 = 'b0000001111;
    x_3 = 'b1111110100;
    x_4 = 'b1111100001;

    h_0 = 'b0000000010;
    h_1 = 'b0000000101;
    h_2 = 'b0000001001;
    h_3 = 'b0000001101;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000011110;
    x_1 = 'b1111101101;
    x_2 = 'b1111101101;
    x_3 = 'b0000011110;
    x_4 = 'b0000000000;

    h_0 = 'b1111110010;
    h_1 = 'b1111100001;
    h_2 = 'b1111100110;
    h_3 = 'b1111111111;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000001000;
    x_1 = 'b1111110000;
    x_2 = 'b0000010110;
    x_3 = 'b1111100101;
    x_4 = 'b0000011111;

    h_0 = 'b1111100110;
    h_1 = 'b1111110110;
    h_2 = 'b0000100000;
    h_3 = 'b1111110110;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111101010;
    x_1 = 'b0000100000;
    x_2 = 'b1111100111;
    x_3 = 'b0000000101;
    x_4 = 'b0000010001;

    h_0 = 'b1111100000;
    h_1 = 'b0000011110;
    h_2 = 'b1111100110;
    h_3 = 'b0000010100;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100000;
    x_1 = 'b1111110101;
    x_2 = 'b0000011100;
    x_3 = 'b0000010100;
    x_4 = 'b1111101011;

    h_0 = 'b1111100010;
    h_1 = 'b0000001110;
    h_2 = 'b0000001001;
    h_3 = 'b1111100101;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111110100;
    x_1 = 'b1111101001;
    x_2 = 'b1111100010;
    x_3 = 'b1111100000;
    x_4 = 'b1111100011;

    h_0 = 'b1111101011;
    h_1 = 'b1111100100;
    h_2 = 'b0000001011;
    h_3 = 'b0000011111;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000010010;
    x_1 = 'b0000011110;
    x_2 = 'b0000011111;
    x_3 = 'b0000010101;
    x_4 = 'b0000000100;

    h_0 = 'b1111111010;
    h_1 = 'b1111101110;
    h_2 = 'b1111100101;
    h_3 = 'b1111100001;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000100000;
    x_1 = 'b1111111110;
    x_2 = 'b1111100000;
    x_3 = 'b0000000100;
    x_4 = 'b0000100000;

    h_0 = 'b0000001001;
    h_1 = 'b0000011001;
    h_2 = 'b0000100000;
    h_3 = 'b0000011100;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000010000;
    x_1 = 'b1111100100;
    x_2 = 'b0000100000;
    x_3 = 'b1111100101;
    x_4 = 'b0000001110;

    h_0 = 'b0000010111;
    h_1 = 'b0000010110;
    h_2 = 'b1111101000;
    h_3 = 'b1111101100;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111110010;
    x_1 = 'b0000011001;
    x_2 = 'b1111100001;
    x_3 = 'b0000011111;
    x_4 = 'b1111101000;

    h_0 = 'b0000011111;
    h_1 = 'b1111101010;
    h_2 = 'b0000000111;
    h_3 = 'b0000001010;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100000;
    x_1 = 'b0000000111;
    x_2 = 'b0000011110;
    x_3 = 'b1111110010;
    x_4 = 'b1111100101;

    h_0 = 'b0000011111;
    h_1 = 'b1111100111;
    h_2 = 'b0000001101;
    h_3 = 'b0000000001;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111101100;
    x_1 = 'b1111100001;
    x_2 = 'b1111100100;
    x_3 = 'b1111110011;
    x_4 = 'b0000001000;

    h_0 = 'b0000011000;
    h_1 = 'b0000010011;
    h_2 = 'b1111100100;
    h_3 = 'b1111110100;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000001010;
    x_1 = 'b0000010011;
    x_2 = 'b0000011010;
    x_3 = 'b0000011111;
    x_4 = 'b0000100000;

    h_0 = 'b0000001011;
    h_1 = 'b0000011011;
    h_2 = 'b0000100000;
    h_3 = 'b0000010110;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000011111;
    x_1 = 'b0000001111;
    x_2 = 'b1111101001;
    x_3 = 'b1111100101;
    x_4 = 'b0000001010;

    h_0 = 'b1111111011;
    h_1 = 'b1111110001;
    h_2 = 'b1111101001;
    h_3 = 'b1111100011;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000010111;
    x_1 = 'b1111100000;
    x_2 = 'b0000010100;
    x_3 = 'b0000000101;
    x_4 = 'b1111100110;

    h_0 = 'b1111101100;
    h_1 = 'b1111100011;
    h_2 = 'b0000000101;
    h_3 = 'b0000100000;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111111010;
    x_1 = 'b0000001011;
    x_2 = 'b1111110000;
    x_3 = 'b0000010101;
    x_4 = 'b1111100111;

    h_0 = 'b1111100011;
    h_1 = 'b0000001011;
    h_2 = 'b0000001111;
    h_3 = 'b1111100001;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100010;
    x_1 = 'b0000010111;
    x_2 = 'b0000001100;
    x_3 = 'b1111100000;
    x_4 = 'b0000001100;

    h_0 = 'b1111100000;
    h_1 = 'b0000011111;
    h_2 = 'b1111100011;
    h_3 = 'b0000011010;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100110;
    x_1 = 'b1111100010;
    x_2 = 'b1111111000;
    x_3 = 'b0000010101;
    x_4 = 'b0000100000;

    h_0 = 'b1111100101;
    h_1 = 'b1111111010;
    h_2 = 'b0000011111;
    h_3 = 'b1111101110;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000000001;
    x_1 = 'b0000000010;
    x_2 = 'b0000000011;
    x_3 = 'b0000000101;
    x_4 = 'b0000000110;

    h_0 = 'b1111110001;
    h_1 = 'b1111100000;
    h_2 = 'b1111101011;
    h_3 = 'b0000000111;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000011100;
    x_1 = 'b0000011100;
    x_2 = 'b0000000001;
    x_3 = 'b1111100101;
    x_4 = 'b1111100011;

    h_0 = 'b0000000001;
    h_1 = 'b0000000010;
    h_2 = 'b0000000011;
    h_3 = 'b0000000100;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000011101;
    x_1 = 'b1111100110;
    x_2 = 'b1111111010;
    x_3 = 'b0000011111;
    x_4 = 'b1111101010;

    h_0 = 'b0000010000;
    h_1 = 'b0000100000;
    h_2 = 'b0000010001;
    h_3 = 'b1111110001;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000000011;
    x_1 = 'b1111111001;
    x_2 = 'b0000001010;
    x_3 = 'b1111110011;
    x_4 = 'b0000010000;

    h_0 = 'b0000011011;
    h_1 = 'b0000000011;
    h_2 = 'b1111100010;
    h_3 = 'b0000011000;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100111;
    x_1 = 'b0000011111;
    x_2 = 'b1111110010;
    x_3 = 'b1111110011;
    x_4 = 'b0000011111;

    h_0 = 'b0000100000;
    h_1 = 'b1111100000;
    h_2 = 'b0000011111;
    h_3 = 'b1111100010;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100010;
    x_1 = 'b1111101101;
    x_2 = 'b0000010010;
    x_3 = 'b0000011111;
    x_4 = 'b0000000001;

    h_0 = 'b0000011101;
    h_1 = 'b1111111001;
    h_2 = 'b1111101100;
    h_3 = 'b0000100000;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111111000;
    x_1 = 'b1111110001;
    x_2 = 'b1111101010;
    x_3 = 'b1111100101;
    x_4 = 'b1111100010;

    h_0 = 'b0000010011;
    h_1 = 'b0000011111;
    h_2 = 'b0000000001;
    h_3 = 'b1111100010;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000010110;
    x_1 = 'b0000100000;
    x_2 = 'b0000011001;
    x_3 = 'b0000000100;
    x_4 = 'b1111101101;

    h_0 = 'b0000000100;
    h_1 = 'b0000001100;
    h_2 = 'b0000010011;
    h_3 = 'b0000011000;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000011111;
    x_1 = 'b1111110101;
    x_2 = 'b1111100101;
    x_3 = 'b0000010101;
    x_4 = 'b0000010100;

    h_0 = 'b1111110100;
    h_1 = 'b1111100011;
    h_2 = 'b1111100010;
    h_3 = 'b1111110000;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000001100;
    x_1 = 'b1111101010;
    x_2 = 'b0000011101;
    x_3 = 'b1111100000;
    x_4 = 'b0000011110;

    h_0 = 'b1111100111;
    h_1 = 'b1111110000;
    h_2 = 'b0000011110;
    h_3 = 'b0000000101;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111101110;
    x_1 = 'b0000011110;
    x_2 = 'b1111100001;
    x_3 = 'b0000010101;
    x_4 = 'b1111111101;

    h_0 = 'b1111100001;
    h_1 = 'b0000011011;
    h_2 = 'b1111101110;
    h_3 = 'b0000000111;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111100000;
    x_1 = 'b1111111101;
    x_2 = 'b0000100000;
    x_3 = 'b0000000101;
    x_4 = 'b1111100001;

    h_0 = 'b1111100001;
    h_1 = 'b0000010011;
    h_2 = 'b1111111111;
    h_3 = 'b1111101111;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b1111110000;
    x_1 = 'b1111100100;
    x_2 = 'b1111100000;
    x_3 = 'b1111100101;
    x_4 = 'b1111110001;

    h_0 = 'b1111101010;
    h_1 = 'b1111101000;
    h_2 = 'b0000010100;
    h_3 = 'b0000011010;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    x_0 = 'b0000001110;
    x_1 = 'b0000011010;
    x_2 = 'b0000100000;
    x_3 = 'b0000011111;
    x_4 = 'b0000010111;

    h_0 = 'b1111111000;
    h_1 = 'b1111101001;
    h_2 = 'b1111100001;
    h_3 = 'b1111100001;
    #20;
    $fdisplay(fd, "%010b %010b %010b %010b", y_0, y_1, y_2, y_3);

    $fclose(fd);    
$finish;
    end
endmodule