`timescale 1ns / 1ps

module gru_tb;

// Parameters
parameter int INT_WIDTH  = 4;
parameter int FRAC_WIDTH = 10;
parameter int WIDTH      = INT_WIDTH + FRAC_WIDTH + 1;
parameter real CLK_PERIOD = 10.0;

// Clock and reset
logic clk;
logic reset;

// Inputs
logic signed [WIDTH-1:0] x_0 = 0;
logic signed [WIDTH-1:0] x_1 = 0;
logic signed [WIDTH-1:0] x_2 = 0;
logic signed [WIDTH-1:0] x_3 = 0;

logic signed [WIDTH-1:0] h_0 = 0;
logic signed [WIDTH-1:0] h_1 = 0;
logic signed [WIDTH-1:0] h_2 = 0;
logic signed [WIDTH-1:0] h_3 = 0;

// Input weights (h×d for each gate)
logic signed [WIDTH-1:0] w_ir_0_0 = 'b00000001010010;
logic signed [WIDTH-1:0] w_ir_0_1 = 'b00000010011100;
logic signed [WIDTH-1:0] w_ir_0_2 = 'b00000001110111;
logic signed [WIDTH-1:0] w_ir_0_3 = 'b00000010001101;
logic signed [WIDTH-1:0] w_ir_1_0 = 'b11111110110101;
logic signed [WIDTH-1:0] w_ir_1_1 = 'b11111101010101;
logic signed [WIDTH-1:0] w_ir_1_2 = 'b00000001110011;
logic signed [WIDTH-1:0] w_ir_1_3 = 'b00000000111110;
logic signed [WIDTH-1:0] w_ir_2_0 = 'b11111100100001;
logic signed [WIDTH-1:0] w_ir_2_1 = 'b00000000010110;
logic signed [WIDTH-1:0] w_ir_2_2 = 'b00000011111011;
logic signed [WIDTH-1:0] w_ir_2_3 = 'b11111111111111;
logic signed [WIDTH-1:0] w_ir_3_0 = 'b00000010100000;
logic signed [WIDTH-1:0] w_ir_3_1 = 'b00000000101100;
logic signed [WIDTH-1:0] w_ir_3_2 = 'b00000000100111;
logic signed [WIDTH-1:0] w_ir_3_3 = 'b00000010111001;

logic signed [WIDTH-1:0] w_iz_0_0 = 'b11111111100000;
logic signed [WIDTH-1:0] w_iz_0_1 = 'b00000011011101;
logic signed [WIDTH-1:0] w_iz_0_2 = 'b11111111100011;
logic signed [WIDTH-1:0] w_iz_0_3 = 'b00000010010001;
logic signed [WIDTH-1:0] w_iz_1_0 = 'b11111111100010;
logic signed [WIDTH-1:0] w_iz_1_1 = 'b00000010000111;
logic signed [WIDTH-1:0] w_iz_1_2 = 'b00000001100010;
logic signed [WIDTH-1:0] w_iz_1_3 = 'b00000001100011;
logic signed [WIDTH-1:0] w_iz_2_0 = 'b11111101011111;
logic signed [WIDTH-1:0] w_iz_2_1 = 'b00000001111000;
logic signed [WIDTH-1:0] w_iz_2_2 = 'b00000010001100;
logic signed [WIDTH-1:0] w_iz_2_3 = 'b00000001011011;
logic signed [WIDTH-1:0] w_iz_3_0 = 'b00000011100011;
logic signed [WIDTH-1:0] w_iz_3_1 = 'b11111100101100;
logic signed [WIDTH-1:0] w_iz_3_2 = 'b11111110110110;
logic signed [WIDTH-1:0] w_iz_3_3 = 'b00000001100111;

logic signed [WIDTH-1:0] w_in_0_0 = 'b00000000110010;
logic signed [WIDTH-1:0] w_in_0_1 = 'b00000001111010;
logic signed [WIDTH-1:0] w_in_0_2 = 'b00000001111010;
logic signed [WIDTH-1:0] w_in_0_3 = 'b00000000011011;
logic signed [WIDTH-1:0] w_in_1_0 = 'b00000011111111;
logic signed [WIDTH-1:0] w_in_1_1 = 'b00000001010001;
logic signed [WIDTH-1:0] w_in_1_2 = 'b11111110111011;
logic signed [WIDTH-1:0] w_in_1_3 = 'b00000000111110;
logic signed [WIDTH-1:0] w_in_2_0 = 'b00000010010110;
logic signed [WIDTH-1:0] w_in_2_1 = 'b11111101000001;
logic signed [WIDTH-1:0] w_in_2_2 = 'b00000000111101;
logic signed [WIDTH-1:0] w_in_2_3 = 'b11111110100001;
logic signed [WIDTH-1:0] w_in_3_0 = 'b11111111111001;
logic signed [WIDTH-1:0] w_in_3_1 = 'b11111101110011;
logic signed [WIDTH-1:0] w_in_3_2 = 'b11111100111010;
logic signed [WIDTH-1:0] w_in_3_3 = 'b00000011011111;

// Recurrent weights (h×h for each gate)
logic signed [WIDTH-1:0] w_hr_0_0 = 'b00000000001110;
logic signed [WIDTH-1:0] w_hr_0_1 = 'b00000000100111;
logic signed [WIDTH-1:0] w_hr_0_2 = 'b00000000111110;
logic signed [WIDTH-1:0] w_hr_0_3 = 'b11111101011100;
logic signed [WIDTH-1:0] w_hr_1_0 = 'b00000100011000;
logic signed [WIDTH-1:0] w_hr_1_1 = 'b00000100101101;
logic signed [WIDTH-1:0] w_hr_1_2 = 'b00000100101011;
logic signed [WIDTH-1:0] w_hr_1_3 = 'b11111011011000;
logic signed [WIDTH-1:0] w_hr_2_0 = 'b00000011111110;
logic signed [WIDTH-1:0] w_hr_2_1 = 'b00000100100000;
logic signed [WIDTH-1:0] w_hr_2_2 = 'b11111101111110;
logic signed [WIDTH-1:0] w_hr_2_3 = 'b11111101100011;
logic signed [WIDTH-1:0] w_hr_3_0 = 'b00000001111101;
logic signed [WIDTH-1:0] w_hr_3_1 = 'b00000010100000;
logic signed [WIDTH-1:0] w_hr_3_2 = 'b00000101101000;
logic signed [WIDTH-1:0] w_hr_3_3 = 'b11111100001101;

logic signed [WIDTH-1:0] w_hz_0_0 = 'b00000011011100;
logic signed [WIDTH-1:0] w_hz_0_1 = 'b00000001110010;
logic signed [WIDTH-1:0] w_hz_0_2 = 'b11111110101100;
logic signed [WIDTH-1:0] w_hz_0_3 = 'b00000010000010;
logic signed [WIDTH-1:0] w_hz_1_0 = 'b00000110100001;
logic signed [WIDTH-1:0] w_hz_1_1 = 'b11111001111001;
logic signed [WIDTH-1:0] w_hz_1_2 = 'b00000000000111;
logic signed [WIDTH-1:0] w_hz_1_3 = 'b00000100011111;
logic signed [WIDTH-1:0] w_hz_2_0 = 'b00000011011001;
logic signed [WIDTH-1:0] w_hz_2_1 = 'b00000000000101;
logic signed [WIDTH-1:0] w_hz_2_2 = 'b11111000001010;
logic signed [WIDTH-1:0] w_hz_2_3 = 'b00000111000111;
logic signed [WIDTH-1:0] w_hz_3_0 = 'b00000101111111;
logic signed [WIDTH-1:0] w_hz_3_1 = 'b00000010001011;
logic signed [WIDTH-1:0] w_hz_3_2 = 'b11111011010011;
logic signed [WIDTH-1:0] w_hz_3_3 = 'b00001010010111;

logic signed [WIDTH-1:0] w_hn_0_0 = 'b11111111010111;
logic signed [WIDTH-1:0] w_hn_0_1 = 'b11111110110011;
logic signed [WIDTH-1:0] w_hn_0_2 = 'b00000010010010;
logic signed [WIDTH-1:0] w_hn_0_3 = 'b11111100110001;
logic signed [WIDTH-1:0] w_hn_1_0 = 'b11111101001011;
logic signed [WIDTH-1:0] w_hn_1_1 = 'b11111111100111;
logic signed [WIDTH-1:0] w_hn_1_2 = 'b00001011101110;
logic signed [WIDTH-1:0] w_hn_1_3 = 'b11111010001000;
logic signed [WIDTH-1:0] w_hn_2_0 = 'b11111111010111;
logic signed [WIDTH-1:0] w_hn_2_1 = 'b00000110110100;
logic signed [WIDTH-1:0] w_hn_2_2 = 'b00001001111100;
logic signed [WIDTH-1:0] w_hn_2_3 = 'b11111001000001;
logic signed [WIDTH-1:0] w_hn_3_0 = 'b11111101011001;
logic signed [WIDTH-1:0] w_hn_3_1 = 'b11111011001100;
logic signed [WIDTH-1:0] w_hn_3_2 = 'b11111100101110;
logic signed [WIDTH-1:0] w_hn_3_3 = 'b00000100111011;

// Biases (h for each gate type)
logic signed [WIDTH-1:0] b_ir_0 = 'b00000000010111;
logic signed [WIDTH-1:0] b_ir_1 = 'b00000100001011;
logic signed [WIDTH-1:0] b_ir_2 = 'b00000111011011;
logic signed [WIDTH-1:0] b_ir_3 = 'b00000010100011;

logic signed [WIDTH-1:0] b_iz_0 = 'b00000011000010;
logic signed [WIDTH-1:0] b_iz_1 = 'b00000010001001;
logic signed [WIDTH-1:0] b_iz_2 = 'b00000111111001;
logic signed [WIDTH-1:0] b_iz_3 = 'b11111111110100;

logic signed [WIDTH-1:0] b_in_0 = 'b00000101010100;
logic signed [WIDTH-1:0] b_in_1 = 'b00000000111010;
logic signed [WIDTH-1:0] b_in_2 = 'b00000111000010;
logic signed [WIDTH-1:0] b_in_3 = 'b00000001001100;

logic signed [WIDTH-1:0] b_hr_0 = 'b00000001001001;
logic signed [WIDTH-1:0] b_hr_1 = 'b00000100111001;
logic signed [WIDTH-1:0] b_hr_2 = 'b00000011011100;
logic signed [WIDTH-1:0] b_hr_3 = 'b00000110100011;

logic signed [WIDTH-1:0] b_hz_0 = 'b00000011010001;
logic signed [WIDTH-1:0] b_hz_1 = 'b00000100100101;
logic signed [WIDTH-1:0] b_hz_2 = 'b00000010100000;
logic signed [WIDTH-1:0] b_hz_3 = 'b00001100111011;

logic signed [WIDTH-1:0] b_hn_0 = 'b00000001100001;
logic signed [WIDTH-1:0] b_hn_1 = 'b00001001100000;
logic signed [WIDTH-1:0] b_hn_2 = 'b00000011101010;
logic signed [WIDTH-1:0] b_hn_3 = 'b11111000010001;

// Outputs (h=4)
logic signed [WIDTH-1:0]  y_0 = 0;
logic signed [WIDTH-1:0]  y_1 = 0;
logic signed [WIDTH-1:0]  y_2 = 0;
logic signed [WIDTH-1:0]  y_3 = 0;

gru #(
        .INT_WIDTH(INT_WIDTH),
        .FRAC_WIDTH(FRAC_WIDTH)
    ) gru_inst (
        .clk(clk),
        .reset(reset),
        // Input features (d=64)
        	
.x_0(x_0), .x_1(x_1), .x_2(x_2), .x_3(x_3), 	
.h_0(h_0), .h_1(h_1), .h_2(h_2), .h_3(h_3), 	
.w_ir_0_0(w_ir_0_0), .w_ir_0_1(w_ir_0_1), .w_ir_0_2(w_ir_0_2), .w_ir_0_3(w_ir_0_3), .w_ir_1_0(w_ir_1_0), .w_ir_1_1(w_ir_1_1), .w_ir_1_2(w_ir_1_2), .w_ir_1_3(w_ir_1_3), .w_ir_2_0(w_ir_2_0), .w_ir_2_1(w_ir_2_1), .w_ir_2_2(w_ir_2_2), .w_ir_2_3(w_ir_2_3), .w_ir_3_0(w_ir_3_0), .w_ir_3_1(w_ir_3_1), .w_ir_3_2(w_ir_3_2), .w_ir_3_3(w_ir_3_3), 	
.w_iz_0_0(w_iz_0_0), .w_iz_0_1(w_iz_0_1), .w_iz_0_2(w_iz_0_2), .w_iz_0_3(w_iz_0_3), .w_iz_1_0(w_iz_1_0), .w_iz_1_1(w_iz_1_1), .w_iz_1_2(w_iz_1_2), .w_iz_1_3(w_iz_1_3), .w_iz_2_0(w_iz_2_0), .w_iz_2_1(w_iz_2_1), .w_iz_2_2(w_iz_2_2), .w_iz_2_3(w_iz_2_3), .w_iz_3_0(w_iz_3_0), .w_iz_3_1(w_iz_3_1), .w_iz_3_2(w_iz_3_2), .w_iz_3_3(w_iz_3_3), 
.w_in_0_0(w_in_0_0), .w_in_0_1(w_in_0_1), .w_in_0_2(w_in_0_2), .w_in_0_3(w_in_0_3), .w_in_1_0(w_in_1_0), .w_in_1_1(w_in_1_1), .w_in_1_2(w_in_1_2), .w_in_1_3(w_in_1_3), .w_in_2_0(w_in_2_0), .w_in_2_1(w_in_2_1), .w_in_2_2(w_in_2_2), .w_in_2_3(w_in_2_3), .w_in_3_0(w_in_3_0), .w_in_3_1(w_in_3_1), .w_in_3_2(w_in_3_2), .w_in_3_3(w_in_3_3), 
.w_hr_0_0(w_hr_0_0), .w_hr_0_1(w_hr_0_1), .w_hr_0_2(w_hr_0_2), .w_hr_0_3(w_hr_0_3), .w_hr_1_0(w_hr_1_0), .w_hr_1_1(w_hr_1_1), .w_hr_1_2(w_hr_1_2), .w_hr_1_3(w_hr_1_3), .w_hr_2_0(w_hr_2_0), .w_hr_2_1(w_hr_2_1), .w_hr_2_2(w_hr_2_2), .w_hr_2_3(w_hr_2_3), .w_hr_3_0(w_hr_3_0), .w_hr_3_1(w_hr_3_1), .w_hr_3_2(w_hr_3_2), .w_hr_3_3(w_hr_3_3), 
.w_hz_0_0(w_hz_0_0), .w_hz_0_1(w_hz_0_1), .w_hz_0_2(w_hz_0_2), .w_hz_0_3(w_hz_0_3), .w_hz_1_0(w_hz_1_0), .w_hz_1_1(w_hz_1_1), .w_hz_1_2(w_hz_1_2), .w_hz_1_3(w_hz_1_3), .w_hz_2_0(w_hz_2_0), .w_hz_2_1(w_hz_2_1), .w_hz_2_2(w_hz_2_2), .w_hz_2_3(w_hz_2_3), .w_hz_3_0(w_hz_3_0), .w_hz_3_1(w_hz_3_1), .w_hz_3_2(w_hz_3_2), .w_hz_3_3(w_hz_3_3), 
.w_hn_0_0(w_hn_0_0), .w_hn_0_1(w_hn_0_1), .w_hn_0_2(w_hn_0_2), .w_hn_0_3(w_hn_0_3), .w_hn_1_0(w_hn_1_0), .w_hn_1_1(w_hn_1_1), .w_hn_1_2(w_hn_1_2), .w_hn_1_3(w_hn_1_3), .w_hn_2_0(w_hn_2_0), .w_hn_2_1(w_hn_2_1), .w_hn_2_2(w_hn_2_2), .w_hn_2_3(w_hn_2_3), .w_hn_3_0(w_hn_3_0), .w_hn_3_1(w_hn_3_1), .w_hn_3_2(w_hn_3_2), .w_hn_3_3(w_hn_3_3), 
.b_ir_0(b_ir_0), .b_ir_1(b_ir_1), .b_ir_2(b_ir_2), .b_ir_3(b_ir_3), 
.b_iz_0(b_iz_0), .b_iz_1(b_iz_1), .b_iz_2(b_iz_2), .b_iz_3(b_iz_3), 
.b_in_0(b_in_0), .b_in_1(b_in_1), .b_in_2(b_in_2), .b_in_3(b_in_3), 
.b_hr_0(b_hr_0), .b_hr_1(b_hr_1), .b_hr_2(b_hr_2), .b_hr_3(b_hr_3), 
.b_hz_0(b_hz_0), .b_hz_1(b_hz_1), .b_hz_2(b_hz_2), .b_hz_3(b_hz_3), 
.b_hn_0(b_hn_0), .b_hn_1(b_hn_1), .b_hn_2(b_hn_2), .b_hn_3(b_hn_3), 
.y_0(y_0), .y_1(y_1), .y_2(y_2), .y_3(y_3)
);

    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end
    
    initial begin
        // Open file for writing (overwrite existing)
        integer fd;
        fd = $fopen("../../../../../output_d4_h4_int4_frac10.txt", "w+");
        if (fd == 0) begin
            $display("ERROR: Failed to open file!");
            $finish;
        end
        x_0 = 'b00001110100011;
    x_1 = 'b11110011111001;
    x_2 = 'b11111011100010;
    x_3 = 'b00001111110101;

    h_0 = 'b00000111101011;
    h_1 = 'b00001111111101;
    h_2 = 'b00001001100101;
    h_3 = 'b11111010011001;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00000010010001;
    x_1 = 'b11111011100010;
    x_2 = 'b00000110100110;
    x_3 = 'b11110111011011;

    h_0 = 'b00001101011110;
    h_1 = 'b00000010010001;
    h_2 = 'b11110000101010;
    h_3 = 'b00001010100001;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110011111001;
    x_1 = 'b00001111110101;
    x_2 = 'b11110111011011;
    x_3 = 'b11111011011001;

    h_0 = 'b00001111111101;
    h_1 = 'b11110000010111;
    h_2 = 'b00001111000001;
    h_3 = 'b11110001111011;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110000101010;
    x_1 = 'b11110111010011;
    x_2 = 'b00001010011010;
    x_3 = 'b00001110100111;

    h_0 = 'b00001110100011;
    h_1 = 'b11111011100010;
    h_2 = 'b11110111010011;
    h_3 = 'b00001111110110;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11111011100010;
    x_1 = 'b11110111011011;
    x_2 = 'b11110011111111;
    x_3 = 'b11110001100001;

    h_0 = 'b00001001100101;
    h_1 = 'b00001111000001;
    h_2 = 'b11111110111100;
    h_3 = 'b11110000011001;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001010100001;
    x_1 = 'b00001111110110;
    x_2 = 'b00001101011001;
    x_3 = 'b00000100010101;

    h_0 = 'b00000010010001;
    h_1 = 'b00000110100110;
    h_2 = 'b00001010011010;
    h_3 = 'b00001101011001;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001111110101;
    x_1 = 'b11111011011001;
    x_2 = 'b11110001100001;
    x_3 = 'b00001000110101;

    h_0 = 'b11111010011001;
    h_1 = 'b11110001111011;
    h_2 = 'b11110000011001;
    h_3 = 'b11110110100010;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00000110100110;
    x_1 = 'b11110011111111;
    x_2 = 'b00001111010011;
    x_3 = 'b11110000001000;

    h_0 = 'b11110011111001;
    h_1 = 'b11110111011011;
    h_2 = 'b00001110100111;
    h_3 = 'b00000100010101;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110111010011;
    x_1 = 'b00001110100111;
    x_2 = 'b11110000001100;
    x_3 = 'b00001011111011;

    h_0 = 'b11110000010111;
    h_1 = 'b00001100110111;
    h_2 = 'b11111000001101;
    h_3 = 'b00000001010110;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110000000000;
    x_1 = 'b11111111110111;
    x_2 = 'b00010000000000;
    x_3 = 'b00000000010010;

    h_0 = 'b11110000101010;
    h_1 = 'b00001010011010;
    h_2 = 'b11111101111000;
    h_3 = 'b11111001001010;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110111011011;
    x_1 = 'b11110001100001;
    x_2 = 'b11110000001000;
    x_3 = 'b11110011101101;

    h_0 = 'b11110100101110;
    h_1 = 'b11110100100111;
    h_2 = 'b00001011001100;
    h_3 = 'b00001011011111;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00000110101110;
    x_1 = 'b00001100001101;
    x_2 = 'b00001111011011;
    x_3 = 'b00001111110010;

    h_0 = 'b11111011100010;
    h_1 = 'b11110011111111;
    h_2 = 'b11110000001100;
    h_3 = 'b11110001010101;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001111110110;
    x_1 = 'b00000100010101;
    x_2 = 'b11110001010101;
    x_3 = 'b11110111101010;

    h_0 = 'b00000011011100;
    h_1 = 'b00001001101100;
    h_2 = 'b00001110001001;
    h_3 = 'b00001111111111;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001010011010;
    x_1 = 'b11110000001100;
    x_2 = 'b00001101100111;
    x_3 = 'b11111011001000;

    h_0 = 'b00001010100001;
    h_1 = 'b00001101011001;
    h_2 = 'b11111001001010;
    h_3 = 'b11110000101111;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11111011011001;
    x_1 = 'b00001000110101;
    x_2 = 'b11110011101101;
    x_3 = 'b00001110101110;

    h_0 = 'b00001111000001;
    h_1 = 'b11111000001101;
    h_2 = 'b11111100110101;
    h_3 = 'b00001100100111;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110000101000;
    x_1 = 'b00001000011110;
    x_2 = 'b00001010101110;
    x_3 = 'b11110001101001;

    h_0 = 'b00001111110101;
    h_1 = 'b11110001100001;
    h_2 = 'b00001011111011;
    h_3 = 'b11110111101010;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110011111111;
    x_1 = 'b11110000001000;
    x_2 = 'b11110111000100;
    x_3 = 'b00000100000100;

    h_0 = 'b00001100110010;
    h_1 = 'b00000101110000;
    h_2 = 'b11110000000100;
    h_3 = 'b00000011000010;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00000010011001;
    x_1 = 'b00000100101111;
    x_2 = 'b00000110111111;
    x_3 = 'b00001001000100;

    h_0 = 'b00000110100110;
    h_1 = 'b00001111010011;
    h_2 = 'b00001101100111;
    h_3 = 'b00000010101011;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001110100111;
    x_1 = 'b00001011111011;
    x_2 = 'b11111011001000;
    x_3 = 'b11110000000110;

    h_0 = 'b11111110110011;
    h_1 = 'b11111100011011;
    h_2 = 'b11111010001000;
    h_3 = 'b11110111111101;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001101011001;
    x_1 = 'b11110001010101;
    x_2 = 'b00000010101011;
    x_3 = 'b00001011101111;

    h_0 = 'b11110111010011;
    h_1 = 'b11110000001100;
    h_2 = 'b11111011110011;
    h_3 = 'b00001100011000;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11111111110111;
    x_1 = 'b00000000010010;
    x_2 = 'b11111111100101;
    x_3 = 'b00000000100100;

    h_0 = 'b11110001111011;
    h_1 = 'b00000001010110;
    h_2 = 'b00001100100111;
    h_3 = 'b11110000110110;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110010011101;
    x_1 = 'b00001110011011;
    x_2 = 'b11111110001010;
    x_3 = 'b11110011100010;

    h_0 = 'b11110000000000;
    h_1 = 'b00010000000000;
    h_2 = 'b11110000000000;
    h_3 = 'b00010000000000;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110001100001;
    x_1 = 'b11110011101101;
    x_2 = 'b00000100000100;
    x_3 = 'b00001111101111;

    h_0 = 'b11110010000000;
    h_1 = 'b00000000111011;
    h_2 = 'b00001101000010;
    h_3 = 'b11110001001101;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11111101111000;
    x_1 = 'b11111011110011;
    x_2 = 'b11111001110011;
    x_3 = 'b11110111111001;

    h_0 = 'b11110111011011;
    h_1 = 'b11110000001000;
    h_2 = 'b11111011001000;
    h_3 = 'b00001011101111;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001100001101;
    x_1 = 'b00001111110010;
    x_2 = 'b00001000001110;
    x_3 = 'b11111010110111;

    h_0 = 'b11111110111100;
    h_1 = 'b11111100110101;
    h_2 = 'b11111010110010;
    h_3 = 'b11111000110101;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001111010011;
    x_1 = 'b11110111000100;
    x_2 = 'b11110101111011;
    x_3 = 'b00001110110101;

    h_0 = 'b00000110101110;
    h_1 = 'b00001111011011;
    h_2 = 'b00001101001111;
    h_3 = 'b00000001101101;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00000100010101;
    x_1 = 'b11110111101010;
    x_2 = 'b00001011101111;
    x_3 = 'b11110001110001;

    h_0 = 'b00001100110111;
    h_1 = 'b00000101010110;
    h_2 = 'b11110000000001;
    h_3 = 'b00000100000000;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110101011000;
    x_1 = 'b00001111111001;
    x_2 = 'b11110010110110;
    x_3 = 'b00000011110010;

    h_0 = 'b00001111110110;
    h_1 = 'b11110001010101;
    h_2 = 'b00001100011000;
    h_3 = 'b11110110110101;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110000001100;
    x_1 = 'b11111011001000;
    x_2 = 'b00001110010011;
    x_3 = 'b00001001010011;

    h_0 = 'b00001110111101;
    h_1 = 'b11111000100101;
    h_2 = 'b11111100001001;
    h_3 = 'b00001101001100;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11111001100010;
    x_1 = 'b11110100001011;
    x_2 = 'b11110000110101;
    x_3 = 'b11110000000100;

    h_0 = 'b00001010011010;
    h_1 = 'b00001101100111;
    h_2 = 'b11111001110011;
    h_3 = 'b11110000011110;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001000110101;
    x_1 = 'b00001110101110;
    x_2 = 'b00001111101111;
    x_3 = 'b00001011100010;

    h_0 = 'b00000011010011;
    h_1 = 'b00001001010110;
    h_2 = 'b00001101110011;
    h_3 = 'b00001111111001;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00010000000000;
    x_1 = 'b11111111100101;
    x_2 = 'b11110000000001;
    x_3 = 'b00000000110110;

    h_0 = 'b11111011011001;
    h_1 = 'b11110011101101;
    h_2 = 'b11110000000110;
    h_3 = 'b11110001110001;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001000011110;
    x_1 = 'b11110001101001;
    x_2 = 'b00001111111011;
    x_3 = 'b11110011010111;

    h_0 = 'b11110100100111;
    h_1 = 'b11110100111010;
    h_2 = 'b00001011101100;
    h_3 = 'b00001010110010;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11111001001010;
    x_1 = 'b00001100011000;
    x_2 = 'b11110000011110;
    x_3 = 'b00001111101100;

    h_0 = 'b11110000101000;
    h_1 = 'b00001010101110;
    h_2 = 'b11111101001100;
    h_3 = 'b11111010000100;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110000001000;
    x_1 = 'b00000100000100;
    x_2 = 'b00001110110101;
    x_3 = 'b11111000001001;

    h_0 = 'b11110000011001;
    h_1 = 'b00001100100111;
    h_2 = 'b11111000110101;
    h_3 = 'b00000000010111;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110101101101;
    x_1 = 'b11110000001111;
    x_2 = 'b11110010001011;
    x_3 = 'b11111010100110;

    h_0 = 'b11110011111111;
    h_1 = 'b11110111000100;
    h_2 = 'b00001110010011;
    h_3 = 'b00000101010010;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00000100101111;
    x_1 = 'b00001001000100;
    x_2 = 'b00001100100100;
    x_3 = 'b00001110111100;

    h_0 = 'b11111010100001;
    h_1 = 'b11110010001000;
    h_2 = 'b11110000010000;
    h_3 = 'b11110101110000;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001111011011;
    x_1 = 'b00001000001110;
    x_2 = 'b11110100111110;
    x_3 = 'b11110001111001;

    h_0 = 'b00000010011001;
    h_1 = 'b00000110111111;
    h_2 = 'b00001010111100;
    h_3 = 'b00001101111010;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001011111011;
    x_1 = 'b11110000000110;
    x_2 = 'b00001001010011;
    x_3 = 'b00000011100001;

    h_0 = 'b00001001101100;
    h_1 = 'b00001110110111;
    h_2 = 'b11111110001111;
    h_3 = 'b11110000001101;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11111101011110;
    x_1 = 'b00000101000001;
    x_2 = 'b11111000101001;
    x_3 = 'b00001001100001;

    h_0 = 'b00001110100111;
    h_1 = 'b11111011001000;
    h_2 = 'b11110111111001;
    h_3 = 'b00001111101100;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110001010101;
    x_1 = 'b00001011101111;
    x_2 = 'b00000101010010;
    x_3 = 'b11110000000011;

    h_0 = 'b00001111111101;
    h_1 = 'b11110000011101;
    h_2 = 'b00001110110000;
    h_3 = 'b11110010011011;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110010101100;
    x_1 = 'b11110001001110;
    x_2 = 'b11111100111010;
    x_3 = 'b00001011010110;

    h_0 = 'b00001101011001;
    h_1 = 'b00000010101011;
    h_2 = 'b11110000011110;
    h_3 = 'b00001001110000;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00000000010010;
    x_1 = 'b00000000100100;
    x_2 = 'b00000000110110;
    x_3 = 'b00000001001000;

    h_0 = 'b00000111100011;
    h_1 = 'b00001111111011;
    h_2 = 'b00001010001001;
    h_3 = 'b11111011010101;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001101100111;
    x_1 = 'b00001110010011;
    x_2 = 'b00000001011010;
    x_3 = 'b11110011001100;

    h_0 = 'b11111111110111;
    h_1 = 'b11111111100101;
    h_2 = 'b11111111010011;
    h_3 = 'b11111111000001;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001110011011;
    x_1 = 'b11110011100010;
    x_2 = 'b11111100010110;
    x_3 = 'b00001111101000;

    h_0 = 'b11111000001101;
    h_1 = 'b11110000000001;
    h_2 = 'b11110111000000;
    h_3 = 'b00000110100010;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00000001111111;
    x_1 = 'b11111100000101;
    x_2 = 'b00000101110100;
    x_3 = 'b11111000011001;

    h_0 = 'b11110010011101;
    h_1 = 'b11111110001010;
    h_2 = 'b00001111001000;
    h_3 = 'b11110100110001;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110011101101;
    x_1 = 'b00001111101111;
    x_2 = 'b11111000001001;
    x_3 = 'b11111010010101;

    h_0 = 'b11110000000010;
    h_1 = 'b00001111101110;
    h_2 = 'b11110000110001;
    h_3 = 'b00001110100001;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110000101111;
    x_1 = 'b11110110110101;
    x_2 = 'b00001001110000;
    x_3 = 'b00001111000010;

    h_0 = 'b11110001100001;
    h_1 = 'b00000100000100;
    h_2 = 'b00001001010011;
    h_3 = 'b11110000000011;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11111011110011;
    x_1 = 'b11110111111001;
    x_2 = 'b11110100100100;
    x_3 = 'b11110010000010;

    h_0 = 'b11110110100010;
    h_1 = 'b11110000110110;
    h_2 = 'b00000000010111;
    h_3 = 'b00001111010111;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001010101110;
    x_1 = 'b00001111111011;
    x_2 = 'b00001100111010;
    x_3 = 'b00000011001111;

    h_0 = 'b11111101111000;
    h_1 = 'b11111001110011;
    h_2 = 'b11110110001001;
    h_3 = 'b11110011001100;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001111110010;
    x_1 = 'b11111010110111;
    x_2 = 'b11110001111001;
    x_3 = 'b00001001110000;

    h_0 = 'b00000101110000;
    h_1 = 'b00001110010001;
    h_2 = 'b00001111011100;
    h_3 = 'b00001000101001;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00000110010101;
    x_1 = 'b11110100010111;
    x_2 = 'b00001111000010;
    x_3 = 'b11110000000010;

    h_0 = 'b00001100001101;
    h_1 = 'b00001000001110;
    h_2 = 'b11110001001000;
    h_3 = 'b11111100101000;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110111000100;
    x_1 = 'b00001110110101;
    x_2 = 'b11110000010110;
    x_3 = 'b00001011001001;

    h_0 = 'b00001111101011;
    h_1 = 'b11110010111001;
    h_2 = 'b00001000011010;
    h_3 = 'b11111101101011;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110000000000;
    x_1 = 'b11111111010011;
    x_2 = 'b00001111111110;
    x_3 = 'b00000001011011;

    h_0 = 'b00001111010011;
    h_1 = 'b11110101111011;
    h_2 = 'b00000001011010;
    h_3 = 'b00000111101111;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110111101010;
    x_1 = 'b11110001110001;
    x_2 = 'b11110000000011;
    x_3 = 'b11110011000001;

    h_0 = 'b00001011001100;
    h_1 = 'b00001011101100;
    h_2 = 'b11110101010101;
    h_3 = 'b11110011110110;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00000110111111;
    x_1 = 'b00001100100100;
    x_2 = 'b00001111101000;
    x_3 = 'b00001111100100;

    h_0 = 'b00000100010101;
    h_1 = 'b00001011101111;
    h_2 = 'b00001111101100;
    h_3 = 'b00001111000010;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001111111001;
    x_1 = 'b00000011110010;
    x_2 = 'b11110001000001;
    x_3 = 'b11111000101001;

    h_0 = 'b11111100011011;
    h_1 = 'b11110101111111;
    h_2 = 'b11110001100011;
    h_3 = 'b11110000000000;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001010001100;
    x_1 = 'b11110000010010;
    x_2 = 'b00001110000011;
    x_3 = 'b11111010000100;

    h_0 = 'b11110101011000;
    h_1 = 'b11110010110110;
    h_2 = 'b00000111011111;
    h_3 = 'b00001110111100;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11111011001000;
    x_1 = 'b00001001010011;
    x_2 = 'b11110011001100;
    x_3 = 'b00001111001000;

    h_0 = 'b11110000111100;
    h_1 = 'b00001000001010;
    h_2 = 'b00000010011110;
    h_3 = 'b11110100000010;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110000100011;
    x_1 = 'b00000111111111;
    x_2 = 'b00001011010110;
    x_3 = 'b11110010001011;

    h_0 = 'b11110000001100;
    h_1 = 'b00001110010011;
    h_2 = 'b11110100100100;
    h_3 = 'b00000111011111;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110100001011;
    x_1 = 'b11110000000100;
    x_2 = 'b11110110011000;
    x_3 = 'b00000010111101;

    h_0 = 'b11110011010100;
    h_1 = 'b11111001110111;
    h_2 = 'b00001111110111;
    h_3 = 'b11111101111101;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00000010101011;
    x_1 = 'b00000101010010;
    x_2 = 'b00000111101111;
    x_3 = 'b00001001111110;

    h_0 = 'b11111001100010;
    h_1 = 'b11110000110101;
    h_2 = 'b11110010000010;
    h_3 = 'b11111100010110;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001110101110;
    x_1 = 'b00001011100010;
    x_2 = 'b11111010010101;
    x_3 = 'b11110000000001;

    h_0 = 'b00000001010110;
    h_1 = 'b00000100000000;
    h_2 = 'b00000110100010;
    h_3 = 'b00001000111000;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001101001111;
    x_1 = 'b11110001001000;
    x_2 = 'b00000011100001;
    x_3 = 'b00001010111100;

    h_0 = 'b00001000110101;
    h_1 = 'b00001111101111;
    h_2 = 'b00000011100001;
    h_3 = 'b11110011000001;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11111111100101;
    x_1 = 'b00000000110110;
    x_2 = 'b11111110101111;
    x_3 = 'b00000001101101;

    h_0 = 'b00001110001001;
    h_1 = 'b11111110001111;
    h_2 = 'b11110011110110;
    h_3 = 'b00001111011100;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110010010100;
    x_1 = 'b00001110001011;
    x_2 = 'b11111111000001;
    x_3 = 'b11110010110110;

    h_0 = 'b00010000000000;
    h_1 = 'b11110000000001;
    h_2 = 'b00001111111110;
    h_3 = 'b11110000000100;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110001101001;
    x_1 = 'b11110011010111;
    x_2 = 'b00000011001111;
    x_3 = 'b00001111100000;

    h_0 = 'b00001101111100;
    h_1 = 'b11111111100000;
    h_2 = 'b11110010100101;
    h_3 = 'b00001110011001;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11111110001010;
    x_1 = 'b11111100010110;
    x_2 = 'b11111010100110;
    x_3 = 'b11111000111001;

    h_0 = 'b00001000011110;
    h_1 = 'b00001111111011;
    h_2 = 'b00000101100011;
    h_3 = 'b11110100111110;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001100011000;
    x_1 = 'b00001111101100;
    x_2 = 'b00000111011111;
    x_3 = 'b11111001110011;

    h_0 = 'b00000000111011;
    h_1 = 'b00000010110000;
    h_2 = 'b00000100100010;
    h_3 = 'b00000110010001;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001111001110;
    x_1 = 'b11110110100110;
    x_2 = 'b11110110100110;
    x_3 = 'b00001111001110;

    h_0 = 'b11111001001010;
    h_1 = 'b11110000011110;
    h_2 = 'b11110011001100;
    h_3 = 'b11111111010011;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00000100000100;
    x_1 = 'b11111000001001;
    x_2 = 'b00001011001001;
    x_3 = 'b11110010010100;

    h_0 = 'b11110011000100;
    h_1 = 'b11111011000100;
    h_2 = 'b00010000000000;
    h_3 = 'b11111011000100;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110101001011;
    x_1 = 'b00001111111100;
    x_2 = 'b11110011010111;
    x_3 = 'b00000010101011;

    h_0 = 'b11110000001000;
    h_1 = 'b00001110110101;
    h_2 = 'b11110011001100;
    h_3 = 'b00001001111110;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110000001111;
    x_1 = 'b11111010100110;
    x_2 = 'b00001101111010;
    x_3 = 'b00001010001100;

    h_0 = 'b11110001000110;
    h_1 = 'b00000111000011;
    h_2 = 'b00000100100010;
    h_3 = 'b11110010010010;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11111001110011;
    x_1 = 'b11110100100100;
    x_2 = 'b11110001001000;
    x_3 = 'b11110000000000;

    h_0 = 'b11110101101101;
    h_1 = 'b11110010001011;
    h_2 = 'b00000101100011;
    h_3 = 'b00001111101111;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001001000100;
    x_1 = 'b00001110111100;
    x_2 = 'b00001111100100;
    x_3 = 'b00001010101110;

    h_0 = 'b11111100110101;
    h_1 = 'b11110111000000;
    h_2 = 'b11110010100101;
    h_3 = 'b11110000010000;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00010000000000;
    x_1 = 'b11111111000001;
    x_2 = 'b11110000000100;
    x_3 = 'b00000001111111;

    h_0 = 'b00000100101111;
    h_1 = 'b00001100100100;
    h_2 = 'b00001111111110;
    h_3 = 'b00001101110001;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001000001110;
    x_1 = 'b11110001111001;
    x_2 = 'b00001111111111;
    x_3 = 'b11110010101100;

    h_0 = 'b00001011011111;
    h_1 = 'b00001010110010;
    h_2 = 'b11110011110110;
    h_3 = 'b11110101111111;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11111000111001;
    x_1 = 'b00001100101111;
    x_2 = 'b11110000010010;
    x_3 = 'b00001111011011;

    h_0 = 'b00001111011011;
    h_1 = 'b11110100111110;
    h_2 = 'b00000011100001;
    h_3 = 'b00000101000001;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110000000110;
    x_1 = 'b00000011100001;
    x_2 = 'b00001111001000;
    x_3 = 'b11111001001010;

    h_0 = 'b00001111100101;
    h_1 = 'b11110011101010;
    h_2 = 'b00000110100010;
    h_3 = 'b00000000101001;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110101111011;
    x_1 = 'b11110000010110;
    x_2 = 'b11110001110001;
    x_3 = 'b11111001100010;

    h_0 = 'b00001011111011;
    h_1 = 'b00001001010011;
    h_2 = 'b11110010000010;
    h_3 = 'b11111001110011;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00000101000001;
    x_1 = 'b00001001100001;
    x_2 = 'b00001101000100;
    x_3 = 'b00001111010011;

    h_0 = 'b00000101010110;
    h_1 = 'b00001101101010;
    h_2 = 'b00001111110111;
    h_3 = 'b00001010111111;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001111100000;
    x_1 = 'b00000111101111;
    x_2 = 'b11110100010111;
    x_3 = 'b11110010011101;

    h_0 = 'b11111101011110;
    h_1 = 'b11111000101001;
    h_2 = 'b11110100100100;
    h_3 = 'b11110001101001;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001011101111;
    x_1 = 'b11110000000011;
    x_2 = 'b00001001111110;
    x_3 = 'b00000010011001;

    h_0 = 'b11110110001101;
    h_1 = 'b11110001010100;
    h_2 = 'b00000010011110;
    h_3 = 'b00001111111011;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11111101001100;
    x_1 = 'b00000101100011;
    x_2 = 'b11110111111001;
    x_3 = 'b00001010011010;

    h_0 = 'b11110001010101;
    h_1 = 'b00000101010010;
    h_2 = 'b00000111011111;
    h_3 = 'b11110000100011;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110001001110;
    x_1 = 'b00001011010110;
    x_2 = 'b00000110000101;
    x_3 = 'b11110000000000;

    h_0 = 'b11110000000100;
    h_1 = 'b00001111011100;
    h_2 = 'b11110001100011;
    h_3 = 'b00001101000010;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110010110110;
    x_1 = 'b11110001000001;
    x_2 = 'b11111100000101;
    x_3 = 'b00001010100001;

    h_0 = 'b11110010101100;
    h_1 = 'b11111100111010;
    h_2 = 'b00001111101100;
    h_3 = 'b11110111000100;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00000000100100;
    x_1 = 'b00000001001000;
    x_2 = 'b00000001101101;
    x_3 = 'b00000010010001;

    h_0 = 'b11111000100101;
    h_1 = 'b11110000001000;
    h_2 = 'b11110101010101;
    h_3 = 'b00000011101110;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001101110001;
    x_1 = 'b00001110000011;
    x_2 = 'b00000000100100;
    x_3 = 'b11110010100010;

    h_0 = 'b00000000010010;
    h_1 = 'b00000000110110;
    h_2 = 'b00000001011011;
    h_3 = 'b00000001111111;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001110010011;
    x_1 = 'b11110011001100;
    x_2 = 'b11111101001100;
    x_3 = 'b00001111010110;

    h_0 = 'b00000111111011;
    h_1 = 'b00010000000000;
    h_2 = 'b00001000011010;
    h_3 = 'b11111000100101;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00000001101101;
    x_1 = 'b11111100101000;
    x_2 = 'b00000101000001;
    x_3 = 'b11111001011010;

    h_0 = 'b00001101100111;
    h_1 = 'b00000001011010;
    h_2 = 'b11110001001000;
    h_3 = 'b00001011111011;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110011100010;
    x_1 = 'b00001111101000;
    x_2 = 'b11111000111001;
    x_3 = 'b11111001010010;

    h_0 = 'b00001111111111;
    h_1 = 'b11110000001101;
    h_2 = 'b00001111011100;
    h_3 = 'b11110001000110;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110000110101;
    x_1 = 'b11110110011000;
    x_2 = 'b00001001000100;
    x_3 = 'b00001111011000;

    h_0 = 'b00001110011011;
    h_1 = 'b11111100010110;
    h_2 = 'b11110110001001;
    h_3 = 'b00010000000000;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11111100000101;
    x_1 = 'b11111000011001;
    x_2 = 'b11110101001011;
    x_3 = 'b11110010100111;

    h_0 = 'b00001001010110;
    h_1 = 'b00001111010010;
    h_2 = 'b00000000010111;
    h_3 = 'b11110000111100;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001010111100;
    x_1 = 'b00001111111110;
    x_2 = 'b00001100011000;
    x_3 = 'b00000010000111;

    h_0 = 'b00000001111111;
    h_1 = 'b00000101110100;
    h_2 = 'b00001001010011;
    h_3 = 'b00001100001101;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00001111101111;
    x_1 = 'b11111010010101;
    x_2 = 'b11110010010100;
    x_3 = 'b00001010101000;

    h_0 = 'b11111010001000;
    h_1 = 'b11110001100011;
    h_2 = 'b11110000110001;
    h_3 = 'b11111000001101;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00000110000101;
    x_1 = 'b11110100110001;
    x_2 = 'b00001110101110;
    x_3 = 'b11110000000000;

    h_0 = 'b11110011101101;
    h_1 = 'b11111000001001;
    h_2 = 'b00001111001000;
    h_3 = 'b00000010011001;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110110110101;
    x_1 = 'b00001111000010;
    x_2 = 'b11110000100011;
    x_3 = 'b00001010010011;

    h_0 = 'b11110000010011;
    h_1 = 'b00001101010110;
    h_2 = 'b11110111000000;
    h_3 = 'b00000011010011;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110000000001;
    x_1 = 'b11111110101111;
    x_2 = 'b00001111111001;
    x_3 = 'b00000010100010;

    h_0 = 'b11110000101111;
    h_1 = 'b00001001110000;
    h_2 = 'b11111111010011;
    h_3 = 'b11110111011011;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b11110111111001;
    x_1 = 'b11110010000010;
    x_2 = 'b11110000000000;
    x_3 = 'b11110010011001;

    h_0 = 'b11110100111010;
    h_1 = 'b11110100000010;
    h_2 = 'b00001010001001;
    h_3 = 'b00001100110010;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    x_0 = 'b00000111001111;
    x_1 = 'b00001100111010;
    x_2 = 'b00001111110010;
    x_3 = 'b00001111010001;

    h_0 = 'b11111011110011;
    h_1 = 'b11110100100100;
    h_2 = 'b11110000011110;
    h_3 = 'b11110000101010;
    #20;
    $fdisplay(fd, "%014b %014b %014b %014b", y_0, y_1, y_2, y_3);

    $fclose(fd);    
$finish;
    end
endmodule