`timescale 1ns / 1ps

module gru_tb;

// Parameters
parameter int D          = 64;
parameter int H          = 16;
parameter int DATA_WIDTH = 21;
parameter int FRAC_BITS  = 11;
parameter int NUM_PARALLEL = 1;
parameter real CLK_PERIOD = 10.0;

// Clock and reset
logic clk;
logic rst_n;
logic start;
logic done;

// Cycle counter
int cycle_count = 0;
int test_start_cycle = 0;
int test_cycles = 0;
int total_cycles = 0;
bit test_timeout = 0;

// Input arrays
logic signed [DATA_WIDTH-1:0] x_t [D-1:0];
logic signed [DATA_WIDTH-1:0] h_t_prev [H-1:0];
logic signed [DATA_WIDTH-1:0] h_t [H-1:0];

// Weight matrices
logic signed [DATA_WIDTH-1:0] W_ir [H-1:0][D-1:0];
logic signed [DATA_WIDTH-1:0] W_hr [H-1:0][H-1:0];
logic signed [DATA_WIDTH-1:0] b_ir [H-1:0];
logic signed [DATA_WIDTH-1:0] b_hr [H-1:0];

logic signed [DATA_WIDTH-1:0] W_iz [H-1:0][D-1:0];
logic signed [DATA_WIDTH-1:0] W_hz [H-1:0][H-1:0];
logic signed [DATA_WIDTH-1:0] b_iz [H-1:0];
logic signed [DATA_WIDTH-1:0] b_hz [H-1:0];

logic signed [DATA_WIDTH-1:0] W_in [H-1:0][D-1:0];
logic signed [DATA_WIDTH-1:0] W_hn [H-1:0][H-1:0];
logic signed [DATA_WIDTH-1:0] b_in [H-1:0];
logic signed [DATA_WIDTH-1:0] b_hn [H-1:0];

// DUT instantiation
gru_cell_parallel #(
    .D(D),
    .H(H),
    .DATA_WIDTH(DATA_WIDTH),
    .FRAC_BITS(FRAC_BITS),
    .NUM_PARALLEL(NUM_PARALLEL)
) dut (
    .clk(clk),
    .rst_n(rst_n),
    .start(start),
    .x_t(x_t),
    .h_t_prev(h_t_prev),
    .W_ir(W_ir),
    .W_hr(W_hr),
    .b_ir(b_ir),
    .b_hr(b_hr),
    .W_iz(W_iz),
    .W_hz(W_hz),
    .b_iz(b_iz),
    .b_hz(b_hz),
    .W_in(W_in),
    .W_hn(W_hn),
    .b_in(b_in),
    .b_hn(b_hn),
    .h_t(h_t),
    .done(done)
);

// Clock generation
initial begin
    clk = 0;
    forever #5 clk = ~clk; // 100MHz clock
end

// Cycle counter
always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        cycle_count <= 0;
    end else begin
        cycle_count <= cycle_count + 1;
    end
end

initial begin
    // Open files for writing
    integer fd_output;
    integer fd_cycles;
    
    fd_output = $fopen("../../../../../output_d64_h16_dw21_fb11_np1.txt", "w+");
    if (fd_output == 0) begin
        $display("ERROR: Failed to open output file!");
        $finish;
    end
    
    fd_cycles = $fopen("../../../../../cycles_d64_h16_dw21_fb11_np1.txt", "w+");
    if (fd_cycles == 0) begin
        $display("ERROR: Failed to open cycles file!");
        $fclose(fd_output);
        $finish;
    end
    
    // Write header to cycles file
    $fdisplay(fd_cycles, "==========================================================");
    $fdisplay(fd_cycles, "GRU Cell Parallel Cycle Count Results");
    $fdisplay(fd_cycles, "==========================================================");
    $fdisplay(fd_cycles, "Parameters:");
    $fdisplay(fd_cycles, "  D (Input Dimension):     64");
    $fdisplay(fd_cycles, "  H (Hidden Dimension):    16");
    $fdisplay(fd_cycles, "  DATA_WIDTH:              21");
    $fdisplay(fd_cycles, "  FRAC_BITS:               11");
    $fdisplay(fd_cycles, "  NUM_PARALLEL:            1");
    $fdisplay(fd_cycles, "  Total Test Vectors:      100");
    $fdisplay(fd_cycles, "==========================================================");
    $fdisplay(fd_cycles, "");
    
    // Initialize weights
    // Initialize W_ir weights
    W_ir[0][0] = 21'b000000000000010100101;
    W_ir[0][1] = 21'b000000000000100111001;
    W_ir[0][2] = 21'b000000000000011101110;
    W_ir[0][3] = 21'b000000000000100011010;
    W_ir[0][4] = 21'b111111111111101101010;
    W_ir[0][5] = 21'b111111111111010101010;
    W_ir[0][6] = 21'b000000000000011100111;
    W_ir[0][7] = 21'b000000000000001111011;
    W_ir[0][8] = 21'b111111111111001000001;
    W_ir[0][9] = 21'b000000000000000101101;
    W_ir[0][10] = 21'b000000000000111110110;
    W_ir[0][11] = 21'b111111111111111111101;
    W_ir[0][12] = 21'b000000000000101000000;
    W_ir[0][13] = 21'b000000000000001011000;
    W_ir[0][14] = 21'b000000000000001001111;
    W_ir[0][15] = 21'b000000000000101110011;
    W_ir[0][16] = 21'b111111111111111000000;
    W_ir[0][17] = 21'b000000000000110111010;
    W_ir[0][18] = 21'b111111111111111000110;
    W_ir[0][19] = 21'b000000000000100100010;
    W_ir[0][20] = 21'b111111111111111000100;
    W_ir[0][21] = 21'b000000000000100001110;
    W_ir[0][22] = 21'b000000000000011000100;
    W_ir[0][23] = 21'b000000000000011000111;
    W_ir[0][24] = 21'b111111111111010111110;
    W_ir[0][25] = 21'b000000000000011110000;
    W_ir[0][26] = 21'b000000000000100010111;
    W_ir[0][27] = 21'b000000000000010110111;
    W_ir[0][28] = 21'b000000000000111000101;
    W_ir[0][29] = 21'b111111111111001011000;
    W_ir[0][30] = 21'b111111111111101101011;
    W_ir[0][31] = 21'b000000000000011001110;
    W_ir[0][32] = 21'b000000000000001100011;
    W_ir[0][33] = 21'b000000000000011110100;
    W_ir[0][34] = 21'b000000000000011110101;
    W_ir[0][35] = 21'b000000000000000110110;
    W_ir[0][36] = 21'b000000000000111111101;
    W_ir[0][37] = 21'b000000000000010100010;
    W_ir[0][38] = 21'b111111111111101110110;
    W_ir[0][39] = 21'b000000000000001111011;
    W_ir[0][40] = 21'b000000000000100101011;
    W_ir[0][41] = 21'b111111111111010000010;
    W_ir[0][42] = 21'b000000000000001111010;
    W_ir[0][43] = 21'b111111111111101000010;
    W_ir[0][44] = 21'b111111111111111110010;
    W_ir[0][45] = 21'b111111111111011100101;
    W_ir[0][46] = 21'b111111111111001110100;
    W_ir[0][47] = 21'b000000000000110111101;
    W_ir[0][48] = 21'b111111111111110001010;
    W_ir[0][49] = 21'b111111111111100111001;
    W_ir[0][50] = 21'b111111111111111001101;
    W_ir[0][51] = 21'b000000000000000000010;
    W_ir[0][52] = 21'b111111111111000110110;
    W_ir[0][53] = 21'b111111111111101010010;
    W_ir[0][54] = 21'b000000000000010000110;
    W_ir[0][55] = 21'b111111111111100111110;
    W_ir[0][56] = 21'b000000000000100110010;
    W_ir[0][57] = 21'b111111111111100101011;
    W_ir[0][58] = 21'b111111111111101011011;
    W_ir[0][59] = 21'b000000000000100010000;
    W_ir[0][60] = 21'b111111111111010101000;
    W_ir[0][61] = 21'b111111111111001101111;
    W_ir[0][62] = 21'b111111111111001100100;
    W_ir[0][63] = 21'b000000000000100001100;
    W_ir[1][0] = 21'b111111111111100010111;
    W_ir[1][1] = 21'b111111111111100110011;
    W_ir[1][2] = 21'b000000000000101111111;
    W_ir[1][3] = 21'b000000000000100101101;
    W_ir[1][4] = 21'b000000000000000101001;
    W_ir[1][5] = 21'b000000000000001111100;
    W_ir[1][6] = 21'b000000000000001101001;
    W_ir[1][7] = 21'b000000000000001000010;
    W_ir[1][8] = 21'b000000000000001010000;
    W_ir[1][9] = 21'b000000000000001001010;
    W_ir[1][10] = 21'b111111111111111000100;
    W_ir[1][11] = 21'b111111111111111111110;
    W_ir[1][12] = 21'b000000000000001011101;
    W_ir[1][13] = 21'b000000000000011100000;
    W_ir[1][14] = 21'b111111111111010101101;
    W_ir[1][15] = 21'b000000000000001000100;
    W_ir[1][16] = 21'b111111111111111111111;
    W_ir[1][17] = 21'b111111111111111111001;
    W_ir[1][18] = 21'b111111111111111100100;
    W_ir[1][19] = 21'b111111111111101100000;
    W_ir[1][20] = 21'b111111111111111100000;
    W_ir[1][21] = 21'b000000000000001011011;
    W_ir[1][22] = 21'b111111111111110000000;
    W_ir[1][23] = 21'b111111111111101000000;
    W_ir[1][24] = 21'b000000000000000000011;
    W_ir[1][25] = 21'b000000000000101110101;
    W_ir[1][26] = 21'b111111111111001100101;
    W_ir[1][27] = 21'b111111111111001110101;
    W_ir[1][28] = 21'b000000000000110101101;
    W_ir[1][29] = 21'b000000000000010000010;
    W_ir[1][30] = 21'b000000000000000011101;
    W_ir[1][31] = 21'b111111111111111111011;
    W_ir[1][32] = 21'b111111111111100001010;
    W_ir[1][33] = 21'b111111111111111101001;
    W_ir[1][34] = 21'b111111111111111011010;
    W_ir[1][35] = 21'b000000000000000011110;
    W_ir[1][36] = 21'b000000000000001111110;
    W_ir[1][37] = 21'b000000000000001001001;
    W_ir[1][38] = 21'b000000000000001100101;
    W_ir[1][39] = 21'b000000000000100000001;
    W_ir[1][40] = 21'b000000000000010011010;
    W_ir[1][41] = 21'b000000000000000000011;
    W_ir[1][42] = 21'b111111111111111101010;
    W_ir[1][43] = 21'b000000000000010000010;
    W_ir[1][44] = 21'b000000000000000110001;
    W_ir[1][45] = 21'b000000000000001100101;
    W_ir[1][46] = 21'b111111111111111100111;
    W_ir[1][47] = 21'b111111111111110111001;
    W_ir[1][48] = 21'b111111111111110110111;
    W_ir[1][49] = 21'b111111111111001010111;
    W_ir[1][50] = 21'b000000000000011110101;
    W_ir[1][51] = 21'b000000000000101010101;
    W_ir[1][52] = 21'b111111111111110011100;
    W_ir[1][53] = 21'b111111111111100111011;
    W_ir[1][54] = 21'b111111111111101000000;
    W_ir[1][55] = 21'b111111111111100100111;
    W_ir[1][56] = 21'b111111111111110000011;
    W_ir[1][57] = 21'b000000000000110010111;
    W_ir[1][58] = 21'b000000000000011101110;
    W_ir[1][59] = 21'b111111111111011111001;
    W_ir[1][60] = 21'b111111111111110111101;
    W_ir[1][61] = 21'b111111111111110010011;
    W_ir[1][62] = 21'b000000000000101011000;
    W_ir[1][63] = 21'b111111111111100111110;
    W_ir[2][0] = 21'b111111111111101001001;
    W_ir[2][1] = 21'b111111111111110000001;
    W_ir[2][2] = 21'b111111111111001001100;
    W_ir[2][3] = 21'b111111111111011110010;
    W_ir[2][4] = 21'b111111111111101101011;
    W_ir[2][5] = 21'b111111111111110111011;
    W_ir[2][6] = 21'b000000000000000101111;
    W_ir[2][7] = 21'b111111111111010111011;
    W_ir[2][8] = 21'b111111111111110101000;
    W_ir[2][9] = 21'b111111111111110101100;
    W_ir[2][10] = 21'b111111111111110100001;
    W_ir[2][11] = 21'b111111111111000101101;
    W_ir[2][12] = 21'b111111111111110110110;
    W_ir[2][13] = 21'b000000000000001101111;
    W_ir[2][14] = 21'b111111111111110101000;
    W_ir[2][15] = 21'b000000000000010110000;
    W_ir[2][16] = 21'b111111111111010110100;
    W_ir[2][17] = 21'b000000000000111001011;
    W_ir[2][18] = 21'b000000000000000011000;
    W_ir[2][19] = 21'b000000000000010011000;
    W_ir[2][20] = 21'b000000000000001101111;
    W_ir[2][21] = 21'b111111111111101110000;
    W_ir[2][22] = 21'b000000000000011110000;
    W_ir[2][23] = 21'b000000000000110101000;
    W_ir[2][24] = 21'b000000000000011011000;
    W_ir[2][25] = 21'b000000000000001000111;
    W_ir[2][26] = 21'b111111111111111100000;
    W_ir[2][27] = 21'b111111111111001011011;
    W_ir[2][28] = 21'b111111111111110001000;
    W_ir[2][29] = 21'b000000000000111100011;
    W_ir[2][30] = 21'b111111111111101000000;
    W_ir[2][31] = 21'b111111111111101000010;
    W_ir[2][32] = 21'b000000000000000010110;
    W_ir[2][33] = 21'b000000000000010111000;
    W_ir[2][34] = 21'b111111111111110100010;
    W_ir[2][35] = 21'b111111111111110010100;
    W_ir[2][36] = 21'b000000000000000011000;
    W_ir[2][37] = 21'b000000000000001010101;
    W_ir[2][38] = 21'b000000000000100000000;
    W_ir[2][39] = 21'b111111111111111111101;
    W_ir[2][40] = 21'b000000000000011100100;
    W_ir[2][41] = 21'b111111111111110010101;
    W_ir[2][42] = 21'b000000000000011101101;
    W_ir[2][43] = 21'b111111111111111100110;
    W_ir[2][44] = 21'b000000000000001011010;
    W_ir[2][45] = 21'b000000000000001111111;
    W_ir[2][46] = 21'b000000000000001100100;
    W_ir[2][47] = 21'b000000000000000110100;
    W_ir[2][48] = 21'b000000000000001100111;
    W_ir[2][49] = 21'b000000000000001010111;
    W_ir[2][50] = 21'b111111111111100001100;
    W_ir[2][51] = 21'b000000000000010101110;
    W_ir[2][52] = 21'b000000000000010100100;
    W_ir[2][53] = 21'b000000000000001110010;
    W_ir[2][54] = 21'b111111111111001001010;
    W_ir[2][55] = 21'b000000000000010010110;
    W_ir[2][56] = 21'b000000000000001100100;
    W_ir[2][57] = 21'b111111111111010111010;
    W_ir[2][58] = 21'b111111111111100001111;
    W_ir[2][59] = 21'b111111111111100101101;
    W_ir[2][60] = 21'b000000000000100110011;
    W_ir[2][61] = 21'b000000000000010001100;
    W_ir[2][62] = 21'b000000000000100111110;
    W_ir[2][63] = 21'b000000000001000110101;
    W_ir[3][0] = 21'b111111111111111101111;
    W_ir[3][1] = 21'b000000000000111111011;
    W_ir[3][2] = 21'b000000000000000000001;
    W_ir[3][3] = 21'b000000000000110010101;
    W_ir[3][4] = 21'b111111111111010010000;
    W_ir[3][5] = 21'b000000000000001010011;
    W_ir[3][6] = 21'b000000000000000111101;
    W_ir[3][7] = 21'b111111111111101100111;
    W_ir[3][8] = 21'b111111111111111000110;
    W_ir[3][9] = 21'b000000000000101001101;
    W_ir[3][10] = 21'b111111111111100010011;
    W_ir[3][11] = 21'b111111111111111010100;
    W_ir[3][12] = 21'b111111111111011111101;
    W_ir[3][13] = 21'b111111111111110101001;
    W_ir[3][14] = 21'b111111111111110001111;
    W_ir[3][15] = 21'b111111111111111000110;
    W_ir[3][16] = 21'b000000000000000010011;
    W_ir[3][17] = 21'b000000000000001010110;
    W_ir[3][18] = 21'b111111111111101001110;
    W_ir[3][19] = 21'b000000000000100000100;
    W_ir[3][20] = 21'b111111111111110011000;
    W_ir[3][21] = 21'b000000000000001100111;
    W_ir[3][22] = 21'b000000000000010101001;
    W_ir[3][23] = 21'b000000000000001101101;
    W_ir[3][24] = 21'b000000000000110101001;
    W_ir[3][25] = 21'b000000000000001011101;
    W_ir[3][26] = 21'b111111111111111000100;
    W_ir[3][27] = 21'b111111111111101100101;
    W_ir[3][28] = 21'b000000000000001011011;
    W_ir[3][29] = 21'b000000000000001001100;
    W_ir[3][30] = 21'b111111111111011110000;
    W_ir[3][31] = 21'b000000000001000010010;
    W_ir[3][32] = 21'b000000000000100010000;
    W_ir[3][33] = 21'b111111111111011000101;
    W_ir[3][34] = 21'b000000000000010000000;
    W_ir[3][35] = 21'b000000000000001001010;
    W_ir[3][36] = 21'b000000000000001011110;
    W_ir[3][37] = 21'b111111111111000111111;
    W_ir[3][38] = 21'b000000000000011000100;
    W_ir[3][39] = 21'b000000000000000011101;
    W_ir[3][40] = 21'b111111111111111110111;
    W_ir[3][41] = 21'b000000000000100101011;
    W_ir[3][42] = 21'b111111111111010110010;
    W_ir[3][43] = 21'b000000000000000110000;
    W_ir[3][44] = 21'b111111111111101010000;
    W_ir[3][45] = 21'b111111111111101110001;
    W_ir[3][46] = 21'b000000000000110001100;
    W_ir[3][47] = 21'b111111111111101000111;
    W_ir[3][48] = 21'b111111111111110010100;
    W_ir[3][49] = 21'b111111111111110110011;
    W_ir[3][50] = 21'b111111111111100100000;
    W_ir[3][51] = 21'b111111111111101000001;
    W_ir[3][52] = 21'b111111111111100101111;
    W_ir[3][53] = 21'b111111111111100010111;
    W_ir[3][54] = 21'b111111111111101111011;
    W_ir[3][55] = 21'b111111111111000110000;
    W_ir[3][56] = 21'b111111111111100100110;
    W_ir[3][57] = 21'b000000000000011111010;
    W_ir[3][58] = 21'b111111111111011100111;
    W_ir[3][59] = 21'b111111111111100111001;
    W_ir[3][60] = 21'b111111111111101000000;
    W_ir[3][61] = 21'b111111111111101011011;
    W_ir[3][62] = 21'b111111111111010000010;
    W_ir[3][63] = 21'b111111111111101100000;
    W_ir[4][0] = 21'b111111111111111100100;
    W_ir[4][1] = 21'b111111111111110011011;
    W_ir[4][2] = 21'b111111111111110110110;
    W_ir[4][3] = 21'b111111111111100111010;
    W_ir[4][4] = 21'b000000000000000001010;
    W_ir[4][5] = 21'b000000000000010111001;
    W_ir[4][6] = 21'b111111111111100011011;
    W_ir[4][7] = 21'b111111111111010111010;
    W_ir[4][8] = 21'b111111111111000101000;
    W_ir[4][9] = 21'b111111111111101001011;
    W_ir[4][10] = 21'b111111111111001011100;
    W_ir[4][11] = 21'b111111111111101111000;
    W_ir[4][12] = 21'b111111111111110110101;
    W_ir[4][13] = 21'b000000000000010111000;
    W_ir[4][14] = 21'b000000000000000110010;
    W_ir[4][15] = 21'b111111111111110110101;
    W_ir[4][16] = 21'b111111111111100000110;
    W_ir[4][17] = 21'b111111111111101000101;
    W_ir[4][18] = 21'b111111111111100001101;
    W_ir[4][19] = 21'b111111111111011010101;
    W_ir[4][20] = 21'b111111111111110111001;
    W_ir[4][21] = 21'b000000000000011010110;
    W_ir[4][22] = 21'b000000000001000011110;
    W_ir[4][23] = 21'b000000000000100101100;
    W_ir[4][24] = 21'b111111111111001000001;
    W_ir[4][25] = 21'b111111111111010010111;
    W_ir[4][26] = 21'b000000000000000011101;
    W_ir[4][27] = 21'b111111111111001000001;
    W_ir[4][28] = 21'b000000000000101111101;
    W_ir[4][29] = 21'b111111111111111101101;
    W_ir[4][30] = 21'b000000000000101101100;
    W_ir[4][31] = 21'b111111111111100001001;
    W_ir[4][32] = 21'b111111111111001100000;
    W_ir[4][33] = 21'b111111111111010010101;
    W_ir[4][34] = 21'b111111111111100001100;
    W_ir[4][35] = 21'b111111111111011110111;
    W_ir[4][36] = 21'b111111111111001101101;
    W_ir[4][37] = 21'b111111111111010101011;
    W_ir[4][38] = 21'b111111111111100100100;
    W_ir[4][39] = 21'b000000000000010001010;
    W_ir[4][40] = 21'b000000000000001100000;
    W_ir[4][41] = 21'b111111111111100011001;
    W_ir[4][42] = 21'b111111111111111011111;
    W_ir[4][43] = 21'b111111111111101001111;
    W_ir[4][44] = 21'b111111111111000010010;
    W_ir[4][45] = 21'b111111111111110101100;
    W_ir[4][46] = 21'b111111111111110101010;
    W_ir[4][47] = 21'b111111111111111000011;
    W_ir[4][48] = 21'b000000000000000000001;
    W_ir[4][49] = 21'b111111111111110010100;
    W_ir[4][50] = 21'b000000000000101001110;
    W_ir[4][51] = 21'b111111111111100111000;
    W_ir[4][52] = 21'b000000000000111010100;
    W_ir[4][53] = 21'b000000000000011100010;
    W_ir[4][54] = 21'b000000000000111101100;
    W_ir[4][55] = 21'b000000000000110011011;
    W_ir[4][56] = 21'b000000000000010100001;
    W_ir[4][57] = 21'b111111111111001000100;
    W_ir[4][58] = 21'b000000000000100000111;
    W_ir[4][59] = 21'b000000000001101110110;
    W_ir[4][60] = 21'b000000000001010010110;
    W_ir[4][61] = 21'b000000000001010111011;
    W_ir[4][62] = 21'b000000000001100111001;
    W_ir[4][63] = 21'b000000000001011100000;
    W_ir[5][0] = 21'b000000000000001010100;
    W_ir[5][1] = 21'b000000000000001011011;
    W_ir[5][2] = 21'b000000000000001101011;
    W_ir[5][3] = 21'b111111111111111000010;
    W_ir[5][4] = 21'b111111111111110111011;
    W_ir[5][5] = 21'b111111111111011011000;
    W_ir[5][6] = 21'b000000000000110001111;
    W_ir[5][7] = 21'b111111111111000101010;
    W_ir[5][8] = 21'b111111111111010010100;
    W_ir[5][9] = 21'b111111111111101111011;
    W_ir[5][10] = 21'b111111111111111110101;
    W_ir[5][11] = 21'b111111111111110110101;
    W_ir[5][12] = 21'b111111111111011100001;
    W_ir[5][13] = 21'b111111111111110101100;
    W_ir[5][14] = 21'b111111111111100001000;
    W_ir[5][15] = 21'b111111111111011111111;
    W_ir[5][16] = 21'b000000000000100101000;
    W_ir[5][17] = 21'b111111111111010111110;
    W_ir[5][18] = 21'b000000000000000111110;
    W_ir[5][19] = 21'b111111111111001101111;
    W_ir[5][20] = 21'b111111111111110110000;
    W_ir[5][21] = 21'b000000000000000001011;
    W_ir[5][22] = 21'b000000000000010100101;
    W_ir[5][23] = 21'b000000000000001100111;
    W_ir[5][24] = 21'b111111111111111011000;
    W_ir[5][25] = 21'b111111111111100111101;
    W_ir[5][26] = 21'b111111111111111011010;
    W_ir[5][27] = 21'b000000000000010111010;
    W_ir[5][28] = 21'b000000000000000101000;
    W_ir[5][29] = 21'b111111111111100010100;
    W_ir[5][30] = 21'b111111111111110001000;
    W_ir[5][31] = 21'b111111111111001000100;
    W_ir[5][32] = 21'b111111111111111100011;
    W_ir[5][33] = 21'b111111111111000000001;
    W_ir[5][34] = 21'b111111111111101111111;
    W_ir[5][35] = 21'b000000000000011111001;
    W_ir[5][36] = 21'b111111111111100000100;
    W_ir[5][37] = 21'b111111111111010001001;
    W_ir[5][38] = 21'b111111111110111010011;
    W_ir[5][39] = 21'b000000000000101000111;
    W_ir[5][40] = 21'b111111111111101011101;
    W_ir[5][41] = 21'b111111111111111000000;
    W_ir[5][42] = 21'b000000000000000011011;
    W_ir[5][43] = 21'b111111111111101001100;
    W_ir[5][44] = 21'b000000000000001000010;
    W_ir[5][45] = 21'b111111111111101010100;
    W_ir[5][46] = 21'b111111111111110110110;
    W_ir[5][47] = 21'b000000000000011110100;
    W_ir[5][48] = 21'b000000000000001111010;
    W_ir[5][49] = 21'b000000000000001100100;
    W_ir[5][50] = 21'b000000000000001010101;
    W_ir[5][51] = 21'b000000000000001011001;
    W_ir[5][52] = 21'b111111111111101110110;
    W_ir[5][53] = 21'b111111111111101011100;
    W_ir[5][54] = 21'b000000000000001110101;
    W_ir[5][55] = 21'b000000000000000000001;
    W_ir[5][56] = 21'b000000000000001011000;
    W_ir[5][57] = 21'b111111111111011011111;
    W_ir[5][58] = 21'b111111111111011110011;
    W_ir[5][59] = 21'b111111111111101101100;
    W_ir[5][60] = 21'b000000000000111011101;
    W_ir[5][61] = 21'b000000000000101000100;
    W_ir[5][62] = 21'b111111111111101100000;
    W_ir[5][63] = 21'b000000000000100100010;
    W_ir[6][0] = 21'b000000000000101110101;
    W_ir[6][1] = 21'b111111111111110011101;
    W_ir[6][2] = 21'b000000000001001010111;
    W_ir[6][3] = 21'b111111111111101100111;
    W_ir[6][4] = 21'b000000000000101010000;
    W_ir[6][5] = 21'b000000000000001001111;
    W_ir[6][6] = 21'b111111111111001011000;
    W_ir[6][7] = 21'b000000000001001011000;
    W_ir[6][8] = 21'b000000000001010110010;
    W_ir[6][9] = 21'b000000000000110010101;
    W_ir[6][10] = 21'b000000000000111101101;
    W_ir[6][11] = 21'b111111111111111110100;
    W_ir[6][12] = 21'b000000000000000000111;
    W_ir[6][13] = 21'b000000000000010010101;
    W_ir[6][14] = 21'b111111111111101110000;
    W_ir[6][15] = 21'b111111111111001011100;
    W_ir[6][16] = 21'b111111111111101010010;
    W_ir[6][17] = 21'b000000000000100111011;
    W_ir[6][18] = 21'b111111111111111110101;
    W_ir[6][19] = 21'b111111111111111101001;
    W_ir[6][20] = 21'b111111111111110100011;
    W_ir[6][21] = 21'b111111111111010101011;
    W_ir[6][22] = 21'b000000000001000101100;
    W_ir[6][23] = 21'b111111111111111101100;
    W_ir[6][24] = 21'b111111111111010111010;
    W_ir[6][25] = 21'b000000000000010100001;
    W_ir[6][26] = 21'b111111111111010011110;
    W_ir[6][27] = 21'b111111111111011110000;
    W_ir[6][28] = 21'b000000000000110000111;
    W_ir[6][29] = 21'b000000000000101010010;
    W_ir[6][30] = 21'b111111111111010110000;
    W_ir[6][31] = 21'b000000000000100110100;
    W_ir[6][32] = 21'b000000000000000011011;
    W_ir[6][33] = 21'b000000000000010100010;
    W_ir[6][34] = 21'b000000000000110101101;
    W_ir[6][35] = 21'b000000000001000000010;
    W_ir[6][36] = 21'b111111111111111011001;
    W_ir[6][37] = 21'b000000000000001111101;
    W_ir[6][38] = 21'b111111111111000001011;
    W_ir[6][39] = 21'b111111111111111001101;
    W_ir[6][40] = 21'b000000000000011111111;
    W_ir[6][41] = 21'b111111111111100111100;
    W_ir[6][42] = 21'b000000000001000111000;
    W_ir[6][43] = 21'b000000000000010001000;
    W_ir[6][44] = 21'b000000000000100010001;
    W_ir[6][45] = 21'b111111111111100010100;
    W_ir[6][46] = 21'b111111111111001011101;
    W_ir[6][47] = 21'b000000000000111111111;
    W_ir[6][48] = 21'b111111111111010000001;
    W_ir[6][49] = 21'b111111111111100010010;
    W_ir[6][50] = 21'b000000000000100000010;
    W_ir[6][51] = 21'b111111111111111011011;
    W_ir[6][52] = 21'b000000000000100010000;
    W_ir[6][53] = 21'b111111111110010011000;
    W_ir[6][54] = 21'b111111111111110001011;
    W_ir[6][55] = 21'b000000000000001001101;
    W_ir[6][56] = 21'b111111111111011001011;
    W_ir[6][57] = 21'b111111111111101110001;
    W_ir[6][58] = 21'b111111111111010111000;
    W_ir[6][59] = 21'b111111111111010000100;
    W_ir[6][60] = 21'b111111111111110001011;
    W_ir[6][61] = 21'b111111111110011110000;
    W_ir[6][62] = 21'b111111111110001010000;
    W_ir[6][63] = 21'b111111111110000011000;
    W_ir[7][0] = 21'b111111111110101001010;
    W_ir[7][1] = 21'b111111111110100110001;
    W_ir[7][2] = 21'b000000000000011000111;
    W_ir[7][3] = 21'b111111111111110011001;
    W_ir[7][4] = 21'b000000000000110001101;
    W_ir[7][5] = 21'b000000000001000011110;
    W_ir[7][6] = 21'b111111111111001001011;
    W_ir[7][7] = 21'b000000000000001101000;
    W_ir[7][8] = 21'b111111111111010111011;
    W_ir[7][9] = 21'b111111111110011100101;
    W_ir[7][10] = 21'b111111111111011101111;
    W_ir[7][11] = 21'b000000000000100111101;
    W_ir[7][12] = 21'b000000000000101111110;
    W_ir[7][13] = 21'b111111111111010011011;
    W_ir[7][14] = 21'b000000000000110000100;
    W_ir[7][15] = 21'b111111111111111111111;
    W_ir[7][16] = 21'b000000000000001001111;
    W_ir[7][17] = 21'b111111111111101000000;
    W_ir[7][18] = 21'b000000000000001001110;
    W_ir[7][19] = 21'b000000000000111010110;
    W_ir[7][20] = 21'b111111111111100011111;
    W_ir[7][21] = 21'b111111111111101000101;
    W_ir[7][22] = 21'b000000000000111111011;
    W_ir[7][23] = 21'b111111111111100101010;
    W_ir[7][24] = 21'b000000000000111001000;
    W_ir[7][25] = 21'b000000000000011011100;
    W_ir[7][26] = 21'b000000000000100010101;
    W_ir[7][27] = 21'b111111111111110001110;
    W_ir[7][28] = 21'b000000000000101101010;
    W_ir[7][29] = 21'b000000000001000100010;
    W_ir[7][30] = 21'b000000000000101100101;
    W_ir[7][31] = 21'b000000000000011000000;
    W_ir[7][32] = 21'b111111111111010111010;
    W_ir[7][33] = 21'b111111111111100111011;
    W_ir[7][34] = 21'b111111111110100011110;
    W_ir[7][35] = 21'b111111111111001101001;
    W_ir[7][36] = 21'b000000000000111100101;
    W_ir[7][37] = 21'b000000000000000000100;
    W_ir[7][38] = 21'b000000000000110011010;
    W_ir[7][39] = 21'b111111111110111011111;
    W_ir[7][40] = 21'b111111111111111101110;
    W_ir[7][41] = 21'b111111111110111110000;
    W_ir[7][42] = 21'b111111111110111001101;
    W_ir[7][43] = 21'b111111111110110111000;
    W_ir[7][44] = 21'b111111111111011010100;
    W_ir[7][45] = 21'b000000000000001001101;
    W_ir[7][46] = 21'b000000000010001100001;
    W_ir[7][47] = 21'b111111111111011010011;
    W_ir[7][48] = 21'b111111111111111001110;
    W_ir[7][49] = 21'b111111111111010110100;
    W_ir[7][50] = 21'b111111111111000010100;
    W_ir[7][51] = 21'b000000000001011101100;
    W_ir[7][52] = 21'b111111111110111010011;
    W_ir[7][53] = 21'b000000000000010110001;
    W_ir[7][54] = 21'b000000000001000111000;
    W_ir[7][55] = 21'b000000000000001011010;
    W_ir[7][56] = 21'b000000000010010001011;
    W_ir[7][57] = 21'b000000000000010010011;
    W_ir[7][58] = 21'b000000000010010100011;
    W_ir[7][59] = 21'b000000000000010111101;
    W_ir[7][60] = 21'b111111111111000010100;
    W_ir[7][61] = 21'b000000000001000111000;
    W_ir[7][62] = 21'b000000000001100000011;
    W_ir[7][63] = 21'b111111111111000010100;
    W_ir[8][0] = 21'b111111111111100011101;
    W_ir[8][1] = 21'b000000000000001111100;
    W_ir[8][2] = 21'b111111111111110011000;
    W_ir[8][3] = 21'b000000000000100011100;
    W_ir[8][4] = 21'b111111111111110110010;
    W_ir[8][5] = 21'b111111111111101110011;
    W_ir[8][6] = 21'b111111111111001000000;
    W_ir[8][7] = 21'b111111111111100001101;
    W_ir[8][8] = 21'b111111111111101110101;
    W_ir[8][9] = 21'b000000000000100101101;
    W_ir[8][10] = 21'b000000000000010001011;
    W_ir[8][11] = 21'b000000000000110111100;
    W_ir[8][12] = 21'b111111111111110001000;
    W_ir[8][13] = 21'b000000000000011100110;
    W_ir[8][14] = 21'b000000000000011100100;
    W_ir[8][15] = 21'b000000000000001100001;
    W_ir[8][16] = 21'b111111111111110101101;
    W_ir[8][17] = 21'b000000000000101011101;
    W_ir[8][18] = 21'b000000000000111111110;
    W_ir[8][19] = 21'b000000000000100011100;
    W_ir[8][20] = 21'b111111111111111001101;
    W_ir[8][21] = 21'b000000000000001011110;
    W_ir[8][22] = 21'b000000000000101100011;
    W_ir[8][23] = 21'b000000000000001010000;
    W_ir[8][24] = 21'b000000000000000011111;
    W_ir[8][25] = 21'b111111111111110101001;
    W_ir[8][26] = 21'b111111111111000100110;
    W_ir[8][27] = 21'b000000000000001101100;
    W_ir[8][28] = 21'b000000000000011111010;
    W_ir[8][29] = 21'b000000000000000010110;
    W_ir[8][30] = 21'b000000000000100111101;
    W_ir[8][31] = 21'b000000000000100001111;
    W_ir[8][32] = 21'b111111111111110110110;
    W_ir[8][33] = 21'b111111111111011011111;
    W_ir[8][34] = 21'b111111111111001110000;
    W_ir[8][35] = 21'b111111111111100111011;
    W_ir[8][36] = 21'b111111111111100100010;
    W_ir[8][37] = 21'b111111111110101101001;
    W_ir[8][38] = 21'b000000000000001110010;
    W_ir[8][39] = 21'b111111111111111011100;
    W_ir[8][40] = 21'b111111111111110100110;
    W_ir[8][41] = 21'b000000000000110110110;
    W_ir[8][42] = 21'b111111111111010101110;
    W_ir[8][43] = 21'b000000000000100010110;
    W_ir[8][44] = 21'b000000000000000000011;
    W_ir[8][45] = 21'b111111111111100000100;
    W_ir[8][46] = 21'b111111111111011010101;
    W_ir[8][47] = 21'b000000000000101010111;
    W_ir[8][48] = 21'b000000000000010001101;
    W_ir[8][49] = 21'b000000000001001011101;
    W_ir[8][50] = 21'b111111111111111111110;
    W_ir[8][51] = 21'b000000000000001111011;
    W_ir[8][52] = 21'b111111111111101101010;
    W_ir[8][53] = 21'b111111111111010001111;
    W_ir[8][54] = 21'b111111111111001011001;
    W_ir[8][55] = 21'b111111111111100101110;
    W_ir[8][56] = 21'b000000000000111011000;
    W_ir[8][57] = 21'b111111111111101101010;
    W_ir[8][58] = 21'b000000000000111100111;
    W_ir[8][59] = 21'b111111111111110010001;
    W_ir[8][60] = 21'b111111111110111010001;
    W_ir[8][61] = 21'b111111111110010010000;
    W_ir[8][62] = 21'b111111111110000000111;
    W_ir[8][63] = 21'b000000000000011011111;
    W_ir[9][0] = 21'b000000000000110010110;
    W_ir[9][1] = 21'b000000000000010001101;
    W_ir[9][2] = 21'b000000000000001011011;
    W_ir[9][3] = 21'b000000000000000000110;
    W_ir[9][4] = 21'b000000000000000111110;
    W_ir[9][5] = 21'b000000000000100110100;
    W_ir[9][6] = 21'b111111111111001101001;
    W_ir[9][7] = 21'b111111111111010110100;
    W_ir[9][8] = 21'b000000000000000001010;
    W_ir[9][9] = 21'b000000000001000000100;
    W_ir[9][10] = 21'b000000000000100001010;
    W_ir[9][11] = 21'b111111111110111100101;
    W_ir[9][12] = 21'b111111111111010111000;
    W_ir[9][13] = 21'b000000000000101011100;
    W_ir[9][14] = 21'b111111111111110010110;
    W_ir[9][15] = 21'b000000000000110011010;
    W_ir[9][16] = 21'b111111111111000011100;
    W_ir[9][17] = 21'b000000000000011101101;
    W_ir[9][18] = 21'b000000000001001000100;
    W_ir[9][19] = 21'b111111111111010100010;
    W_ir[9][20] = 21'b111111111111011001101;
    W_ir[9][21] = 21'b111111111111000100001;
    W_ir[9][22] = 21'b000000000000100011011;
    W_ir[9][23] = 21'b000000000001010011111;
    W_ir[9][24] = 21'b000000000000011111000;
    W_ir[9][25] = 21'b111111111111100001011;
    W_ir[9][26] = 21'b111111111111100110000;
    W_ir[9][27] = 21'b111111111111011110110;
    W_ir[9][28] = 21'b111111111111101010100;
    W_ir[9][29] = 21'b111111111111001101100;
    W_ir[9][30] = 21'b111111111111110001111;
    W_ir[9][31] = 21'b111111111111001100111;
    W_ir[9][32] = 21'b000000000000100111010;
    W_ir[9][33] = 21'b111111111111101111101;
    W_ir[9][34] = 21'b111111111111011111100;
    W_ir[9][35] = 21'b000000000000101001011;
    W_ir[9][36] = 21'b111111111110110110111;
    W_ir[9][37] = 21'b000000000000001010100;
    W_ir[9][38] = 21'b111111111111111110010;
    W_ir[9][39] = 21'b111111111111011111100;
    W_ir[9][40] = 21'b000000000000101101101;
    W_ir[9][41] = 21'b000000000000010111000;
    W_ir[9][42] = 21'b000000000000111011111;
    W_ir[9][43] = 21'b000000000000110011011;
    W_ir[9][44] = 21'b000000000000000011001;
    W_ir[9][45] = 21'b000000000000111010101;
    W_ir[9][46] = 21'b000000000000010000011;
    W_ir[9][47] = 21'b111111111111110010011;
    W_ir[9][48] = 21'b111111111111010001010;
    W_ir[9][49] = 21'b111111111111110110110;
    W_ir[9][50] = 21'b111111111111100101001;
    W_ir[9][51] = 21'b000000000000011101001;
    W_ir[9][52] = 21'b000000000000101011100;
    W_ir[9][53] = 21'b000000000000011000100;
    W_ir[9][54] = 21'b111111111111000011000;
    W_ir[9][55] = 21'b000000000001001100110;
    W_ir[9][56] = 21'b000000000000100110100;
    W_ir[9][57] = 21'b111111111111110000101;
    W_ir[9][58] = 21'b111111111111111011100;
    W_ir[9][59] = 21'b000000000000110111110;
    W_ir[9][60] = 21'b111111111110111011100;
    W_ir[9][61] = 21'b111111111111111100110;
    W_ir[9][62] = 21'b111111111111100100100;
    W_ir[9][63] = 21'b111111111111101000000;
    W_ir[10][0] = 21'b000000000000010110111;
    W_ir[10][1] = 21'b000000000000011111101;
    W_ir[10][2] = 21'b111111111111110100001;
    W_ir[10][3] = 21'b000000000000001100011;
    W_ir[10][4] = 21'b000000000000110011010;
    W_ir[10][5] = 21'b000000000000010110010;
    W_ir[10][6] = 21'b111111111110110110100;
    W_ir[10][7] = 21'b000000000000010111001;
    W_ir[10][8] = 21'b111111111110100000110;
    W_ir[10][9] = 21'b111111111111110011010;
    W_ir[10][10] = 21'b111111111111111110111;
    W_ir[10][11] = 21'b111111111111100011111;
    W_ir[10][12] = 21'b111111111111001000100;
    W_ir[10][13] = 21'b000000000000011001010;
    W_ir[10][14] = 21'b111111111111111100100;
    W_ir[10][15] = 21'b111111111110101001101;
    W_ir[10][16] = 21'b000000000000100001001;
    W_ir[10][17] = 21'b000000000000100101001;
    W_ir[10][18] = 21'b111111111110100001000;
    W_ir[10][19] = 21'b111111111110111100111;
    W_ir[10][20] = 21'b000000000000110100111;
    W_ir[10][21] = 21'b111111111111001101111;
    W_ir[10][22] = 21'b000000000000010101101;
    W_ir[10][23] = 21'b111111111111010000011;
    W_ir[10][24] = 21'b000000000000011001011;
    W_ir[10][25] = 21'b111111111111010100111;
    W_ir[10][26] = 21'b000000000001001010111;
    W_ir[10][27] = 21'b111111111111110011111;
    W_ir[10][28] = 21'b000000000000101101000;
    W_ir[10][29] = 21'b000000000001000110111;
    W_ir[10][30] = 21'b111111111111110110001;
    W_ir[10][31] = 21'b000000000000000000010;
    W_ir[10][32] = 21'b000000000001010111000;
    W_ir[10][33] = 21'b111111111110111110100;
    W_ir[10][34] = 21'b111111111111000010111;
    W_ir[10][35] = 21'b111111111111100010110;
    W_ir[10][36] = 21'b000000000001010000110;
    W_ir[10][37] = 21'b000000000001000010111;
    W_ir[10][38] = 21'b111111111111010110100;
    W_ir[10][39] = 21'b111111111110101011101;
    W_ir[10][40] = 21'b000000000000100011100;
    W_ir[10][41] = 21'b111111111111111011010;
    W_ir[10][42] = 21'b111111111111000011101;
    W_ir[10][43] = 21'b000000000000001011001;
    W_ir[10][44] = 21'b111111111111101011011;
    W_ir[10][45] = 21'b000000000000100110100;
    W_ir[10][46] = 21'b111111111111110001110;
    W_ir[10][47] = 21'b111111111111110001100;
    W_ir[10][48] = 21'b111111111111100111111;
    W_ir[10][49] = 21'b111111111111111111001;
    W_ir[10][50] = 21'b111111111111000011100;
    W_ir[10][51] = 21'b111111111111100110101;
    W_ir[10][52] = 21'b111111111110111111000;
    W_ir[10][53] = 21'b000000000000110110101;
    W_ir[10][54] = 21'b111111111111111000000;
    W_ir[10][55] = 21'b111111111111100011100;
    W_ir[10][56] = 21'b111111111111100100101;
    W_ir[10][57] = 21'b000000000000111001101;
    W_ir[10][58] = 21'b000000000000111101110;
    W_ir[10][59] = 21'b000000000001001101101;
    W_ir[10][60] = 21'b000000000001111001011;
    W_ir[10][61] = 21'b000000000001010001011;
    W_ir[10][62] = 21'b000000000010001011110;
    W_ir[10][63] = 21'b000000000001100111101;
    W_ir[11][0] = 21'b111111111110100110010;
    W_ir[11][1] = 21'b000000000001000001011;
    W_ir[11][2] = 21'b000000000000000100111;
    W_ir[11][3] = 21'b000000000001000111000;
    W_ir[11][4] = 21'b111111111110101110010;
    W_ir[11][5] = 21'b000000000000010001101;
    W_ir[11][6] = 21'b111111111110111000010;
    W_ir[11][7] = 21'b000000000000100111101;
    W_ir[11][8] = 21'b111111111110010001110;
    W_ir[11][9] = 21'b111111111110100110000;
    W_ir[11][10] = 21'b000000000001001010001;
    W_ir[11][11] = 21'b111111111110100110001;
    W_ir[11][12] = 21'b111111111110101000111;
    W_ir[11][13] = 21'b000000000000100101001;
    W_ir[11][14] = 21'b000000000000011111101;
    W_ir[11][15] = 21'b000000000000011111110;
    W_ir[11][16] = 21'b000000000001010101001;
    W_ir[11][17] = 21'b111111111111101110010;
    W_ir[11][18] = 21'b111111111111111111101;
    W_ir[11][19] = 21'b000000000001100101100;
    W_ir[11][20] = 21'b111111111111110000100;
    W_ir[11][21] = 21'b111111111111000011100;
    W_ir[11][22] = 21'b111111111111101001011;
    W_ir[11][23] = 21'b111111111111100010111;
    W_ir[11][24] = 21'b111111111110110000110;
    W_ir[11][25] = 21'b111111111111110001011;
    W_ir[11][26] = 21'b111111111110111111011;
    W_ir[11][27] = 21'b111111111110101111111;
    W_ir[11][28] = 21'b000000000001101001110;
    W_ir[11][29] = 21'b000000000000100011011;
    W_ir[11][30] = 21'b000000000000000110011;
    W_ir[11][31] = 21'b000000000000111010101;
    W_ir[11][32] = 21'b000000000000100010100;
    W_ir[11][33] = 21'b111111111111110000001;
    W_ir[11][34] = 21'b000000000000111001010;
    W_ir[11][35] = 21'b000000000000011100110;
    W_ir[11][36] = 21'b111111111110111011110;
    W_ir[11][37] = 21'b111111111110101101110;
    W_ir[11][38] = 21'b000000000000100010011;
    W_ir[11][39] = 21'b111111111111111101010;
    W_ir[11][40] = 21'b111111111110100000101;
    W_ir[11][41] = 21'b111111111110101100110;
    W_ir[11][42] = 21'b000000000001000001011;
    W_ir[11][43] = 21'b000000000000000101111;
    W_ir[11][44] = 21'b000000000000010110001;
    W_ir[11][45] = 21'b000000000001100011100;
    W_ir[11][46] = 21'b111111111111110111000;
    W_ir[11][47] = 21'b000000000001010000001;
    W_ir[11][48] = 21'b000000000000001001100;
    W_ir[11][49] = 21'b111111111111110110110;
    W_ir[11][50] = 21'b111111111111010100111;
    W_ir[11][51] = 21'b000000000000101100110;
    W_ir[11][52] = 21'b111111111111101100001;
    W_ir[11][53] = 21'b111111111110101111001;
    W_ir[11][54] = 21'b000000000001100010010;
    W_ir[11][55] = 21'b000000000000001111001;
    W_ir[11][56] = 21'b111111111111010001101;
    W_ir[11][57] = 21'b000000000000101101100;
    W_ir[11][58] = 21'b111111111111011001111;
    W_ir[11][59] = 21'b000000000001011000101;
    W_ir[11][60] = 21'b000000000001010111010;
    W_ir[11][61] = 21'b000000000000010100110;
    W_ir[11][62] = 21'b000000000000000111001;
    W_ir[11][63] = 21'b000000000001001011111;
    W_ir[12][0] = 21'b000000000000010100101;
    W_ir[12][1] = 21'b000000000000100111001;
    W_ir[12][2] = 21'b000000000000011101110;
    W_ir[12][3] = 21'b000000000000100011010;
    W_ir[12][4] = 21'b111111111111101101010;
    W_ir[12][5] = 21'b111111111111010101010;
    W_ir[12][6] = 21'b000000000000011100111;
    W_ir[12][7] = 21'b000000000000001111011;
    W_ir[12][8] = 21'b111111111111001000001;
    W_ir[12][9] = 21'b000000000000000101101;
    W_ir[12][10] = 21'b000000000000111110110;
    W_ir[12][11] = 21'b111111111111111111101;
    W_ir[12][12] = 21'b000000000000101000000;
    W_ir[12][13] = 21'b000000000000001011000;
    W_ir[12][14] = 21'b000000000000001001111;
    W_ir[12][15] = 21'b000000000000101110011;
    W_ir[12][16] = 21'b111111111111111000000;
    W_ir[12][17] = 21'b000000000000110111010;
    W_ir[12][18] = 21'b111111111111111000110;
    W_ir[12][19] = 21'b000000000000100100010;
    W_ir[12][20] = 21'b111111111111111000100;
    W_ir[12][21] = 21'b000000000000100001110;
    W_ir[12][22] = 21'b000000000000011000100;
    W_ir[12][23] = 21'b000000000000011000111;
    W_ir[12][24] = 21'b111111111111010111110;
    W_ir[12][25] = 21'b000000000000011110000;
    W_ir[12][26] = 21'b000000000000100010111;
    W_ir[12][27] = 21'b000000000000010110111;
    W_ir[12][28] = 21'b000000000000111000101;
    W_ir[12][29] = 21'b111111111111001011000;
    W_ir[12][30] = 21'b111111111111101101011;
    W_ir[12][31] = 21'b000000000000011001110;
    W_ir[12][32] = 21'b000000000000001100011;
    W_ir[12][33] = 21'b000000000000011110100;
    W_ir[12][34] = 21'b000000000000011110101;
    W_ir[12][35] = 21'b000000000000000110110;
    W_ir[12][36] = 21'b000000000000111111101;
    W_ir[12][37] = 21'b000000000000010100010;
    W_ir[12][38] = 21'b111111111111101110110;
    W_ir[12][39] = 21'b000000000000001111011;
    W_ir[12][40] = 21'b000000000000100101011;
    W_ir[12][41] = 21'b111111111111010000010;
    W_ir[12][42] = 21'b000000000000001111010;
    W_ir[12][43] = 21'b111111111111101000010;
    W_ir[12][44] = 21'b111111111111111110010;
    W_ir[12][45] = 21'b111111111111011100101;
    W_ir[12][46] = 21'b111111111111001110100;
    W_ir[12][47] = 21'b000000000000110111101;
    W_ir[12][48] = 21'b111111111111110001010;
    W_ir[12][49] = 21'b111111111111100111001;
    W_ir[12][50] = 21'b111111111111111001101;
    W_ir[12][51] = 21'b000000000000000000010;
    W_ir[12][52] = 21'b111111111111000110110;
    W_ir[12][53] = 21'b111111111111101010010;
    W_ir[12][54] = 21'b000000000000010000110;
    W_ir[12][55] = 21'b111111111111100111110;
    W_ir[12][56] = 21'b000000000000100110010;
    W_ir[12][57] = 21'b111111111111100101011;
    W_ir[12][58] = 21'b111111111111101011011;
    W_ir[12][59] = 21'b000000000000100010000;
    W_ir[12][60] = 21'b111111111111010101000;
    W_ir[12][61] = 21'b111111111111001101111;
    W_ir[12][62] = 21'b111111111111001100100;
    W_ir[12][63] = 21'b000000000000100001100;
    W_ir[13][0] = 21'b111111111111100010111;
    W_ir[13][1] = 21'b111111111111100110011;
    W_ir[13][2] = 21'b000000000000101111111;
    W_ir[13][3] = 21'b000000000000100101101;
    W_ir[13][4] = 21'b000000000000000101001;
    W_ir[13][5] = 21'b000000000000001111100;
    W_ir[13][6] = 21'b000000000000001101001;
    W_ir[13][7] = 21'b000000000000001000010;
    W_ir[13][8] = 21'b000000000000001010000;
    W_ir[13][9] = 21'b000000000000001001010;
    W_ir[13][10] = 21'b111111111111111000100;
    W_ir[13][11] = 21'b111111111111111111110;
    W_ir[13][12] = 21'b000000000000001011101;
    W_ir[13][13] = 21'b000000000000011100000;
    W_ir[13][14] = 21'b111111111111010101101;
    W_ir[13][15] = 21'b000000000000001000100;
    W_ir[13][16] = 21'b111111111111111111111;
    W_ir[13][17] = 21'b111111111111111111001;
    W_ir[13][18] = 21'b111111111111111100100;
    W_ir[13][19] = 21'b111111111111101100000;
    W_ir[13][20] = 21'b111111111111111100000;
    W_ir[13][21] = 21'b000000000000001011011;
    W_ir[13][22] = 21'b111111111111110000000;
    W_ir[13][23] = 21'b111111111111101000000;
    W_ir[13][24] = 21'b000000000000000000011;
    W_ir[13][25] = 21'b000000000000101110101;
    W_ir[13][26] = 21'b111111111111001100101;
    W_ir[13][27] = 21'b111111111111001110101;
    W_ir[13][28] = 21'b000000000000110101101;
    W_ir[13][29] = 21'b000000000000010000010;
    W_ir[13][30] = 21'b000000000000000011101;
    W_ir[13][31] = 21'b111111111111111111011;
    W_ir[13][32] = 21'b111111111111100001010;
    W_ir[13][33] = 21'b111111111111111101001;
    W_ir[13][34] = 21'b111111111111111011010;
    W_ir[13][35] = 21'b000000000000000011110;
    W_ir[13][36] = 21'b000000000000001111110;
    W_ir[13][37] = 21'b000000000000001001001;
    W_ir[13][38] = 21'b000000000000001100101;
    W_ir[13][39] = 21'b000000000000100000001;
    W_ir[13][40] = 21'b000000000000010011010;
    W_ir[13][41] = 21'b000000000000000000011;
    W_ir[13][42] = 21'b111111111111111101010;
    W_ir[13][43] = 21'b000000000000010000010;
    W_ir[13][44] = 21'b000000000000000110001;
    W_ir[13][45] = 21'b000000000000001100101;
    W_ir[13][46] = 21'b111111111111111100111;
    W_ir[13][47] = 21'b111111111111110111001;
    W_ir[13][48] = 21'b111111111111110110111;
    W_ir[13][49] = 21'b111111111111001010111;
    W_ir[13][50] = 21'b000000000000011110101;
    W_ir[13][51] = 21'b000000000000101010101;
    W_ir[13][52] = 21'b111111111111110011100;
    W_ir[13][53] = 21'b111111111111100111011;
    W_ir[13][54] = 21'b111111111111101000000;
    W_ir[13][55] = 21'b111111111111100100111;
    W_ir[13][56] = 21'b111111111111110000011;
    W_ir[13][57] = 21'b000000000000110010111;
    W_ir[13][58] = 21'b000000000000011101110;
    W_ir[13][59] = 21'b111111111111011111001;
    W_ir[13][60] = 21'b111111111111110111101;
    W_ir[13][61] = 21'b111111111111110010011;
    W_ir[13][62] = 21'b000000000000101011000;
    W_ir[13][63] = 21'b111111111111100111110;
    W_ir[14][0] = 21'b111111111111101001001;
    W_ir[14][1] = 21'b111111111111110000001;
    W_ir[14][2] = 21'b111111111111001001100;
    W_ir[14][3] = 21'b111111111111011110010;
    W_ir[14][4] = 21'b111111111111101101011;
    W_ir[14][5] = 21'b111111111111110111011;
    W_ir[14][6] = 21'b000000000000000101111;
    W_ir[14][7] = 21'b111111111111010111011;
    W_ir[14][8] = 21'b111111111111110101000;
    W_ir[14][9] = 21'b111111111111110101100;
    W_ir[14][10] = 21'b111111111111110100001;
    W_ir[14][11] = 21'b111111111111000101101;
    W_ir[14][12] = 21'b111111111111110110110;
    W_ir[14][13] = 21'b000000000000001101111;
    W_ir[14][14] = 21'b111111111111110101000;
    W_ir[14][15] = 21'b000000000000010110000;
    W_ir[14][16] = 21'b111111111111010110100;
    W_ir[14][17] = 21'b000000000000111001011;
    W_ir[14][18] = 21'b000000000000000011000;
    W_ir[14][19] = 21'b000000000000010011000;
    W_ir[14][20] = 21'b000000000000001101111;
    W_ir[14][21] = 21'b111111111111101110000;
    W_ir[14][22] = 21'b000000000000011110000;
    W_ir[14][23] = 21'b000000000000110101000;
    W_ir[14][24] = 21'b000000000000011011000;
    W_ir[14][25] = 21'b000000000000001000111;
    W_ir[14][26] = 21'b111111111111111100000;
    W_ir[14][27] = 21'b111111111111001011011;
    W_ir[14][28] = 21'b111111111111110001000;
    W_ir[14][29] = 21'b000000000000111100011;
    W_ir[14][30] = 21'b111111111111101000000;
    W_ir[14][31] = 21'b111111111111101000010;
    W_ir[14][32] = 21'b000000000000000010110;
    W_ir[14][33] = 21'b000000000000010111000;
    W_ir[14][34] = 21'b111111111111110100010;
    W_ir[14][35] = 21'b111111111111110010100;
    W_ir[14][36] = 21'b000000000000000011000;
    W_ir[14][37] = 21'b000000000000001010101;
    W_ir[14][38] = 21'b000000000000100000000;
    W_ir[14][39] = 21'b111111111111111111101;
    W_ir[14][40] = 21'b000000000000011100100;
    W_ir[14][41] = 21'b111111111111110010101;
    W_ir[14][42] = 21'b000000000000011101101;
    W_ir[14][43] = 21'b111111111111111100110;
    W_ir[14][44] = 21'b000000000000001011010;
    W_ir[14][45] = 21'b000000000000001111111;
    W_ir[14][46] = 21'b000000000000001100100;
    W_ir[14][47] = 21'b000000000000000110100;
    W_ir[14][48] = 21'b000000000000001100111;
    W_ir[14][49] = 21'b000000000000001010111;
    W_ir[14][50] = 21'b111111111111100001100;
    W_ir[14][51] = 21'b000000000000010101110;
    W_ir[14][52] = 21'b000000000000010100100;
    W_ir[14][53] = 21'b000000000000001110010;
    W_ir[14][54] = 21'b111111111111001001010;
    W_ir[14][55] = 21'b000000000000010010110;
    W_ir[14][56] = 21'b000000000000001100100;
    W_ir[14][57] = 21'b111111111111010111010;
    W_ir[14][58] = 21'b111111111111100001111;
    W_ir[14][59] = 21'b111111111111100101101;
    W_ir[14][60] = 21'b000000000000100110011;
    W_ir[14][61] = 21'b000000000000010001100;
    W_ir[14][62] = 21'b000000000000100111110;
    W_ir[14][63] = 21'b000000000001000110101;
    W_ir[15][0] = 21'b111111111111111101111;
    W_ir[15][1] = 21'b000000000000111111011;
    W_ir[15][2] = 21'b000000000000000000001;
    W_ir[15][3] = 21'b000000000000110010101;
    W_ir[15][4] = 21'b111111111111010010000;
    W_ir[15][5] = 21'b000000000000001010011;
    W_ir[15][6] = 21'b000000000000000111101;
    W_ir[15][7] = 21'b111111111111101100111;
    W_ir[15][8] = 21'b111111111111111000110;
    W_ir[15][9] = 21'b000000000000101001101;
    W_ir[15][10] = 21'b111111111111100010011;
    W_ir[15][11] = 21'b111111111111111010100;
    W_ir[15][12] = 21'b111111111111011111101;
    W_ir[15][13] = 21'b111111111111110101001;
    W_ir[15][14] = 21'b111111111111110001111;
    W_ir[15][15] = 21'b111111111111111000110;
    W_ir[15][16] = 21'b000000000000000010011;
    W_ir[15][17] = 21'b000000000000001010110;
    W_ir[15][18] = 21'b111111111111101001110;
    W_ir[15][19] = 21'b000000000000100000100;
    W_ir[15][20] = 21'b111111111111110011000;
    W_ir[15][21] = 21'b000000000000001100111;
    W_ir[15][22] = 21'b000000000000010101001;
    W_ir[15][23] = 21'b000000000000001101101;
    W_ir[15][24] = 21'b000000000000110101001;
    W_ir[15][25] = 21'b000000000000001011101;
    W_ir[15][26] = 21'b111111111111111000100;
    W_ir[15][27] = 21'b111111111111101100101;
    W_ir[15][28] = 21'b000000000000001011011;
    W_ir[15][29] = 21'b000000000000001001100;
    W_ir[15][30] = 21'b111111111111011110000;
    W_ir[15][31] = 21'b000000000001000010010;
    W_ir[15][32] = 21'b000000000000100010000;
    W_ir[15][33] = 21'b111111111111011000101;
    W_ir[15][34] = 21'b000000000000010000000;
    W_ir[15][35] = 21'b000000000000001001010;
    W_ir[15][36] = 21'b000000000000001011110;
    W_ir[15][37] = 21'b111111111111000111111;
    W_ir[15][38] = 21'b000000000000011000100;
    W_ir[15][39] = 21'b000000000000000011101;
    W_ir[15][40] = 21'b111111111111111110111;
    W_ir[15][41] = 21'b000000000000100101011;
    W_ir[15][42] = 21'b111111111111010110010;
    W_ir[15][43] = 21'b000000000000000110000;
    W_ir[15][44] = 21'b111111111111101010000;
    W_ir[15][45] = 21'b111111111111101110001;
    W_ir[15][46] = 21'b000000000000110001100;
    W_ir[15][47] = 21'b111111111111101000111;
    W_ir[15][48] = 21'b111111111111110010100;
    W_ir[15][49] = 21'b111111111111110110011;
    W_ir[15][50] = 21'b111111111111100100000;
    W_ir[15][51] = 21'b111111111111101000001;
    W_ir[15][52] = 21'b111111111111100101111;
    W_ir[15][53] = 21'b111111111111100010111;
    W_ir[15][54] = 21'b111111111111101111011;
    W_ir[15][55] = 21'b111111111111000110000;
    W_ir[15][56] = 21'b111111111111100100110;
    W_ir[15][57] = 21'b000000000000011111010;
    W_ir[15][58] = 21'b111111111111011100111;
    W_ir[15][59] = 21'b111111111111100111001;
    W_ir[15][60] = 21'b111111111111101000000;
    W_ir[15][61] = 21'b111111111111101011011;
    W_ir[15][62] = 21'b111111111111010000010;
    W_ir[15][63] = 21'b111111111111101100000;

    // Initialize W_iz weights
    W_iz[0][0] = 21'b111111111111111100100;
    W_iz[0][1] = 21'b111111111111110011011;
    W_iz[0][2] = 21'b111111111111110110110;
    W_iz[0][3] = 21'b111111111111100111010;
    W_iz[0][4] = 21'b000000000000000001010;
    W_iz[0][5] = 21'b000000000000010111001;
    W_iz[0][6] = 21'b111111111111100011011;
    W_iz[0][7] = 21'b111111111111010111010;
    W_iz[0][8] = 21'b111111111111000101000;
    W_iz[0][9] = 21'b111111111111101001011;
    W_iz[0][10] = 21'b111111111111001011100;
    W_iz[0][11] = 21'b111111111111101111000;
    W_iz[0][12] = 21'b111111111111110110101;
    W_iz[0][13] = 21'b000000000000010111000;
    W_iz[0][14] = 21'b000000000000000110010;
    W_iz[0][15] = 21'b111111111111110110101;
    W_iz[0][16] = 21'b111111111111100000110;
    W_iz[0][17] = 21'b111111111111101000101;
    W_iz[0][18] = 21'b111111111111100001101;
    W_iz[0][19] = 21'b111111111111011010101;
    W_iz[0][20] = 21'b111111111111110111001;
    W_iz[0][21] = 21'b000000000000011010110;
    W_iz[0][22] = 21'b000000000001000011110;
    W_iz[0][23] = 21'b000000000000100101100;
    W_iz[0][24] = 21'b111111111111001000001;
    W_iz[0][25] = 21'b111111111111010010111;
    W_iz[0][26] = 21'b000000000000000011101;
    W_iz[0][27] = 21'b111111111111001000001;
    W_iz[0][28] = 21'b000000000000101111101;
    W_iz[0][29] = 21'b111111111111111101101;
    W_iz[0][30] = 21'b000000000000101101100;
    W_iz[0][31] = 21'b111111111111100001001;
    W_iz[0][32] = 21'b111111111111001100000;
    W_iz[0][33] = 21'b111111111111010010101;
    W_iz[0][34] = 21'b111111111111100001100;
    W_iz[0][35] = 21'b111111111111011110111;
    W_iz[0][36] = 21'b111111111111001101101;
    W_iz[0][37] = 21'b111111111111010101011;
    W_iz[0][38] = 21'b111111111111100100100;
    W_iz[0][39] = 21'b000000000000010001010;
    W_iz[0][40] = 21'b000000000000001100000;
    W_iz[0][41] = 21'b111111111111100011001;
    W_iz[0][42] = 21'b111111111111111011111;
    W_iz[0][43] = 21'b111111111111101001111;
    W_iz[0][44] = 21'b111111111111000010010;
    W_iz[0][45] = 21'b111111111111110101100;
    W_iz[0][46] = 21'b111111111111110101010;
    W_iz[0][47] = 21'b111111111111111000011;
    W_iz[0][48] = 21'b000000000000000000001;
    W_iz[0][49] = 21'b111111111111110010100;
    W_iz[0][50] = 21'b000000000000101001110;
    W_iz[0][51] = 21'b111111111111100111000;
    W_iz[0][52] = 21'b000000000000111010100;
    W_iz[0][53] = 21'b000000000000011100010;
    W_iz[0][54] = 21'b000000000000111101100;
    W_iz[0][55] = 21'b000000000000110011011;
    W_iz[0][56] = 21'b000000000000010100001;
    W_iz[0][57] = 21'b111111111111001000100;
    W_iz[0][58] = 21'b000000000000100000111;
    W_iz[0][59] = 21'b000000000001101110110;
    W_iz[0][60] = 21'b000000000001010010110;
    W_iz[0][61] = 21'b000000000001010111011;
    W_iz[0][62] = 21'b000000000001100111001;
    W_iz[0][63] = 21'b000000000001011100000;
    W_iz[1][0] = 21'b000000000000001010100;
    W_iz[1][1] = 21'b000000000000001011011;
    W_iz[1][2] = 21'b000000000000001101011;
    W_iz[1][3] = 21'b111111111111111000010;
    W_iz[1][4] = 21'b111111111111110111011;
    W_iz[1][5] = 21'b111111111111011011000;
    W_iz[1][6] = 21'b000000000000110001111;
    W_iz[1][7] = 21'b111111111111000101010;
    W_iz[1][8] = 21'b111111111111010010100;
    W_iz[1][9] = 21'b111111111111101111011;
    W_iz[1][10] = 21'b111111111111111110101;
    W_iz[1][11] = 21'b111111111111110110101;
    W_iz[1][12] = 21'b111111111111011100001;
    W_iz[1][13] = 21'b111111111111110101100;
    W_iz[1][14] = 21'b111111111111100001000;
    W_iz[1][15] = 21'b111111111111011111111;
    W_iz[1][16] = 21'b000000000000100101000;
    W_iz[1][17] = 21'b111111111111010111110;
    W_iz[1][18] = 21'b000000000000000111110;
    W_iz[1][19] = 21'b111111111111001101111;
    W_iz[1][20] = 21'b111111111111110110000;
    W_iz[1][21] = 21'b000000000000000001011;
    W_iz[1][22] = 21'b000000000000010100101;
    W_iz[1][23] = 21'b000000000000001100111;
    W_iz[1][24] = 21'b111111111111111011000;
    W_iz[1][25] = 21'b111111111111100111101;
    W_iz[1][26] = 21'b111111111111111011010;
    W_iz[1][27] = 21'b000000000000010111010;
    W_iz[1][28] = 21'b000000000000000101000;
    W_iz[1][29] = 21'b111111111111100010100;
    W_iz[1][30] = 21'b111111111111110001000;
    W_iz[1][31] = 21'b111111111111001000100;
    W_iz[1][32] = 21'b111111111111111100011;
    W_iz[1][33] = 21'b111111111111000000001;
    W_iz[1][34] = 21'b111111111111101111111;
    W_iz[1][35] = 21'b000000000000011111001;
    W_iz[1][36] = 21'b111111111111100000100;
    W_iz[1][37] = 21'b111111111111010001001;
    W_iz[1][38] = 21'b111111111110111010011;
    W_iz[1][39] = 21'b000000000000101000111;
    W_iz[1][40] = 21'b111111111111101011101;
    W_iz[1][41] = 21'b111111111111111000000;
    W_iz[1][42] = 21'b000000000000000011011;
    W_iz[1][43] = 21'b111111111111101001100;
    W_iz[1][44] = 21'b000000000000001000010;
    W_iz[1][45] = 21'b111111111111101010100;
    W_iz[1][46] = 21'b111111111111110110110;
    W_iz[1][47] = 21'b000000000000011110100;
    W_iz[1][48] = 21'b000000000000001111010;
    W_iz[1][49] = 21'b000000000000001100100;
    W_iz[1][50] = 21'b000000000000001010101;
    W_iz[1][51] = 21'b000000000000001011001;
    W_iz[1][52] = 21'b111111111111101110110;
    W_iz[1][53] = 21'b111111111111101011100;
    W_iz[1][54] = 21'b000000000000001110101;
    W_iz[1][55] = 21'b000000000000000000001;
    W_iz[1][56] = 21'b000000000000001011000;
    W_iz[1][57] = 21'b111111111111011011111;
    W_iz[1][58] = 21'b111111111111011110011;
    W_iz[1][59] = 21'b111111111111101101100;
    W_iz[1][60] = 21'b000000000000111011101;
    W_iz[1][61] = 21'b000000000000101000100;
    W_iz[1][62] = 21'b111111111111101100000;
    W_iz[1][63] = 21'b000000000000100100010;
    W_iz[2][0] = 21'b000000000000101110101;
    W_iz[2][1] = 21'b111111111111110011101;
    W_iz[2][2] = 21'b000000000001001010111;
    W_iz[2][3] = 21'b111111111111101100111;
    W_iz[2][4] = 21'b000000000000101010000;
    W_iz[2][5] = 21'b000000000000001001111;
    W_iz[2][6] = 21'b111111111111001011000;
    W_iz[2][7] = 21'b000000000001001011000;
    W_iz[2][8] = 21'b000000000001010110010;
    W_iz[2][9] = 21'b000000000000110010101;
    W_iz[2][10] = 21'b000000000000111101101;
    W_iz[2][11] = 21'b111111111111111110100;
    W_iz[2][12] = 21'b000000000000000000111;
    W_iz[2][13] = 21'b000000000000010010101;
    W_iz[2][14] = 21'b111111111111101110000;
    W_iz[2][15] = 21'b111111111111001011100;
    W_iz[2][16] = 21'b111111111111101010010;
    W_iz[2][17] = 21'b000000000000100111011;
    W_iz[2][18] = 21'b111111111111111110101;
    W_iz[2][19] = 21'b111111111111111101001;
    W_iz[2][20] = 21'b111111111111110100011;
    W_iz[2][21] = 21'b111111111111010101011;
    W_iz[2][22] = 21'b000000000001000101100;
    W_iz[2][23] = 21'b111111111111111101100;
    W_iz[2][24] = 21'b111111111111010111010;
    W_iz[2][25] = 21'b000000000000010100001;
    W_iz[2][26] = 21'b111111111111010011110;
    W_iz[2][27] = 21'b111111111111011110000;
    W_iz[2][28] = 21'b000000000000110000111;
    W_iz[2][29] = 21'b000000000000101010010;
    W_iz[2][30] = 21'b111111111111010110000;
    W_iz[2][31] = 21'b000000000000100110100;
    W_iz[2][32] = 21'b000000000000000011011;
    W_iz[2][33] = 21'b000000000000010100010;
    W_iz[2][34] = 21'b000000000000110101101;
    W_iz[2][35] = 21'b000000000001000000010;
    W_iz[2][36] = 21'b111111111111111011001;
    W_iz[2][37] = 21'b000000000000001111101;
    W_iz[2][38] = 21'b111111111111000001011;
    W_iz[2][39] = 21'b111111111111111001101;
    W_iz[2][40] = 21'b000000000000011111111;
    W_iz[2][41] = 21'b111111111111100111100;
    W_iz[2][42] = 21'b000000000001000111000;
    W_iz[2][43] = 21'b000000000000010001000;
    W_iz[2][44] = 21'b000000000000100010001;
    W_iz[2][45] = 21'b111111111111100010100;
    W_iz[2][46] = 21'b111111111111001011101;
    W_iz[2][47] = 21'b000000000000111111111;
    W_iz[2][48] = 21'b111111111111010000001;
    W_iz[2][49] = 21'b111111111111100010010;
    W_iz[2][50] = 21'b000000000000100000010;
    W_iz[2][51] = 21'b111111111111111011011;
    W_iz[2][52] = 21'b000000000000100010000;
    W_iz[2][53] = 21'b111111111110010011000;
    W_iz[2][54] = 21'b111111111111110001011;
    W_iz[2][55] = 21'b000000000000001001101;
    W_iz[2][56] = 21'b111111111111011001011;
    W_iz[2][57] = 21'b111111111111101110001;
    W_iz[2][58] = 21'b111111111111010111000;
    W_iz[2][59] = 21'b111111111111010000100;
    W_iz[2][60] = 21'b111111111111110001011;
    W_iz[2][61] = 21'b111111111110011110000;
    W_iz[2][62] = 21'b111111111110001010000;
    W_iz[2][63] = 21'b111111111110000011000;
    W_iz[3][0] = 21'b111111111110101001010;
    W_iz[3][1] = 21'b111111111110100110001;
    W_iz[3][2] = 21'b000000000000011000111;
    W_iz[3][3] = 21'b111111111111110011001;
    W_iz[3][4] = 21'b000000000000110001101;
    W_iz[3][5] = 21'b000000000001000011110;
    W_iz[3][6] = 21'b111111111111001001011;
    W_iz[3][7] = 21'b000000000000001101000;
    W_iz[3][8] = 21'b111111111111010111011;
    W_iz[3][9] = 21'b111111111110011100101;
    W_iz[3][10] = 21'b111111111111011101111;
    W_iz[3][11] = 21'b000000000000100111101;
    W_iz[3][12] = 21'b000000000000101111110;
    W_iz[3][13] = 21'b111111111111010011011;
    W_iz[3][14] = 21'b000000000000110000100;
    W_iz[3][15] = 21'b111111111111111111111;
    W_iz[3][16] = 21'b000000000000001001111;
    W_iz[3][17] = 21'b111111111111101000000;
    W_iz[3][18] = 21'b000000000000001001110;
    W_iz[3][19] = 21'b000000000000111010110;
    W_iz[3][20] = 21'b111111111111100011111;
    W_iz[3][21] = 21'b111111111111101000101;
    W_iz[3][22] = 21'b000000000000111111011;
    W_iz[3][23] = 21'b111111111111100101010;
    W_iz[3][24] = 21'b000000000000111001000;
    W_iz[3][25] = 21'b000000000000011011100;
    W_iz[3][26] = 21'b000000000000100010101;
    W_iz[3][27] = 21'b111111111111110001110;
    W_iz[3][28] = 21'b000000000000101101010;
    W_iz[3][29] = 21'b000000000001000100010;
    W_iz[3][30] = 21'b000000000000101100101;
    W_iz[3][31] = 21'b000000000000011000000;
    W_iz[3][32] = 21'b111111111111010111010;
    W_iz[3][33] = 21'b111111111111100111011;
    W_iz[3][34] = 21'b111111111110100011110;
    W_iz[3][35] = 21'b111111111111001101001;
    W_iz[3][36] = 21'b000000000000111100101;
    W_iz[3][37] = 21'b000000000000000000100;
    W_iz[3][38] = 21'b000000000000110011010;
    W_iz[3][39] = 21'b111111111110111011111;
    W_iz[3][40] = 21'b111111111111111101110;
    W_iz[3][41] = 21'b111111111110111110000;
    W_iz[3][42] = 21'b111111111110111001101;
    W_iz[3][43] = 21'b111111111110110111000;
    W_iz[3][44] = 21'b111111111111011010100;
    W_iz[3][45] = 21'b000000000000001001101;
    W_iz[3][46] = 21'b000000000010001100001;
    W_iz[3][47] = 21'b111111111111011010011;
    W_iz[3][48] = 21'b111111111111111001110;
    W_iz[3][49] = 21'b111111111111010110100;
    W_iz[3][50] = 21'b111111111111000010100;
    W_iz[3][51] = 21'b000000000001011101100;
    W_iz[3][52] = 21'b111111111110111010011;
    W_iz[3][53] = 21'b000000000000010110001;
    W_iz[3][54] = 21'b000000000001000111000;
    W_iz[3][55] = 21'b000000000000001011010;
    W_iz[3][56] = 21'b000000000010010001011;
    W_iz[3][57] = 21'b000000000000010010011;
    W_iz[3][58] = 21'b000000000010010100011;
    W_iz[3][59] = 21'b000000000000010111101;
    W_iz[3][60] = 21'b111111111111000010100;
    W_iz[3][61] = 21'b000000000001000111000;
    W_iz[3][62] = 21'b000000000001100000011;
    W_iz[3][63] = 21'b111111111111000010100;
    W_iz[4][0] = 21'b111111111111100011101;
    W_iz[4][1] = 21'b000000000000001111100;
    W_iz[4][2] = 21'b111111111111110011000;
    W_iz[4][3] = 21'b000000000000100011100;
    W_iz[4][4] = 21'b111111111111110110010;
    W_iz[4][5] = 21'b111111111111101110011;
    W_iz[4][6] = 21'b111111111111001000000;
    W_iz[4][7] = 21'b111111111111100001101;
    W_iz[4][8] = 21'b111111111111101110101;
    W_iz[4][9] = 21'b000000000000100101101;
    W_iz[4][10] = 21'b000000000000010001011;
    W_iz[4][11] = 21'b000000000000110111100;
    W_iz[4][12] = 21'b111111111111110001000;
    W_iz[4][13] = 21'b000000000000011100110;
    W_iz[4][14] = 21'b000000000000011100100;
    W_iz[4][15] = 21'b000000000000001100001;
    W_iz[4][16] = 21'b111111111111110101101;
    W_iz[4][17] = 21'b000000000000101011101;
    W_iz[4][18] = 21'b000000000000111111110;
    W_iz[4][19] = 21'b000000000000100011100;
    W_iz[4][20] = 21'b111111111111111001101;
    W_iz[4][21] = 21'b000000000000001011110;
    W_iz[4][22] = 21'b000000000000101100011;
    W_iz[4][23] = 21'b000000000000001010000;
    W_iz[4][24] = 21'b000000000000000011111;
    W_iz[4][25] = 21'b111111111111110101001;
    W_iz[4][26] = 21'b111111111111000100110;
    W_iz[4][27] = 21'b000000000000001101100;
    W_iz[4][28] = 21'b000000000000011111010;
    W_iz[4][29] = 21'b000000000000000010110;
    W_iz[4][30] = 21'b000000000000100111101;
    W_iz[4][31] = 21'b000000000000100001111;
    W_iz[4][32] = 21'b111111111111110110110;
    W_iz[4][33] = 21'b111111111111011011111;
    W_iz[4][34] = 21'b111111111111001110000;
    W_iz[4][35] = 21'b111111111111100111011;
    W_iz[4][36] = 21'b111111111111100100010;
    W_iz[4][37] = 21'b111111111110101101001;
    W_iz[4][38] = 21'b000000000000001110010;
    W_iz[4][39] = 21'b111111111111111011100;
    W_iz[4][40] = 21'b111111111111110100110;
    W_iz[4][41] = 21'b000000000000110110110;
    W_iz[4][42] = 21'b111111111111010101110;
    W_iz[4][43] = 21'b000000000000100010110;
    W_iz[4][44] = 21'b000000000000000000011;
    W_iz[4][45] = 21'b111111111111100000100;
    W_iz[4][46] = 21'b111111111111011010101;
    W_iz[4][47] = 21'b000000000000101010111;
    W_iz[4][48] = 21'b000000000000010001101;
    W_iz[4][49] = 21'b000000000001001011101;
    W_iz[4][50] = 21'b111111111111111111110;
    W_iz[4][51] = 21'b000000000000001111011;
    W_iz[4][52] = 21'b111111111111101101010;
    W_iz[4][53] = 21'b111111111111010001111;
    W_iz[4][54] = 21'b111111111111001011001;
    W_iz[4][55] = 21'b111111111111100101110;
    W_iz[4][56] = 21'b000000000000111011000;
    W_iz[4][57] = 21'b111111111111101101010;
    W_iz[4][58] = 21'b000000000000111100111;
    W_iz[4][59] = 21'b111111111111110010001;
    W_iz[4][60] = 21'b111111111110111010001;
    W_iz[4][61] = 21'b111111111110010010000;
    W_iz[4][62] = 21'b111111111110000000111;
    W_iz[4][63] = 21'b000000000000011011111;
    W_iz[5][0] = 21'b000000000000110010110;
    W_iz[5][1] = 21'b000000000000010001101;
    W_iz[5][2] = 21'b000000000000001011011;
    W_iz[5][3] = 21'b000000000000000000110;
    W_iz[5][4] = 21'b000000000000000111110;
    W_iz[5][5] = 21'b000000000000100110100;
    W_iz[5][6] = 21'b111111111111001101001;
    W_iz[5][7] = 21'b111111111111010110100;
    W_iz[5][8] = 21'b000000000000000001010;
    W_iz[5][9] = 21'b000000000001000000100;
    W_iz[5][10] = 21'b000000000000100001010;
    W_iz[5][11] = 21'b111111111110111100101;
    W_iz[5][12] = 21'b111111111111010111000;
    W_iz[5][13] = 21'b000000000000101011100;
    W_iz[5][14] = 21'b111111111111110010110;
    W_iz[5][15] = 21'b000000000000110011010;
    W_iz[5][16] = 21'b111111111111000011100;
    W_iz[5][17] = 21'b000000000000011101101;
    W_iz[5][18] = 21'b000000000001001000100;
    W_iz[5][19] = 21'b111111111111010100010;
    W_iz[5][20] = 21'b111111111111011001101;
    W_iz[5][21] = 21'b111111111111000100001;
    W_iz[5][22] = 21'b000000000000100011011;
    W_iz[5][23] = 21'b000000000001010011111;
    W_iz[5][24] = 21'b000000000000011111000;
    W_iz[5][25] = 21'b111111111111100001011;
    W_iz[5][26] = 21'b111111111111100110000;
    W_iz[5][27] = 21'b111111111111011110110;
    W_iz[5][28] = 21'b111111111111101010100;
    W_iz[5][29] = 21'b111111111111001101100;
    W_iz[5][30] = 21'b111111111111110001111;
    W_iz[5][31] = 21'b111111111111001100111;
    W_iz[5][32] = 21'b000000000000100111010;
    W_iz[5][33] = 21'b111111111111101111101;
    W_iz[5][34] = 21'b111111111111011111100;
    W_iz[5][35] = 21'b000000000000101001011;
    W_iz[5][36] = 21'b111111111110110110111;
    W_iz[5][37] = 21'b000000000000001010100;
    W_iz[5][38] = 21'b111111111111111110010;
    W_iz[5][39] = 21'b111111111111011111100;
    W_iz[5][40] = 21'b000000000000101101101;
    W_iz[5][41] = 21'b000000000000010111000;
    W_iz[5][42] = 21'b000000000000111011111;
    W_iz[5][43] = 21'b000000000000110011011;
    W_iz[5][44] = 21'b000000000000000011001;
    W_iz[5][45] = 21'b000000000000111010101;
    W_iz[5][46] = 21'b000000000000010000011;
    W_iz[5][47] = 21'b111111111111110010011;
    W_iz[5][48] = 21'b111111111111010001010;
    W_iz[5][49] = 21'b111111111111110110110;
    W_iz[5][50] = 21'b111111111111100101001;
    W_iz[5][51] = 21'b000000000000011101001;
    W_iz[5][52] = 21'b000000000000101011100;
    W_iz[5][53] = 21'b000000000000011000100;
    W_iz[5][54] = 21'b111111111111000011000;
    W_iz[5][55] = 21'b000000000001001100110;
    W_iz[5][56] = 21'b000000000000100110100;
    W_iz[5][57] = 21'b111111111111110000101;
    W_iz[5][58] = 21'b111111111111111011100;
    W_iz[5][59] = 21'b000000000000110111110;
    W_iz[5][60] = 21'b111111111110111011100;
    W_iz[5][61] = 21'b111111111111111100110;
    W_iz[5][62] = 21'b111111111111100100100;
    W_iz[5][63] = 21'b111111111111101000000;
    W_iz[6][0] = 21'b000000000000010110111;
    W_iz[6][1] = 21'b000000000000011111101;
    W_iz[6][2] = 21'b111111111111110100001;
    W_iz[6][3] = 21'b000000000000001100011;
    W_iz[6][4] = 21'b000000000000110011010;
    W_iz[6][5] = 21'b000000000000010110010;
    W_iz[6][6] = 21'b111111111110110110100;
    W_iz[6][7] = 21'b000000000000010111001;
    W_iz[6][8] = 21'b111111111110100000110;
    W_iz[6][9] = 21'b111111111111110011010;
    W_iz[6][10] = 21'b111111111111111110111;
    W_iz[6][11] = 21'b111111111111100011111;
    W_iz[6][12] = 21'b111111111111001000100;
    W_iz[6][13] = 21'b000000000000011001010;
    W_iz[6][14] = 21'b111111111111111100100;
    W_iz[6][15] = 21'b111111111110101001101;
    W_iz[6][16] = 21'b000000000000100001001;
    W_iz[6][17] = 21'b000000000000100101001;
    W_iz[6][18] = 21'b111111111110100001000;
    W_iz[6][19] = 21'b111111111110111100111;
    W_iz[6][20] = 21'b000000000000110100111;
    W_iz[6][21] = 21'b111111111111001101111;
    W_iz[6][22] = 21'b000000000000010101101;
    W_iz[6][23] = 21'b111111111111010000011;
    W_iz[6][24] = 21'b000000000000011001011;
    W_iz[6][25] = 21'b111111111111010100111;
    W_iz[6][26] = 21'b000000000001001010111;
    W_iz[6][27] = 21'b111111111111110011111;
    W_iz[6][28] = 21'b000000000000101101000;
    W_iz[6][29] = 21'b000000000001000110111;
    W_iz[6][30] = 21'b111111111111110110001;
    W_iz[6][31] = 21'b000000000000000000010;
    W_iz[6][32] = 21'b000000000001010111000;
    W_iz[6][33] = 21'b111111111110111110100;
    W_iz[6][34] = 21'b111111111111000010111;
    W_iz[6][35] = 21'b111111111111100010110;
    W_iz[6][36] = 21'b000000000001010000110;
    W_iz[6][37] = 21'b000000000001000010111;
    W_iz[6][38] = 21'b111111111111010110100;
    W_iz[6][39] = 21'b111111111110101011101;
    W_iz[6][40] = 21'b000000000000100011100;
    W_iz[6][41] = 21'b111111111111111011010;
    W_iz[6][42] = 21'b111111111111000011101;
    W_iz[6][43] = 21'b000000000000001011001;
    W_iz[6][44] = 21'b111111111111101011011;
    W_iz[6][45] = 21'b000000000000100110100;
    W_iz[6][46] = 21'b111111111111110001110;
    W_iz[6][47] = 21'b111111111111110001100;
    W_iz[6][48] = 21'b111111111111100111111;
    W_iz[6][49] = 21'b111111111111111111001;
    W_iz[6][50] = 21'b111111111111000011100;
    W_iz[6][51] = 21'b111111111111100110101;
    W_iz[6][52] = 21'b111111111110111111000;
    W_iz[6][53] = 21'b000000000000110110101;
    W_iz[6][54] = 21'b111111111111111000000;
    W_iz[6][55] = 21'b111111111111100011100;
    W_iz[6][56] = 21'b111111111111100100101;
    W_iz[6][57] = 21'b000000000000111001101;
    W_iz[6][58] = 21'b000000000000111101110;
    W_iz[6][59] = 21'b000000000001001101101;
    W_iz[6][60] = 21'b000000000001111001011;
    W_iz[6][61] = 21'b000000000001010001011;
    W_iz[6][62] = 21'b000000000010001011110;
    W_iz[6][63] = 21'b000000000001100111101;
    W_iz[7][0] = 21'b111111111110100110010;
    W_iz[7][1] = 21'b000000000001000001011;
    W_iz[7][2] = 21'b000000000000000100111;
    W_iz[7][3] = 21'b000000000001000111000;
    W_iz[7][4] = 21'b111111111110101110010;
    W_iz[7][5] = 21'b000000000000010001101;
    W_iz[7][6] = 21'b111111111110111000010;
    W_iz[7][7] = 21'b000000000000100111101;
    W_iz[7][8] = 21'b111111111110010001110;
    W_iz[7][9] = 21'b111111111110100110000;
    W_iz[7][10] = 21'b000000000001001010001;
    W_iz[7][11] = 21'b111111111110100110001;
    W_iz[7][12] = 21'b111111111110101000111;
    W_iz[7][13] = 21'b000000000000100101001;
    W_iz[7][14] = 21'b000000000000011111101;
    W_iz[7][15] = 21'b000000000000011111110;
    W_iz[7][16] = 21'b000000000001010101001;
    W_iz[7][17] = 21'b111111111111101110010;
    W_iz[7][18] = 21'b111111111111111111101;
    W_iz[7][19] = 21'b000000000001100101100;
    W_iz[7][20] = 21'b111111111111110000100;
    W_iz[7][21] = 21'b111111111111000011100;
    W_iz[7][22] = 21'b111111111111101001011;
    W_iz[7][23] = 21'b111111111111100010111;
    W_iz[7][24] = 21'b111111111110110000110;
    W_iz[7][25] = 21'b111111111111110001011;
    W_iz[7][26] = 21'b111111111110111111011;
    W_iz[7][27] = 21'b111111111110101111111;
    W_iz[7][28] = 21'b000000000001101001110;
    W_iz[7][29] = 21'b000000000000100011011;
    W_iz[7][30] = 21'b000000000000000110011;
    W_iz[7][31] = 21'b000000000000111010101;
    W_iz[7][32] = 21'b000000000000100010100;
    W_iz[7][33] = 21'b111111111111110000001;
    W_iz[7][34] = 21'b000000000000111001010;
    W_iz[7][35] = 21'b000000000000011100110;
    W_iz[7][36] = 21'b111111111110111011110;
    W_iz[7][37] = 21'b111111111110101101110;
    W_iz[7][38] = 21'b000000000000100010011;
    W_iz[7][39] = 21'b111111111111111101010;
    W_iz[7][40] = 21'b111111111110100000101;
    W_iz[7][41] = 21'b111111111110101100110;
    W_iz[7][42] = 21'b000000000001000001011;
    W_iz[7][43] = 21'b000000000000000101111;
    W_iz[7][44] = 21'b000000000000010110001;
    W_iz[7][45] = 21'b000000000001100011100;
    W_iz[7][46] = 21'b111111111111110111000;
    W_iz[7][47] = 21'b000000000001010000001;
    W_iz[7][48] = 21'b000000000000001001100;
    W_iz[7][49] = 21'b111111111111110110110;
    W_iz[7][50] = 21'b111111111111010100111;
    W_iz[7][51] = 21'b000000000000101100110;
    W_iz[7][52] = 21'b111111111111101100001;
    W_iz[7][53] = 21'b111111111110101111001;
    W_iz[7][54] = 21'b000000000001100010010;
    W_iz[7][55] = 21'b000000000000001111001;
    W_iz[7][56] = 21'b111111111111010001101;
    W_iz[7][57] = 21'b000000000000101101100;
    W_iz[7][58] = 21'b111111111111011001111;
    W_iz[7][59] = 21'b000000000001011000101;
    W_iz[7][60] = 21'b000000000001010111010;
    W_iz[7][61] = 21'b000000000000010100110;
    W_iz[7][62] = 21'b000000000000000111001;
    W_iz[7][63] = 21'b000000000001001011111;
    W_iz[8][0] = 21'b000000000000010100101;
    W_iz[8][1] = 21'b000000000000100111001;
    W_iz[8][2] = 21'b000000000000011101110;
    W_iz[8][3] = 21'b000000000000100011010;
    W_iz[8][4] = 21'b111111111111101101010;
    W_iz[8][5] = 21'b111111111111010101010;
    W_iz[8][6] = 21'b000000000000011100111;
    W_iz[8][7] = 21'b000000000000001111011;
    W_iz[8][8] = 21'b111111111111001000001;
    W_iz[8][9] = 21'b000000000000000101101;
    W_iz[8][10] = 21'b000000000000111110110;
    W_iz[8][11] = 21'b111111111111111111101;
    W_iz[8][12] = 21'b000000000000101000000;
    W_iz[8][13] = 21'b000000000000001011000;
    W_iz[8][14] = 21'b000000000000001001111;
    W_iz[8][15] = 21'b000000000000101110011;
    W_iz[8][16] = 21'b111111111111111000000;
    W_iz[8][17] = 21'b000000000000110111010;
    W_iz[8][18] = 21'b111111111111111000110;
    W_iz[8][19] = 21'b000000000000100100010;
    W_iz[8][20] = 21'b111111111111111000100;
    W_iz[8][21] = 21'b000000000000100001110;
    W_iz[8][22] = 21'b000000000000011000100;
    W_iz[8][23] = 21'b000000000000011000111;
    W_iz[8][24] = 21'b111111111111010111110;
    W_iz[8][25] = 21'b000000000000011110000;
    W_iz[8][26] = 21'b000000000000100010111;
    W_iz[8][27] = 21'b000000000000010110111;
    W_iz[8][28] = 21'b000000000000111000101;
    W_iz[8][29] = 21'b111111111111001011000;
    W_iz[8][30] = 21'b111111111111101101011;
    W_iz[8][31] = 21'b000000000000011001110;
    W_iz[8][32] = 21'b000000000000001100011;
    W_iz[8][33] = 21'b000000000000011110100;
    W_iz[8][34] = 21'b000000000000011110101;
    W_iz[8][35] = 21'b000000000000000110110;
    W_iz[8][36] = 21'b000000000000111111101;
    W_iz[8][37] = 21'b000000000000010100010;
    W_iz[8][38] = 21'b111111111111101110110;
    W_iz[8][39] = 21'b000000000000001111011;
    W_iz[8][40] = 21'b000000000000100101011;
    W_iz[8][41] = 21'b111111111111010000010;
    W_iz[8][42] = 21'b000000000000001111010;
    W_iz[8][43] = 21'b111111111111101000010;
    W_iz[8][44] = 21'b111111111111111110010;
    W_iz[8][45] = 21'b111111111111011100101;
    W_iz[8][46] = 21'b111111111111001110100;
    W_iz[8][47] = 21'b000000000000110111101;
    W_iz[8][48] = 21'b111111111111110001010;
    W_iz[8][49] = 21'b111111111111100111001;
    W_iz[8][50] = 21'b111111111111111001101;
    W_iz[8][51] = 21'b000000000000000000010;
    W_iz[8][52] = 21'b111111111111000110110;
    W_iz[8][53] = 21'b111111111111101010010;
    W_iz[8][54] = 21'b000000000000010000110;
    W_iz[8][55] = 21'b111111111111100111110;
    W_iz[8][56] = 21'b000000000000100110010;
    W_iz[8][57] = 21'b111111111111100101011;
    W_iz[8][58] = 21'b111111111111101011011;
    W_iz[8][59] = 21'b000000000000100010000;
    W_iz[8][60] = 21'b111111111111010101000;
    W_iz[8][61] = 21'b111111111111001101111;
    W_iz[8][62] = 21'b111111111111001100100;
    W_iz[8][63] = 21'b000000000000100001100;
    W_iz[9][0] = 21'b111111111111100010111;
    W_iz[9][1] = 21'b111111111111100110011;
    W_iz[9][2] = 21'b000000000000101111111;
    W_iz[9][3] = 21'b000000000000100101101;
    W_iz[9][4] = 21'b000000000000000101001;
    W_iz[9][5] = 21'b000000000000001111100;
    W_iz[9][6] = 21'b000000000000001101001;
    W_iz[9][7] = 21'b000000000000001000010;
    W_iz[9][8] = 21'b000000000000001010000;
    W_iz[9][9] = 21'b000000000000001001010;
    W_iz[9][10] = 21'b111111111111111000100;
    W_iz[9][11] = 21'b111111111111111111110;
    W_iz[9][12] = 21'b000000000000001011101;
    W_iz[9][13] = 21'b000000000000011100000;
    W_iz[9][14] = 21'b111111111111010101101;
    W_iz[9][15] = 21'b000000000000001000100;
    W_iz[9][16] = 21'b111111111111111111111;
    W_iz[9][17] = 21'b111111111111111111001;
    W_iz[9][18] = 21'b111111111111111100100;
    W_iz[9][19] = 21'b111111111111101100000;
    W_iz[9][20] = 21'b111111111111111100000;
    W_iz[9][21] = 21'b000000000000001011011;
    W_iz[9][22] = 21'b111111111111110000000;
    W_iz[9][23] = 21'b111111111111101000000;
    W_iz[9][24] = 21'b000000000000000000011;
    W_iz[9][25] = 21'b000000000000101110101;
    W_iz[9][26] = 21'b111111111111001100101;
    W_iz[9][27] = 21'b111111111111001110101;
    W_iz[9][28] = 21'b000000000000110101101;
    W_iz[9][29] = 21'b000000000000010000010;
    W_iz[9][30] = 21'b000000000000000011101;
    W_iz[9][31] = 21'b111111111111111111011;
    W_iz[9][32] = 21'b111111111111100001010;
    W_iz[9][33] = 21'b111111111111111101001;
    W_iz[9][34] = 21'b111111111111111011010;
    W_iz[9][35] = 21'b000000000000000011110;
    W_iz[9][36] = 21'b000000000000001111110;
    W_iz[9][37] = 21'b000000000000001001001;
    W_iz[9][38] = 21'b000000000000001100101;
    W_iz[9][39] = 21'b000000000000100000001;
    W_iz[9][40] = 21'b000000000000010011010;
    W_iz[9][41] = 21'b000000000000000000011;
    W_iz[9][42] = 21'b111111111111111101010;
    W_iz[9][43] = 21'b000000000000010000010;
    W_iz[9][44] = 21'b000000000000000110001;
    W_iz[9][45] = 21'b000000000000001100101;
    W_iz[9][46] = 21'b111111111111111100111;
    W_iz[9][47] = 21'b111111111111110111001;
    W_iz[9][48] = 21'b111111111111110110111;
    W_iz[9][49] = 21'b111111111111001010111;
    W_iz[9][50] = 21'b000000000000011110101;
    W_iz[9][51] = 21'b000000000000101010101;
    W_iz[9][52] = 21'b111111111111110011100;
    W_iz[9][53] = 21'b111111111111100111011;
    W_iz[9][54] = 21'b111111111111101000000;
    W_iz[9][55] = 21'b111111111111100100111;
    W_iz[9][56] = 21'b111111111111110000011;
    W_iz[9][57] = 21'b000000000000110010111;
    W_iz[9][58] = 21'b000000000000011101110;
    W_iz[9][59] = 21'b111111111111011111001;
    W_iz[9][60] = 21'b111111111111110111101;
    W_iz[9][61] = 21'b111111111111110010011;
    W_iz[9][62] = 21'b000000000000101011000;
    W_iz[9][63] = 21'b111111111111100111110;
    W_iz[10][0] = 21'b111111111111101001001;
    W_iz[10][1] = 21'b111111111111110000001;
    W_iz[10][2] = 21'b111111111111001001100;
    W_iz[10][3] = 21'b111111111111011110010;
    W_iz[10][4] = 21'b111111111111101101011;
    W_iz[10][5] = 21'b111111111111110111011;
    W_iz[10][6] = 21'b000000000000000101111;
    W_iz[10][7] = 21'b111111111111010111011;
    W_iz[10][8] = 21'b111111111111110101000;
    W_iz[10][9] = 21'b111111111111110101100;
    W_iz[10][10] = 21'b111111111111110100001;
    W_iz[10][11] = 21'b111111111111000101101;
    W_iz[10][12] = 21'b111111111111110110110;
    W_iz[10][13] = 21'b000000000000001101111;
    W_iz[10][14] = 21'b111111111111110101000;
    W_iz[10][15] = 21'b000000000000010110000;
    W_iz[10][16] = 21'b111111111111010110100;
    W_iz[10][17] = 21'b000000000000111001011;
    W_iz[10][18] = 21'b000000000000000011000;
    W_iz[10][19] = 21'b000000000000010011000;
    W_iz[10][20] = 21'b000000000000001101111;
    W_iz[10][21] = 21'b111111111111101110000;
    W_iz[10][22] = 21'b000000000000011110000;
    W_iz[10][23] = 21'b000000000000110101000;
    W_iz[10][24] = 21'b000000000000011011000;
    W_iz[10][25] = 21'b000000000000001000111;
    W_iz[10][26] = 21'b111111111111111100000;
    W_iz[10][27] = 21'b111111111111001011011;
    W_iz[10][28] = 21'b111111111111110001000;
    W_iz[10][29] = 21'b000000000000111100011;
    W_iz[10][30] = 21'b111111111111101000000;
    W_iz[10][31] = 21'b111111111111101000010;
    W_iz[10][32] = 21'b000000000000000010110;
    W_iz[10][33] = 21'b000000000000010111000;
    W_iz[10][34] = 21'b111111111111110100010;
    W_iz[10][35] = 21'b111111111111110010100;
    W_iz[10][36] = 21'b000000000000000011000;
    W_iz[10][37] = 21'b000000000000001010101;
    W_iz[10][38] = 21'b000000000000100000000;
    W_iz[10][39] = 21'b111111111111111111101;
    W_iz[10][40] = 21'b000000000000011100100;
    W_iz[10][41] = 21'b111111111111110010101;
    W_iz[10][42] = 21'b000000000000011101101;
    W_iz[10][43] = 21'b111111111111111100110;
    W_iz[10][44] = 21'b000000000000001011010;
    W_iz[10][45] = 21'b000000000000001111111;
    W_iz[10][46] = 21'b000000000000001100100;
    W_iz[10][47] = 21'b000000000000000110100;
    W_iz[10][48] = 21'b000000000000001100111;
    W_iz[10][49] = 21'b000000000000001010111;
    W_iz[10][50] = 21'b111111111111100001100;
    W_iz[10][51] = 21'b000000000000010101110;
    W_iz[10][52] = 21'b000000000000010100100;
    W_iz[10][53] = 21'b000000000000001110010;
    W_iz[10][54] = 21'b111111111111001001010;
    W_iz[10][55] = 21'b000000000000010010110;
    W_iz[10][56] = 21'b000000000000001100100;
    W_iz[10][57] = 21'b111111111111010111010;
    W_iz[10][58] = 21'b111111111111100001111;
    W_iz[10][59] = 21'b111111111111100101101;
    W_iz[10][60] = 21'b000000000000100110011;
    W_iz[10][61] = 21'b000000000000010001100;
    W_iz[10][62] = 21'b000000000000100111110;
    W_iz[10][63] = 21'b000000000001000110101;
    W_iz[11][0] = 21'b111111111111111101111;
    W_iz[11][1] = 21'b000000000000111111011;
    W_iz[11][2] = 21'b000000000000000000001;
    W_iz[11][3] = 21'b000000000000110010101;
    W_iz[11][4] = 21'b111111111111010010000;
    W_iz[11][5] = 21'b000000000000001010011;
    W_iz[11][6] = 21'b000000000000000111101;
    W_iz[11][7] = 21'b111111111111101100111;
    W_iz[11][8] = 21'b111111111111111000110;
    W_iz[11][9] = 21'b000000000000101001101;
    W_iz[11][10] = 21'b111111111111100010011;
    W_iz[11][11] = 21'b111111111111111010100;
    W_iz[11][12] = 21'b111111111111011111101;
    W_iz[11][13] = 21'b111111111111110101001;
    W_iz[11][14] = 21'b111111111111110001111;
    W_iz[11][15] = 21'b111111111111111000110;
    W_iz[11][16] = 21'b000000000000000010011;
    W_iz[11][17] = 21'b000000000000001010110;
    W_iz[11][18] = 21'b111111111111101001110;
    W_iz[11][19] = 21'b000000000000100000100;
    W_iz[11][20] = 21'b111111111111110011000;
    W_iz[11][21] = 21'b000000000000001100111;
    W_iz[11][22] = 21'b000000000000010101001;
    W_iz[11][23] = 21'b000000000000001101101;
    W_iz[11][24] = 21'b000000000000110101001;
    W_iz[11][25] = 21'b000000000000001011101;
    W_iz[11][26] = 21'b111111111111111000100;
    W_iz[11][27] = 21'b111111111111101100101;
    W_iz[11][28] = 21'b000000000000001011011;
    W_iz[11][29] = 21'b000000000000001001100;
    W_iz[11][30] = 21'b111111111111011110000;
    W_iz[11][31] = 21'b000000000001000010010;
    W_iz[11][32] = 21'b000000000000100010000;
    W_iz[11][33] = 21'b111111111111011000101;
    W_iz[11][34] = 21'b000000000000010000000;
    W_iz[11][35] = 21'b000000000000001001010;
    W_iz[11][36] = 21'b000000000000001011110;
    W_iz[11][37] = 21'b111111111111000111111;
    W_iz[11][38] = 21'b000000000000011000100;
    W_iz[11][39] = 21'b000000000000000011101;
    W_iz[11][40] = 21'b111111111111111110111;
    W_iz[11][41] = 21'b000000000000100101011;
    W_iz[11][42] = 21'b111111111111010110010;
    W_iz[11][43] = 21'b000000000000000110000;
    W_iz[11][44] = 21'b111111111111101010000;
    W_iz[11][45] = 21'b111111111111101110001;
    W_iz[11][46] = 21'b000000000000110001100;
    W_iz[11][47] = 21'b111111111111101000111;
    W_iz[11][48] = 21'b111111111111110010100;
    W_iz[11][49] = 21'b111111111111110110011;
    W_iz[11][50] = 21'b111111111111100100000;
    W_iz[11][51] = 21'b111111111111101000001;
    W_iz[11][52] = 21'b111111111111100101111;
    W_iz[11][53] = 21'b111111111111100010111;
    W_iz[11][54] = 21'b111111111111101111011;
    W_iz[11][55] = 21'b111111111111000110000;
    W_iz[11][56] = 21'b111111111111100100110;
    W_iz[11][57] = 21'b000000000000011111010;
    W_iz[11][58] = 21'b111111111111011100111;
    W_iz[11][59] = 21'b111111111111100111001;
    W_iz[11][60] = 21'b111111111111101000000;
    W_iz[11][61] = 21'b111111111111101011011;
    W_iz[11][62] = 21'b111111111111010000010;
    W_iz[11][63] = 21'b111111111111101100000;
    W_iz[12][0] = 21'b111111111111111100100;
    W_iz[12][1] = 21'b111111111111110011011;
    W_iz[12][2] = 21'b111111111111110110110;
    W_iz[12][3] = 21'b111111111111100111010;
    W_iz[12][4] = 21'b000000000000000001010;
    W_iz[12][5] = 21'b000000000000010111001;
    W_iz[12][6] = 21'b111111111111100011011;
    W_iz[12][7] = 21'b111111111111010111010;
    W_iz[12][8] = 21'b111111111111000101000;
    W_iz[12][9] = 21'b111111111111101001011;
    W_iz[12][10] = 21'b111111111111001011100;
    W_iz[12][11] = 21'b111111111111101111000;
    W_iz[12][12] = 21'b111111111111110110101;
    W_iz[12][13] = 21'b000000000000010111000;
    W_iz[12][14] = 21'b000000000000000110010;
    W_iz[12][15] = 21'b111111111111110110101;
    W_iz[12][16] = 21'b111111111111100000110;
    W_iz[12][17] = 21'b111111111111101000101;
    W_iz[12][18] = 21'b111111111111100001101;
    W_iz[12][19] = 21'b111111111111011010101;
    W_iz[12][20] = 21'b111111111111110111001;
    W_iz[12][21] = 21'b000000000000011010110;
    W_iz[12][22] = 21'b000000000001000011110;
    W_iz[12][23] = 21'b000000000000100101100;
    W_iz[12][24] = 21'b111111111111001000001;
    W_iz[12][25] = 21'b111111111111010010111;
    W_iz[12][26] = 21'b000000000000000011101;
    W_iz[12][27] = 21'b111111111111001000001;
    W_iz[12][28] = 21'b000000000000101111101;
    W_iz[12][29] = 21'b111111111111111101101;
    W_iz[12][30] = 21'b000000000000101101100;
    W_iz[12][31] = 21'b111111111111100001001;
    W_iz[12][32] = 21'b111111111111001100000;
    W_iz[12][33] = 21'b111111111111010010101;
    W_iz[12][34] = 21'b111111111111100001100;
    W_iz[12][35] = 21'b111111111111011110111;
    W_iz[12][36] = 21'b111111111111001101101;
    W_iz[12][37] = 21'b111111111111010101011;
    W_iz[12][38] = 21'b111111111111100100100;
    W_iz[12][39] = 21'b000000000000010001010;
    W_iz[12][40] = 21'b000000000000001100000;
    W_iz[12][41] = 21'b111111111111100011001;
    W_iz[12][42] = 21'b111111111111111011111;
    W_iz[12][43] = 21'b111111111111101001111;
    W_iz[12][44] = 21'b111111111111000010010;
    W_iz[12][45] = 21'b111111111111110101100;
    W_iz[12][46] = 21'b111111111111110101010;
    W_iz[12][47] = 21'b111111111111111000011;
    W_iz[12][48] = 21'b000000000000000000001;
    W_iz[12][49] = 21'b111111111111110010100;
    W_iz[12][50] = 21'b000000000000101001110;
    W_iz[12][51] = 21'b111111111111100111000;
    W_iz[12][52] = 21'b000000000000111010100;
    W_iz[12][53] = 21'b000000000000011100010;
    W_iz[12][54] = 21'b000000000000111101100;
    W_iz[12][55] = 21'b000000000000110011011;
    W_iz[12][56] = 21'b000000000000010100001;
    W_iz[12][57] = 21'b111111111111001000100;
    W_iz[12][58] = 21'b000000000000100000111;
    W_iz[12][59] = 21'b000000000001101110110;
    W_iz[12][60] = 21'b000000000001010010110;
    W_iz[12][61] = 21'b000000000001010111011;
    W_iz[12][62] = 21'b000000000001100111001;
    W_iz[12][63] = 21'b000000000001011100000;
    W_iz[13][0] = 21'b000000000000001010100;
    W_iz[13][1] = 21'b000000000000001011011;
    W_iz[13][2] = 21'b000000000000001101011;
    W_iz[13][3] = 21'b111111111111111000010;
    W_iz[13][4] = 21'b111111111111110111011;
    W_iz[13][5] = 21'b111111111111011011000;
    W_iz[13][6] = 21'b000000000000110001111;
    W_iz[13][7] = 21'b111111111111000101010;
    W_iz[13][8] = 21'b111111111111010010100;
    W_iz[13][9] = 21'b111111111111101111011;
    W_iz[13][10] = 21'b111111111111111110101;
    W_iz[13][11] = 21'b111111111111110110101;
    W_iz[13][12] = 21'b111111111111011100001;
    W_iz[13][13] = 21'b111111111111110101100;
    W_iz[13][14] = 21'b111111111111100001000;
    W_iz[13][15] = 21'b111111111111011111111;
    W_iz[13][16] = 21'b000000000000100101000;
    W_iz[13][17] = 21'b111111111111010111110;
    W_iz[13][18] = 21'b000000000000000111110;
    W_iz[13][19] = 21'b111111111111001101111;
    W_iz[13][20] = 21'b111111111111110110000;
    W_iz[13][21] = 21'b000000000000000001011;
    W_iz[13][22] = 21'b000000000000010100101;
    W_iz[13][23] = 21'b000000000000001100111;
    W_iz[13][24] = 21'b111111111111111011000;
    W_iz[13][25] = 21'b111111111111100111101;
    W_iz[13][26] = 21'b111111111111111011010;
    W_iz[13][27] = 21'b000000000000010111010;
    W_iz[13][28] = 21'b000000000000000101000;
    W_iz[13][29] = 21'b111111111111100010100;
    W_iz[13][30] = 21'b111111111111110001000;
    W_iz[13][31] = 21'b111111111111001000100;
    W_iz[13][32] = 21'b111111111111111100011;
    W_iz[13][33] = 21'b111111111111000000001;
    W_iz[13][34] = 21'b111111111111101111111;
    W_iz[13][35] = 21'b000000000000011111001;
    W_iz[13][36] = 21'b111111111111100000100;
    W_iz[13][37] = 21'b111111111111010001001;
    W_iz[13][38] = 21'b111111111110111010011;
    W_iz[13][39] = 21'b000000000000101000111;
    W_iz[13][40] = 21'b111111111111101011101;
    W_iz[13][41] = 21'b111111111111111000000;
    W_iz[13][42] = 21'b000000000000000011011;
    W_iz[13][43] = 21'b111111111111101001100;
    W_iz[13][44] = 21'b000000000000001000010;
    W_iz[13][45] = 21'b111111111111101010100;
    W_iz[13][46] = 21'b111111111111110110110;
    W_iz[13][47] = 21'b000000000000011110100;
    W_iz[13][48] = 21'b000000000000001111010;
    W_iz[13][49] = 21'b000000000000001100100;
    W_iz[13][50] = 21'b000000000000001010101;
    W_iz[13][51] = 21'b000000000000001011001;
    W_iz[13][52] = 21'b111111111111101110110;
    W_iz[13][53] = 21'b111111111111101011100;
    W_iz[13][54] = 21'b000000000000001110101;
    W_iz[13][55] = 21'b000000000000000000001;
    W_iz[13][56] = 21'b000000000000001011000;
    W_iz[13][57] = 21'b111111111111011011111;
    W_iz[13][58] = 21'b111111111111011110011;
    W_iz[13][59] = 21'b111111111111101101100;
    W_iz[13][60] = 21'b000000000000111011101;
    W_iz[13][61] = 21'b000000000000101000100;
    W_iz[13][62] = 21'b111111111111101100000;
    W_iz[13][63] = 21'b000000000000100100010;
    W_iz[14][0] = 21'b000000000000101110101;
    W_iz[14][1] = 21'b111111111111110011101;
    W_iz[14][2] = 21'b000000000001001010111;
    W_iz[14][3] = 21'b111111111111101100111;
    W_iz[14][4] = 21'b000000000000101010000;
    W_iz[14][5] = 21'b000000000000001001111;
    W_iz[14][6] = 21'b111111111111001011000;
    W_iz[14][7] = 21'b000000000001001011000;
    W_iz[14][8] = 21'b000000000001010110010;
    W_iz[14][9] = 21'b000000000000110010101;
    W_iz[14][10] = 21'b000000000000111101101;
    W_iz[14][11] = 21'b111111111111111110100;
    W_iz[14][12] = 21'b000000000000000000111;
    W_iz[14][13] = 21'b000000000000010010101;
    W_iz[14][14] = 21'b111111111111101110000;
    W_iz[14][15] = 21'b111111111111001011100;
    W_iz[14][16] = 21'b111111111111101010010;
    W_iz[14][17] = 21'b000000000000100111011;
    W_iz[14][18] = 21'b111111111111111110101;
    W_iz[14][19] = 21'b111111111111111101001;
    W_iz[14][20] = 21'b111111111111110100011;
    W_iz[14][21] = 21'b111111111111010101011;
    W_iz[14][22] = 21'b000000000001000101100;
    W_iz[14][23] = 21'b111111111111111101100;
    W_iz[14][24] = 21'b111111111111010111010;
    W_iz[14][25] = 21'b000000000000010100001;
    W_iz[14][26] = 21'b111111111111010011110;
    W_iz[14][27] = 21'b111111111111011110000;
    W_iz[14][28] = 21'b000000000000110000111;
    W_iz[14][29] = 21'b000000000000101010010;
    W_iz[14][30] = 21'b111111111111010110000;
    W_iz[14][31] = 21'b000000000000100110100;
    W_iz[14][32] = 21'b000000000000000011011;
    W_iz[14][33] = 21'b000000000000010100010;
    W_iz[14][34] = 21'b000000000000110101101;
    W_iz[14][35] = 21'b000000000001000000010;
    W_iz[14][36] = 21'b111111111111111011001;
    W_iz[14][37] = 21'b000000000000001111101;
    W_iz[14][38] = 21'b111111111111000001011;
    W_iz[14][39] = 21'b111111111111111001101;
    W_iz[14][40] = 21'b000000000000011111111;
    W_iz[14][41] = 21'b111111111111100111100;
    W_iz[14][42] = 21'b000000000001000111000;
    W_iz[14][43] = 21'b000000000000010001000;
    W_iz[14][44] = 21'b000000000000100010001;
    W_iz[14][45] = 21'b111111111111100010100;
    W_iz[14][46] = 21'b111111111111001011101;
    W_iz[14][47] = 21'b000000000000111111111;
    W_iz[14][48] = 21'b111111111111010000001;
    W_iz[14][49] = 21'b111111111111100010010;
    W_iz[14][50] = 21'b000000000000100000010;
    W_iz[14][51] = 21'b111111111111111011011;
    W_iz[14][52] = 21'b000000000000100010000;
    W_iz[14][53] = 21'b111111111110010011000;
    W_iz[14][54] = 21'b111111111111110001011;
    W_iz[14][55] = 21'b000000000000001001101;
    W_iz[14][56] = 21'b111111111111011001011;
    W_iz[14][57] = 21'b111111111111101110001;
    W_iz[14][58] = 21'b111111111111010111000;
    W_iz[14][59] = 21'b111111111111010000100;
    W_iz[14][60] = 21'b111111111111110001011;
    W_iz[14][61] = 21'b111111111110011110000;
    W_iz[14][62] = 21'b111111111110001010000;
    W_iz[14][63] = 21'b111111111110000011000;
    W_iz[15][0] = 21'b111111111110101001010;
    W_iz[15][1] = 21'b111111111110100110001;
    W_iz[15][2] = 21'b000000000000011000111;
    W_iz[15][3] = 21'b111111111111110011001;
    W_iz[15][4] = 21'b000000000000110001101;
    W_iz[15][5] = 21'b000000000001000011110;
    W_iz[15][6] = 21'b111111111111001001011;
    W_iz[15][7] = 21'b000000000000001101000;
    W_iz[15][8] = 21'b111111111111010111011;
    W_iz[15][9] = 21'b111111111110011100101;
    W_iz[15][10] = 21'b111111111111011101111;
    W_iz[15][11] = 21'b000000000000100111101;
    W_iz[15][12] = 21'b000000000000101111110;
    W_iz[15][13] = 21'b111111111111010011011;
    W_iz[15][14] = 21'b000000000000110000100;
    W_iz[15][15] = 21'b111111111111111111111;
    W_iz[15][16] = 21'b000000000000001001111;
    W_iz[15][17] = 21'b111111111111101000000;
    W_iz[15][18] = 21'b000000000000001001110;
    W_iz[15][19] = 21'b000000000000111010110;
    W_iz[15][20] = 21'b111111111111100011111;
    W_iz[15][21] = 21'b111111111111101000101;
    W_iz[15][22] = 21'b000000000000111111011;
    W_iz[15][23] = 21'b111111111111100101010;
    W_iz[15][24] = 21'b000000000000111001000;
    W_iz[15][25] = 21'b000000000000011011100;
    W_iz[15][26] = 21'b000000000000100010101;
    W_iz[15][27] = 21'b111111111111110001110;
    W_iz[15][28] = 21'b000000000000101101010;
    W_iz[15][29] = 21'b000000000001000100010;
    W_iz[15][30] = 21'b000000000000101100101;
    W_iz[15][31] = 21'b000000000000011000000;
    W_iz[15][32] = 21'b111111111111010111010;
    W_iz[15][33] = 21'b111111111111100111011;
    W_iz[15][34] = 21'b111111111110100011110;
    W_iz[15][35] = 21'b111111111111001101001;
    W_iz[15][36] = 21'b000000000000111100101;
    W_iz[15][37] = 21'b000000000000000000100;
    W_iz[15][38] = 21'b000000000000110011010;
    W_iz[15][39] = 21'b111111111110111011111;
    W_iz[15][40] = 21'b111111111111111101110;
    W_iz[15][41] = 21'b111111111110111110000;
    W_iz[15][42] = 21'b111111111110111001101;
    W_iz[15][43] = 21'b111111111110110111000;
    W_iz[15][44] = 21'b111111111111011010100;
    W_iz[15][45] = 21'b000000000000001001101;
    W_iz[15][46] = 21'b000000000010001100001;
    W_iz[15][47] = 21'b111111111111011010011;
    W_iz[15][48] = 21'b111111111111111001110;
    W_iz[15][49] = 21'b111111111111010110100;
    W_iz[15][50] = 21'b111111111111000010100;
    W_iz[15][51] = 21'b000000000001011101100;
    W_iz[15][52] = 21'b111111111110111010011;
    W_iz[15][53] = 21'b000000000000010110001;
    W_iz[15][54] = 21'b000000000001000111000;
    W_iz[15][55] = 21'b000000000000001011010;
    W_iz[15][56] = 21'b000000000010010001011;
    W_iz[15][57] = 21'b000000000000010010011;
    W_iz[15][58] = 21'b000000000010010100011;
    W_iz[15][59] = 21'b000000000000010111101;
    W_iz[15][60] = 21'b111111111111000010100;
    W_iz[15][61] = 21'b000000000001000111000;
    W_iz[15][62] = 21'b000000000001100000011;
    W_iz[15][63] = 21'b111111111111000010100;

    // Initialize W_in weights
    W_in[0][0] = 21'b111111111111100011101;
    W_in[0][1] = 21'b000000000000001111100;
    W_in[0][2] = 21'b111111111111110011000;
    W_in[0][3] = 21'b000000000000100011100;
    W_in[0][4] = 21'b111111111111110110010;
    W_in[0][5] = 21'b111111111111101110011;
    W_in[0][6] = 21'b111111111111001000000;
    W_in[0][7] = 21'b111111111111100001101;
    W_in[0][8] = 21'b111111111111101110101;
    W_in[0][9] = 21'b000000000000100101101;
    W_in[0][10] = 21'b000000000000010001011;
    W_in[0][11] = 21'b000000000000110111100;
    W_in[0][12] = 21'b111111111111110001000;
    W_in[0][13] = 21'b000000000000011100110;
    W_in[0][14] = 21'b000000000000011100100;
    W_in[0][15] = 21'b000000000000001100001;
    W_in[0][16] = 21'b111111111111110101101;
    W_in[0][17] = 21'b000000000000101011101;
    W_in[0][18] = 21'b000000000000111111110;
    W_in[0][19] = 21'b000000000000100011100;
    W_in[0][20] = 21'b111111111111111001101;
    W_in[0][21] = 21'b000000000000001011110;
    W_in[0][22] = 21'b000000000000101100011;
    W_in[0][23] = 21'b000000000000001010000;
    W_in[0][24] = 21'b000000000000000011111;
    W_in[0][25] = 21'b111111111111110101001;
    W_in[0][26] = 21'b111111111111000100110;
    W_in[0][27] = 21'b000000000000001101100;
    W_in[0][28] = 21'b000000000000011111010;
    W_in[0][29] = 21'b000000000000000010110;
    W_in[0][30] = 21'b000000000000100111101;
    W_in[0][31] = 21'b000000000000100001111;
    W_in[0][32] = 21'b111111111111110110110;
    W_in[0][33] = 21'b111111111111011011111;
    W_in[0][34] = 21'b111111111111001110000;
    W_in[0][35] = 21'b111111111111100111011;
    W_in[0][36] = 21'b111111111111100100010;
    W_in[0][37] = 21'b111111111110101101001;
    W_in[0][38] = 21'b000000000000001110010;
    W_in[0][39] = 21'b111111111111111011100;
    W_in[0][40] = 21'b111111111111110100110;
    W_in[0][41] = 21'b000000000000110110110;
    W_in[0][42] = 21'b111111111111010101110;
    W_in[0][43] = 21'b000000000000100010110;
    W_in[0][44] = 21'b000000000000000000011;
    W_in[0][45] = 21'b111111111111100000100;
    W_in[0][46] = 21'b111111111111011010101;
    W_in[0][47] = 21'b000000000000101010111;
    W_in[0][48] = 21'b000000000000010001101;
    W_in[0][49] = 21'b000000000001001011101;
    W_in[0][50] = 21'b111111111111111111110;
    W_in[0][51] = 21'b000000000000001111011;
    W_in[0][52] = 21'b111111111111101101010;
    W_in[0][53] = 21'b111111111111010001111;
    W_in[0][54] = 21'b111111111111001011001;
    W_in[0][55] = 21'b111111111111100101110;
    W_in[0][56] = 21'b000000000000111011000;
    W_in[0][57] = 21'b111111111111101101010;
    W_in[0][58] = 21'b000000000000111100111;
    W_in[0][59] = 21'b111111111111110010001;
    W_in[0][60] = 21'b111111111110111010001;
    W_in[0][61] = 21'b111111111110010010000;
    W_in[0][62] = 21'b111111111110000000111;
    W_in[0][63] = 21'b000000000000011011111;
    W_in[1][0] = 21'b000000000000110010110;
    W_in[1][1] = 21'b000000000000010001101;
    W_in[1][2] = 21'b000000000000001011011;
    W_in[1][3] = 21'b000000000000000000110;
    W_in[1][4] = 21'b000000000000000111110;
    W_in[1][5] = 21'b000000000000100110100;
    W_in[1][6] = 21'b111111111111001101001;
    W_in[1][7] = 21'b111111111111010110100;
    W_in[1][8] = 21'b000000000000000001010;
    W_in[1][9] = 21'b000000000001000000100;
    W_in[1][10] = 21'b000000000000100001010;
    W_in[1][11] = 21'b111111111110111100101;
    W_in[1][12] = 21'b111111111111010111000;
    W_in[1][13] = 21'b000000000000101011100;
    W_in[1][14] = 21'b111111111111110010110;
    W_in[1][15] = 21'b000000000000110011010;
    W_in[1][16] = 21'b111111111111000011100;
    W_in[1][17] = 21'b000000000000011101101;
    W_in[1][18] = 21'b000000000001001000100;
    W_in[1][19] = 21'b111111111111010100010;
    W_in[1][20] = 21'b111111111111011001101;
    W_in[1][21] = 21'b111111111111000100001;
    W_in[1][22] = 21'b000000000000100011011;
    W_in[1][23] = 21'b000000000001010011111;
    W_in[1][24] = 21'b000000000000011111000;
    W_in[1][25] = 21'b111111111111100001011;
    W_in[1][26] = 21'b111111111111100110000;
    W_in[1][27] = 21'b111111111111011110110;
    W_in[1][28] = 21'b111111111111101010100;
    W_in[1][29] = 21'b111111111111001101100;
    W_in[1][30] = 21'b111111111111110001111;
    W_in[1][31] = 21'b111111111111001100111;
    W_in[1][32] = 21'b000000000000100111010;
    W_in[1][33] = 21'b111111111111101111101;
    W_in[1][34] = 21'b111111111111011111100;
    W_in[1][35] = 21'b000000000000101001011;
    W_in[1][36] = 21'b111111111110110110111;
    W_in[1][37] = 21'b000000000000001010100;
    W_in[1][38] = 21'b111111111111111110010;
    W_in[1][39] = 21'b111111111111011111100;
    W_in[1][40] = 21'b000000000000101101101;
    W_in[1][41] = 21'b000000000000010111000;
    W_in[1][42] = 21'b000000000000111011111;
    W_in[1][43] = 21'b000000000000110011011;
    W_in[1][44] = 21'b000000000000000011001;
    W_in[1][45] = 21'b000000000000111010101;
    W_in[1][46] = 21'b000000000000010000011;
    W_in[1][47] = 21'b111111111111110010011;
    W_in[1][48] = 21'b111111111111010001010;
    W_in[1][49] = 21'b111111111111110110110;
    W_in[1][50] = 21'b111111111111100101001;
    W_in[1][51] = 21'b000000000000011101001;
    W_in[1][52] = 21'b000000000000101011100;
    W_in[1][53] = 21'b000000000000011000100;
    W_in[1][54] = 21'b111111111111000011000;
    W_in[1][55] = 21'b000000000001001100110;
    W_in[1][56] = 21'b000000000000100110100;
    W_in[1][57] = 21'b111111111111110000101;
    W_in[1][58] = 21'b111111111111111011100;
    W_in[1][59] = 21'b000000000000110111110;
    W_in[1][60] = 21'b111111111110111011100;
    W_in[1][61] = 21'b111111111111111100110;
    W_in[1][62] = 21'b111111111111100100100;
    W_in[1][63] = 21'b111111111111101000000;
    W_in[2][0] = 21'b000000000000010110111;
    W_in[2][1] = 21'b000000000000011111101;
    W_in[2][2] = 21'b111111111111110100001;
    W_in[2][3] = 21'b000000000000001100011;
    W_in[2][4] = 21'b000000000000110011010;
    W_in[2][5] = 21'b000000000000010110010;
    W_in[2][6] = 21'b111111111110110110100;
    W_in[2][7] = 21'b000000000000010111001;
    W_in[2][8] = 21'b111111111110100000110;
    W_in[2][9] = 21'b111111111111110011010;
    W_in[2][10] = 21'b111111111111111110111;
    W_in[2][11] = 21'b111111111111100011111;
    W_in[2][12] = 21'b111111111111001000100;
    W_in[2][13] = 21'b000000000000011001010;
    W_in[2][14] = 21'b111111111111111100100;
    W_in[2][15] = 21'b111111111110101001101;
    W_in[2][16] = 21'b000000000000100001001;
    W_in[2][17] = 21'b000000000000100101001;
    W_in[2][18] = 21'b111111111110100001000;
    W_in[2][19] = 21'b111111111110111100111;
    W_in[2][20] = 21'b000000000000110100111;
    W_in[2][21] = 21'b111111111111001101111;
    W_in[2][22] = 21'b000000000000010101101;
    W_in[2][23] = 21'b111111111111010000011;
    W_in[2][24] = 21'b000000000000011001011;
    W_in[2][25] = 21'b111111111111010100111;
    W_in[2][26] = 21'b000000000001001010111;
    W_in[2][27] = 21'b111111111111110011111;
    W_in[2][28] = 21'b000000000000101101000;
    W_in[2][29] = 21'b000000000001000110111;
    W_in[2][30] = 21'b111111111111110110001;
    W_in[2][31] = 21'b000000000000000000010;
    W_in[2][32] = 21'b000000000001010111000;
    W_in[2][33] = 21'b111111111110111110100;
    W_in[2][34] = 21'b111111111111000010111;
    W_in[2][35] = 21'b111111111111100010110;
    W_in[2][36] = 21'b000000000001010000110;
    W_in[2][37] = 21'b000000000001000010111;
    W_in[2][38] = 21'b111111111111010110100;
    W_in[2][39] = 21'b111111111110101011101;
    W_in[2][40] = 21'b000000000000100011100;
    W_in[2][41] = 21'b111111111111111011010;
    W_in[2][42] = 21'b111111111111000011101;
    W_in[2][43] = 21'b000000000000001011001;
    W_in[2][44] = 21'b111111111111101011011;
    W_in[2][45] = 21'b000000000000100110100;
    W_in[2][46] = 21'b111111111111110001110;
    W_in[2][47] = 21'b111111111111110001100;
    W_in[2][48] = 21'b111111111111100111111;
    W_in[2][49] = 21'b111111111111111111001;
    W_in[2][50] = 21'b111111111111000011100;
    W_in[2][51] = 21'b111111111111100110101;
    W_in[2][52] = 21'b111111111110111111000;
    W_in[2][53] = 21'b000000000000110110101;
    W_in[2][54] = 21'b111111111111111000000;
    W_in[2][55] = 21'b111111111111100011100;
    W_in[2][56] = 21'b111111111111100100101;
    W_in[2][57] = 21'b000000000000111001101;
    W_in[2][58] = 21'b000000000000111101110;
    W_in[2][59] = 21'b000000000001001101101;
    W_in[2][60] = 21'b000000000001111001011;
    W_in[2][61] = 21'b000000000001010001011;
    W_in[2][62] = 21'b000000000010001011110;
    W_in[2][63] = 21'b000000000001100111101;
    W_in[3][0] = 21'b111111111110100110010;
    W_in[3][1] = 21'b000000000001000001011;
    W_in[3][2] = 21'b000000000000000100111;
    W_in[3][3] = 21'b000000000001000111000;
    W_in[3][4] = 21'b111111111110101110010;
    W_in[3][5] = 21'b000000000000010001101;
    W_in[3][6] = 21'b111111111110111000010;
    W_in[3][7] = 21'b000000000000100111101;
    W_in[3][8] = 21'b111111111110010001110;
    W_in[3][9] = 21'b111111111110100110000;
    W_in[3][10] = 21'b000000000001001010001;
    W_in[3][11] = 21'b111111111110100110001;
    W_in[3][12] = 21'b111111111110101000111;
    W_in[3][13] = 21'b000000000000100101001;
    W_in[3][14] = 21'b000000000000011111101;
    W_in[3][15] = 21'b000000000000011111110;
    W_in[3][16] = 21'b000000000001010101001;
    W_in[3][17] = 21'b111111111111101110010;
    W_in[3][18] = 21'b111111111111111111101;
    W_in[3][19] = 21'b000000000001100101100;
    W_in[3][20] = 21'b111111111111110000100;
    W_in[3][21] = 21'b111111111111000011100;
    W_in[3][22] = 21'b111111111111101001011;
    W_in[3][23] = 21'b111111111111100010111;
    W_in[3][24] = 21'b111111111110110000110;
    W_in[3][25] = 21'b111111111111110001011;
    W_in[3][26] = 21'b111111111110111111011;
    W_in[3][27] = 21'b111111111110101111111;
    W_in[3][28] = 21'b000000000001101001110;
    W_in[3][29] = 21'b000000000000100011011;
    W_in[3][30] = 21'b000000000000000110011;
    W_in[3][31] = 21'b000000000000111010101;
    W_in[3][32] = 21'b000000000000100010100;
    W_in[3][33] = 21'b111111111111110000001;
    W_in[3][34] = 21'b000000000000111001010;
    W_in[3][35] = 21'b000000000000011100110;
    W_in[3][36] = 21'b111111111110111011110;
    W_in[3][37] = 21'b111111111110101101110;
    W_in[3][38] = 21'b000000000000100010011;
    W_in[3][39] = 21'b111111111111111101010;
    W_in[3][40] = 21'b111111111110100000101;
    W_in[3][41] = 21'b111111111110101100110;
    W_in[3][42] = 21'b000000000001000001011;
    W_in[3][43] = 21'b000000000000000101111;
    W_in[3][44] = 21'b000000000000010110001;
    W_in[3][45] = 21'b000000000001100011100;
    W_in[3][46] = 21'b111111111111110111000;
    W_in[3][47] = 21'b000000000001010000001;
    W_in[3][48] = 21'b000000000000001001100;
    W_in[3][49] = 21'b111111111111110110110;
    W_in[3][50] = 21'b111111111111010100111;
    W_in[3][51] = 21'b000000000000101100110;
    W_in[3][52] = 21'b111111111111101100001;
    W_in[3][53] = 21'b111111111110101111001;
    W_in[3][54] = 21'b000000000001100010010;
    W_in[3][55] = 21'b000000000000001111001;
    W_in[3][56] = 21'b111111111111010001101;
    W_in[3][57] = 21'b000000000000101101100;
    W_in[3][58] = 21'b111111111111011001111;
    W_in[3][59] = 21'b000000000001011000101;
    W_in[3][60] = 21'b000000000001010111010;
    W_in[3][61] = 21'b000000000000010100110;
    W_in[3][62] = 21'b000000000000000111001;
    W_in[3][63] = 21'b000000000001001011111;
    W_in[4][0] = 21'b000000000000010100101;
    W_in[4][1] = 21'b000000000000100111001;
    W_in[4][2] = 21'b000000000000011101110;
    W_in[4][3] = 21'b000000000000100011010;
    W_in[4][4] = 21'b111111111111101101010;
    W_in[4][5] = 21'b111111111111010101010;
    W_in[4][6] = 21'b000000000000011100111;
    W_in[4][7] = 21'b000000000000001111011;
    W_in[4][8] = 21'b111111111111001000001;
    W_in[4][9] = 21'b000000000000000101101;
    W_in[4][10] = 21'b000000000000111110110;
    W_in[4][11] = 21'b111111111111111111101;
    W_in[4][12] = 21'b000000000000101000000;
    W_in[4][13] = 21'b000000000000001011000;
    W_in[4][14] = 21'b000000000000001001111;
    W_in[4][15] = 21'b000000000000101110011;
    W_in[4][16] = 21'b111111111111111000000;
    W_in[4][17] = 21'b000000000000110111010;
    W_in[4][18] = 21'b111111111111111000110;
    W_in[4][19] = 21'b000000000000100100010;
    W_in[4][20] = 21'b111111111111111000100;
    W_in[4][21] = 21'b000000000000100001110;
    W_in[4][22] = 21'b000000000000011000100;
    W_in[4][23] = 21'b000000000000011000111;
    W_in[4][24] = 21'b111111111111010111110;
    W_in[4][25] = 21'b000000000000011110000;
    W_in[4][26] = 21'b000000000000100010111;
    W_in[4][27] = 21'b000000000000010110111;
    W_in[4][28] = 21'b000000000000111000101;
    W_in[4][29] = 21'b111111111111001011000;
    W_in[4][30] = 21'b111111111111101101011;
    W_in[4][31] = 21'b000000000000011001110;
    W_in[4][32] = 21'b000000000000001100011;
    W_in[4][33] = 21'b000000000000011110100;
    W_in[4][34] = 21'b000000000000011110101;
    W_in[4][35] = 21'b000000000000000110110;
    W_in[4][36] = 21'b000000000000111111101;
    W_in[4][37] = 21'b000000000000010100010;
    W_in[4][38] = 21'b111111111111101110110;
    W_in[4][39] = 21'b000000000000001111011;
    W_in[4][40] = 21'b000000000000100101011;
    W_in[4][41] = 21'b111111111111010000010;
    W_in[4][42] = 21'b000000000000001111010;
    W_in[4][43] = 21'b111111111111101000010;
    W_in[4][44] = 21'b111111111111111110010;
    W_in[4][45] = 21'b111111111111011100101;
    W_in[4][46] = 21'b111111111111001110100;
    W_in[4][47] = 21'b000000000000110111101;
    W_in[4][48] = 21'b111111111111110001010;
    W_in[4][49] = 21'b111111111111100111001;
    W_in[4][50] = 21'b111111111111111001101;
    W_in[4][51] = 21'b000000000000000000010;
    W_in[4][52] = 21'b111111111111000110110;
    W_in[4][53] = 21'b111111111111101010010;
    W_in[4][54] = 21'b000000000000010000110;
    W_in[4][55] = 21'b111111111111100111110;
    W_in[4][56] = 21'b000000000000100110010;
    W_in[4][57] = 21'b111111111111100101011;
    W_in[4][58] = 21'b111111111111101011011;
    W_in[4][59] = 21'b000000000000100010000;
    W_in[4][60] = 21'b111111111111010101000;
    W_in[4][61] = 21'b111111111111001101111;
    W_in[4][62] = 21'b111111111111001100100;
    W_in[4][63] = 21'b000000000000100001100;
    W_in[5][0] = 21'b111111111111100010111;
    W_in[5][1] = 21'b111111111111100110011;
    W_in[5][2] = 21'b000000000000101111111;
    W_in[5][3] = 21'b000000000000100101101;
    W_in[5][4] = 21'b000000000000000101001;
    W_in[5][5] = 21'b000000000000001111100;
    W_in[5][6] = 21'b000000000000001101001;
    W_in[5][7] = 21'b000000000000001000010;
    W_in[5][8] = 21'b000000000000001010000;
    W_in[5][9] = 21'b000000000000001001010;
    W_in[5][10] = 21'b111111111111111000100;
    W_in[5][11] = 21'b111111111111111111110;
    W_in[5][12] = 21'b000000000000001011101;
    W_in[5][13] = 21'b000000000000011100000;
    W_in[5][14] = 21'b111111111111010101101;
    W_in[5][15] = 21'b000000000000001000100;
    W_in[5][16] = 21'b111111111111111111111;
    W_in[5][17] = 21'b111111111111111111001;
    W_in[5][18] = 21'b111111111111111100100;
    W_in[5][19] = 21'b111111111111101100000;
    W_in[5][20] = 21'b111111111111111100000;
    W_in[5][21] = 21'b000000000000001011011;
    W_in[5][22] = 21'b111111111111110000000;
    W_in[5][23] = 21'b111111111111101000000;
    W_in[5][24] = 21'b000000000000000000011;
    W_in[5][25] = 21'b000000000000101110101;
    W_in[5][26] = 21'b111111111111001100101;
    W_in[5][27] = 21'b111111111111001110101;
    W_in[5][28] = 21'b000000000000110101101;
    W_in[5][29] = 21'b000000000000010000010;
    W_in[5][30] = 21'b000000000000000011101;
    W_in[5][31] = 21'b111111111111111111011;
    W_in[5][32] = 21'b111111111111100001010;
    W_in[5][33] = 21'b111111111111111101001;
    W_in[5][34] = 21'b111111111111111011010;
    W_in[5][35] = 21'b000000000000000011110;
    W_in[5][36] = 21'b000000000000001111110;
    W_in[5][37] = 21'b000000000000001001001;
    W_in[5][38] = 21'b000000000000001100101;
    W_in[5][39] = 21'b000000000000100000001;
    W_in[5][40] = 21'b000000000000010011010;
    W_in[5][41] = 21'b000000000000000000011;
    W_in[5][42] = 21'b111111111111111101010;
    W_in[5][43] = 21'b000000000000010000010;
    W_in[5][44] = 21'b000000000000000110001;
    W_in[5][45] = 21'b000000000000001100101;
    W_in[5][46] = 21'b111111111111111100111;
    W_in[5][47] = 21'b111111111111110111001;
    W_in[5][48] = 21'b111111111111110110111;
    W_in[5][49] = 21'b111111111111001010111;
    W_in[5][50] = 21'b000000000000011110101;
    W_in[5][51] = 21'b000000000000101010101;
    W_in[5][52] = 21'b111111111111110011100;
    W_in[5][53] = 21'b111111111111100111011;
    W_in[5][54] = 21'b111111111111101000000;
    W_in[5][55] = 21'b111111111111100100111;
    W_in[5][56] = 21'b111111111111110000011;
    W_in[5][57] = 21'b000000000000110010111;
    W_in[5][58] = 21'b000000000000011101110;
    W_in[5][59] = 21'b111111111111011111001;
    W_in[5][60] = 21'b111111111111110111101;
    W_in[5][61] = 21'b111111111111110010011;
    W_in[5][62] = 21'b000000000000101011000;
    W_in[5][63] = 21'b111111111111100111110;
    W_in[6][0] = 21'b111111111111101001001;
    W_in[6][1] = 21'b111111111111110000001;
    W_in[6][2] = 21'b111111111111001001100;
    W_in[6][3] = 21'b111111111111011110010;
    W_in[6][4] = 21'b111111111111101101011;
    W_in[6][5] = 21'b111111111111110111011;
    W_in[6][6] = 21'b000000000000000101111;
    W_in[6][7] = 21'b111111111111010111011;
    W_in[6][8] = 21'b111111111111110101000;
    W_in[6][9] = 21'b111111111111110101100;
    W_in[6][10] = 21'b111111111111110100001;
    W_in[6][11] = 21'b111111111111000101101;
    W_in[6][12] = 21'b111111111111110110110;
    W_in[6][13] = 21'b000000000000001101111;
    W_in[6][14] = 21'b111111111111110101000;
    W_in[6][15] = 21'b000000000000010110000;
    W_in[6][16] = 21'b111111111111010110100;
    W_in[6][17] = 21'b000000000000111001011;
    W_in[6][18] = 21'b000000000000000011000;
    W_in[6][19] = 21'b000000000000010011000;
    W_in[6][20] = 21'b000000000000001101111;
    W_in[6][21] = 21'b111111111111101110000;
    W_in[6][22] = 21'b000000000000011110000;
    W_in[6][23] = 21'b000000000000110101000;
    W_in[6][24] = 21'b000000000000011011000;
    W_in[6][25] = 21'b000000000000001000111;
    W_in[6][26] = 21'b111111111111111100000;
    W_in[6][27] = 21'b111111111111001011011;
    W_in[6][28] = 21'b111111111111110001000;
    W_in[6][29] = 21'b000000000000111100011;
    W_in[6][30] = 21'b111111111111101000000;
    W_in[6][31] = 21'b111111111111101000010;
    W_in[6][32] = 21'b000000000000000010110;
    W_in[6][33] = 21'b000000000000010111000;
    W_in[6][34] = 21'b111111111111110100010;
    W_in[6][35] = 21'b111111111111110010100;
    W_in[6][36] = 21'b000000000000000011000;
    W_in[6][37] = 21'b000000000000001010101;
    W_in[6][38] = 21'b000000000000100000000;
    W_in[6][39] = 21'b111111111111111111101;
    W_in[6][40] = 21'b000000000000011100100;
    W_in[6][41] = 21'b111111111111110010101;
    W_in[6][42] = 21'b000000000000011101101;
    W_in[6][43] = 21'b111111111111111100110;
    W_in[6][44] = 21'b000000000000001011010;
    W_in[6][45] = 21'b000000000000001111111;
    W_in[6][46] = 21'b000000000000001100100;
    W_in[6][47] = 21'b000000000000000110100;
    W_in[6][48] = 21'b000000000000001100111;
    W_in[6][49] = 21'b000000000000001010111;
    W_in[6][50] = 21'b111111111111100001100;
    W_in[6][51] = 21'b000000000000010101110;
    W_in[6][52] = 21'b000000000000010100100;
    W_in[6][53] = 21'b000000000000001110010;
    W_in[6][54] = 21'b111111111111001001010;
    W_in[6][55] = 21'b000000000000010010110;
    W_in[6][56] = 21'b000000000000001100100;
    W_in[6][57] = 21'b111111111111010111010;
    W_in[6][58] = 21'b111111111111100001111;
    W_in[6][59] = 21'b111111111111100101101;
    W_in[6][60] = 21'b000000000000100110011;
    W_in[6][61] = 21'b000000000000010001100;
    W_in[6][62] = 21'b000000000000100111110;
    W_in[6][63] = 21'b000000000001000110101;
    W_in[7][0] = 21'b111111111111111101111;
    W_in[7][1] = 21'b000000000000111111011;
    W_in[7][2] = 21'b000000000000000000001;
    W_in[7][3] = 21'b000000000000110010101;
    W_in[7][4] = 21'b111111111111010010000;
    W_in[7][5] = 21'b000000000000001010011;
    W_in[7][6] = 21'b000000000000000111101;
    W_in[7][7] = 21'b111111111111101100111;
    W_in[7][8] = 21'b111111111111111000110;
    W_in[7][9] = 21'b000000000000101001101;
    W_in[7][10] = 21'b111111111111100010011;
    W_in[7][11] = 21'b111111111111111010100;
    W_in[7][12] = 21'b111111111111011111101;
    W_in[7][13] = 21'b111111111111110101001;
    W_in[7][14] = 21'b111111111111110001111;
    W_in[7][15] = 21'b111111111111111000110;
    W_in[7][16] = 21'b000000000000000010011;
    W_in[7][17] = 21'b000000000000001010110;
    W_in[7][18] = 21'b111111111111101001110;
    W_in[7][19] = 21'b000000000000100000100;
    W_in[7][20] = 21'b111111111111110011000;
    W_in[7][21] = 21'b000000000000001100111;
    W_in[7][22] = 21'b000000000000010101001;
    W_in[7][23] = 21'b000000000000001101101;
    W_in[7][24] = 21'b000000000000110101001;
    W_in[7][25] = 21'b000000000000001011101;
    W_in[7][26] = 21'b111111111111111000100;
    W_in[7][27] = 21'b111111111111101100101;
    W_in[7][28] = 21'b000000000000001011011;
    W_in[7][29] = 21'b000000000000001001100;
    W_in[7][30] = 21'b111111111111011110000;
    W_in[7][31] = 21'b000000000001000010010;
    W_in[7][32] = 21'b000000000000100010000;
    W_in[7][33] = 21'b111111111111011000101;
    W_in[7][34] = 21'b000000000000010000000;
    W_in[7][35] = 21'b000000000000001001010;
    W_in[7][36] = 21'b000000000000001011110;
    W_in[7][37] = 21'b111111111111000111111;
    W_in[7][38] = 21'b000000000000011000100;
    W_in[7][39] = 21'b000000000000000011101;
    W_in[7][40] = 21'b111111111111111110111;
    W_in[7][41] = 21'b000000000000100101011;
    W_in[7][42] = 21'b111111111111010110010;
    W_in[7][43] = 21'b000000000000000110000;
    W_in[7][44] = 21'b111111111111101010000;
    W_in[7][45] = 21'b111111111111101110001;
    W_in[7][46] = 21'b000000000000110001100;
    W_in[7][47] = 21'b111111111111101000111;
    W_in[7][48] = 21'b111111111111110010100;
    W_in[7][49] = 21'b111111111111110110011;
    W_in[7][50] = 21'b111111111111100100000;
    W_in[7][51] = 21'b111111111111101000001;
    W_in[7][52] = 21'b111111111111100101111;
    W_in[7][53] = 21'b111111111111100010111;
    W_in[7][54] = 21'b111111111111101111011;
    W_in[7][55] = 21'b111111111111000110000;
    W_in[7][56] = 21'b111111111111100100110;
    W_in[7][57] = 21'b000000000000011111010;
    W_in[7][58] = 21'b111111111111011100111;
    W_in[7][59] = 21'b111111111111100111001;
    W_in[7][60] = 21'b111111111111101000000;
    W_in[7][61] = 21'b111111111111101011011;
    W_in[7][62] = 21'b111111111111010000010;
    W_in[7][63] = 21'b111111111111101100000;
    W_in[8][0] = 21'b111111111111111100100;
    W_in[8][1] = 21'b111111111111110011011;
    W_in[8][2] = 21'b111111111111110110110;
    W_in[8][3] = 21'b111111111111100111010;
    W_in[8][4] = 21'b000000000000000001010;
    W_in[8][5] = 21'b000000000000010111001;
    W_in[8][6] = 21'b111111111111100011011;
    W_in[8][7] = 21'b111111111111010111010;
    W_in[8][8] = 21'b111111111111000101000;
    W_in[8][9] = 21'b111111111111101001011;
    W_in[8][10] = 21'b111111111111001011100;
    W_in[8][11] = 21'b111111111111101111000;
    W_in[8][12] = 21'b111111111111110110101;
    W_in[8][13] = 21'b000000000000010111000;
    W_in[8][14] = 21'b000000000000000110010;
    W_in[8][15] = 21'b111111111111110110101;
    W_in[8][16] = 21'b111111111111100000110;
    W_in[8][17] = 21'b111111111111101000101;
    W_in[8][18] = 21'b111111111111100001101;
    W_in[8][19] = 21'b111111111111011010101;
    W_in[8][20] = 21'b111111111111110111001;
    W_in[8][21] = 21'b000000000000011010110;
    W_in[8][22] = 21'b000000000001000011110;
    W_in[8][23] = 21'b000000000000100101100;
    W_in[8][24] = 21'b111111111111001000001;
    W_in[8][25] = 21'b111111111111010010111;
    W_in[8][26] = 21'b000000000000000011101;
    W_in[8][27] = 21'b111111111111001000001;
    W_in[8][28] = 21'b000000000000101111101;
    W_in[8][29] = 21'b111111111111111101101;
    W_in[8][30] = 21'b000000000000101101100;
    W_in[8][31] = 21'b111111111111100001001;
    W_in[8][32] = 21'b111111111111001100000;
    W_in[8][33] = 21'b111111111111010010101;
    W_in[8][34] = 21'b111111111111100001100;
    W_in[8][35] = 21'b111111111111011110111;
    W_in[8][36] = 21'b111111111111001101101;
    W_in[8][37] = 21'b111111111111010101011;
    W_in[8][38] = 21'b111111111111100100100;
    W_in[8][39] = 21'b000000000000010001010;
    W_in[8][40] = 21'b000000000000001100000;
    W_in[8][41] = 21'b111111111111100011001;
    W_in[8][42] = 21'b111111111111111011111;
    W_in[8][43] = 21'b111111111111101001111;
    W_in[8][44] = 21'b111111111111000010010;
    W_in[8][45] = 21'b111111111111110101100;
    W_in[8][46] = 21'b111111111111110101010;
    W_in[8][47] = 21'b111111111111111000011;
    W_in[8][48] = 21'b000000000000000000001;
    W_in[8][49] = 21'b111111111111110010100;
    W_in[8][50] = 21'b000000000000101001110;
    W_in[8][51] = 21'b111111111111100111000;
    W_in[8][52] = 21'b000000000000111010100;
    W_in[8][53] = 21'b000000000000011100010;
    W_in[8][54] = 21'b000000000000111101100;
    W_in[8][55] = 21'b000000000000110011011;
    W_in[8][56] = 21'b000000000000010100001;
    W_in[8][57] = 21'b111111111111001000100;
    W_in[8][58] = 21'b000000000000100000111;
    W_in[8][59] = 21'b000000000001101110110;
    W_in[8][60] = 21'b000000000001010010110;
    W_in[8][61] = 21'b000000000001010111011;
    W_in[8][62] = 21'b000000000001100111001;
    W_in[8][63] = 21'b000000000001011100000;
    W_in[9][0] = 21'b000000000000001010100;
    W_in[9][1] = 21'b000000000000001011011;
    W_in[9][2] = 21'b000000000000001101011;
    W_in[9][3] = 21'b111111111111111000010;
    W_in[9][4] = 21'b111111111111110111011;
    W_in[9][5] = 21'b111111111111011011000;
    W_in[9][6] = 21'b000000000000110001111;
    W_in[9][7] = 21'b111111111111000101010;
    W_in[9][8] = 21'b111111111111010010100;
    W_in[9][9] = 21'b111111111111101111011;
    W_in[9][10] = 21'b111111111111111110101;
    W_in[9][11] = 21'b111111111111110110101;
    W_in[9][12] = 21'b111111111111011100001;
    W_in[9][13] = 21'b111111111111110101100;
    W_in[9][14] = 21'b111111111111100001000;
    W_in[9][15] = 21'b111111111111011111111;
    W_in[9][16] = 21'b000000000000100101000;
    W_in[9][17] = 21'b111111111111010111110;
    W_in[9][18] = 21'b000000000000000111110;
    W_in[9][19] = 21'b111111111111001101111;
    W_in[9][20] = 21'b111111111111110110000;
    W_in[9][21] = 21'b000000000000000001011;
    W_in[9][22] = 21'b000000000000010100101;
    W_in[9][23] = 21'b000000000000001100111;
    W_in[9][24] = 21'b111111111111111011000;
    W_in[9][25] = 21'b111111111111100111101;
    W_in[9][26] = 21'b111111111111111011010;
    W_in[9][27] = 21'b000000000000010111010;
    W_in[9][28] = 21'b000000000000000101000;
    W_in[9][29] = 21'b111111111111100010100;
    W_in[9][30] = 21'b111111111111110001000;
    W_in[9][31] = 21'b111111111111001000100;
    W_in[9][32] = 21'b111111111111111100011;
    W_in[9][33] = 21'b111111111111000000001;
    W_in[9][34] = 21'b111111111111101111111;
    W_in[9][35] = 21'b000000000000011111001;
    W_in[9][36] = 21'b111111111111100000100;
    W_in[9][37] = 21'b111111111111010001001;
    W_in[9][38] = 21'b111111111110111010011;
    W_in[9][39] = 21'b000000000000101000111;
    W_in[9][40] = 21'b111111111111101011101;
    W_in[9][41] = 21'b111111111111111000000;
    W_in[9][42] = 21'b000000000000000011011;
    W_in[9][43] = 21'b111111111111101001100;
    W_in[9][44] = 21'b000000000000001000010;
    W_in[9][45] = 21'b111111111111101010100;
    W_in[9][46] = 21'b111111111111110110110;
    W_in[9][47] = 21'b000000000000011110100;
    W_in[9][48] = 21'b000000000000001111010;
    W_in[9][49] = 21'b000000000000001100100;
    W_in[9][50] = 21'b000000000000001010101;
    W_in[9][51] = 21'b000000000000001011001;
    W_in[9][52] = 21'b111111111111101110110;
    W_in[9][53] = 21'b111111111111101011100;
    W_in[9][54] = 21'b000000000000001110101;
    W_in[9][55] = 21'b000000000000000000001;
    W_in[9][56] = 21'b000000000000001011000;
    W_in[9][57] = 21'b111111111111011011111;
    W_in[9][58] = 21'b111111111111011110011;
    W_in[9][59] = 21'b111111111111101101100;
    W_in[9][60] = 21'b000000000000111011101;
    W_in[9][61] = 21'b000000000000101000100;
    W_in[9][62] = 21'b111111111111101100000;
    W_in[9][63] = 21'b000000000000100100010;
    W_in[10][0] = 21'b000000000000101110101;
    W_in[10][1] = 21'b111111111111110011101;
    W_in[10][2] = 21'b000000000001001010111;
    W_in[10][3] = 21'b111111111111101100111;
    W_in[10][4] = 21'b000000000000101010000;
    W_in[10][5] = 21'b000000000000001001111;
    W_in[10][6] = 21'b111111111111001011000;
    W_in[10][7] = 21'b000000000001001011000;
    W_in[10][8] = 21'b000000000001010110010;
    W_in[10][9] = 21'b000000000000110010101;
    W_in[10][10] = 21'b000000000000111101101;
    W_in[10][11] = 21'b111111111111111110100;
    W_in[10][12] = 21'b000000000000000000111;
    W_in[10][13] = 21'b000000000000010010101;
    W_in[10][14] = 21'b111111111111101110000;
    W_in[10][15] = 21'b111111111111001011100;
    W_in[10][16] = 21'b111111111111101010010;
    W_in[10][17] = 21'b000000000000100111011;
    W_in[10][18] = 21'b111111111111111110101;
    W_in[10][19] = 21'b111111111111111101001;
    W_in[10][20] = 21'b111111111111110100011;
    W_in[10][21] = 21'b111111111111010101011;
    W_in[10][22] = 21'b000000000001000101100;
    W_in[10][23] = 21'b111111111111111101100;
    W_in[10][24] = 21'b111111111111010111010;
    W_in[10][25] = 21'b000000000000010100001;
    W_in[10][26] = 21'b111111111111010011110;
    W_in[10][27] = 21'b111111111111011110000;
    W_in[10][28] = 21'b000000000000110000111;
    W_in[10][29] = 21'b000000000000101010010;
    W_in[10][30] = 21'b111111111111010110000;
    W_in[10][31] = 21'b000000000000100110100;
    W_in[10][32] = 21'b000000000000000011011;
    W_in[10][33] = 21'b000000000000010100010;
    W_in[10][34] = 21'b000000000000110101101;
    W_in[10][35] = 21'b000000000001000000010;
    W_in[10][36] = 21'b111111111111111011001;
    W_in[10][37] = 21'b000000000000001111101;
    W_in[10][38] = 21'b111111111111000001011;
    W_in[10][39] = 21'b111111111111111001101;
    W_in[10][40] = 21'b000000000000011111111;
    W_in[10][41] = 21'b111111111111100111100;
    W_in[10][42] = 21'b000000000001000111000;
    W_in[10][43] = 21'b000000000000010001000;
    W_in[10][44] = 21'b000000000000100010001;
    W_in[10][45] = 21'b111111111111100010100;
    W_in[10][46] = 21'b111111111111001011101;
    W_in[10][47] = 21'b000000000000111111111;
    W_in[10][48] = 21'b111111111111010000001;
    W_in[10][49] = 21'b111111111111100010010;
    W_in[10][50] = 21'b000000000000100000010;
    W_in[10][51] = 21'b111111111111111011011;
    W_in[10][52] = 21'b000000000000100010000;
    W_in[10][53] = 21'b111111111110010011000;
    W_in[10][54] = 21'b111111111111110001011;
    W_in[10][55] = 21'b000000000000001001101;
    W_in[10][56] = 21'b111111111111011001011;
    W_in[10][57] = 21'b111111111111101110001;
    W_in[10][58] = 21'b111111111111010111000;
    W_in[10][59] = 21'b111111111111010000100;
    W_in[10][60] = 21'b111111111111110001011;
    W_in[10][61] = 21'b111111111110011110000;
    W_in[10][62] = 21'b111111111110001010000;
    W_in[10][63] = 21'b111111111110000011000;
    W_in[11][0] = 21'b111111111110101001010;
    W_in[11][1] = 21'b111111111110100110001;
    W_in[11][2] = 21'b000000000000011000111;
    W_in[11][3] = 21'b111111111111110011001;
    W_in[11][4] = 21'b000000000000110001101;
    W_in[11][5] = 21'b000000000001000011110;
    W_in[11][6] = 21'b111111111111001001011;
    W_in[11][7] = 21'b000000000000001101000;
    W_in[11][8] = 21'b111111111111010111011;
    W_in[11][9] = 21'b111111111110011100101;
    W_in[11][10] = 21'b111111111111011101111;
    W_in[11][11] = 21'b000000000000100111101;
    W_in[11][12] = 21'b000000000000101111110;
    W_in[11][13] = 21'b111111111111010011011;
    W_in[11][14] = 21'b000000000000110000100;
    W_in[11][15] = 21'b111111111111111111111;
    W_in[11][16] = 21'b000000000000001001111;
    W_in[11][17] = 21'b111111111111101000000;
    W_in[11][18] = 21'b000000000000001001110;
    W_in[11][19] = 21'b000000000000111010110;
    W_in[11][20] = 21'b111111111111100011111;
    W_in[11][21] = 21'b111111111111101000101;
    W_in[11][22] = 21'b000000000000111111011;
    W_in[11][23] = 21'b111111111111100101010;
    W_in[11][24] = 21'b000000000000111001000;
    W_in[11][25] = 21'b000000000000011011100;
    W_in[11][26] = 21'b000000000000100010101;
    W_in[11][27] = 21'b111111111111110001110;
    W_in[11][28] = 21'b000000000000101101010;
    W_in[11][29] = 21'b000000000001000100010;
    W_in[11][30] = 21'b000000000000101100101;
    W_in[11][31] = 21'b000000000000011000000;
    W_in[11][32] = 21'b111111111111010111010;
    W_in[11][33] = 21'b111111111111100111011;
    W_in[11][34] = 21'b111111111110100011110;
    W_in[11][35] = 21'b111111111111001101001;
    W_in[11][36] = 21'b000000000000111100101;
    W_in[11][37] = 21'b000000000000000000100;
    W_in[11][38] = 21'b000000000000110011010;
    W_in[11][39] = 21'b111111111110111011111;
    W_in[11][40] = 21'b111111111111111101110;
    W_in[11][41] = 21'b111111111110111110000;
    W_in[11][42] = 21'b111111111110111001101;
    W_in[11][43] = 21'b111111111110110111000;
    W_in[11][44] = 21'b111111111111011010100;
    W_in[11][45] = 21'b000000000000001001101;
    W_in[11][46] = 21'b000000000010001100001;
    W_in[11][47] = 21'b111111111111011010011;
    W_in[11][48] = 21'b111111111111111001110;
    W_in[11][49] = 21'b111111111111010110100;
    W_in[11][50] = 21'b111111111111000010100;
    W_in[11][51] = 21'b000000000001011101100;
    W_in[11][52] = 21'b111111111110111010011;
    W_in[11][53] = 21'b000000000000010110001;
    W_in[11][54] = 21'b000000000001000111000;
    W_in[11][55] = 21'b000000000000001011010;
    W_in[11][56] = 21'b000000000010010001011;
    W_in[11][57] = 21'b000000000000010010011;
    W_in[11][58] = 21'b000000000010010100011;
    W_in[11][59] = 21'b000000000000010111101;
    W_in[11][60] = 21'b111111111111000010100;
    W_in[11][61] = 21'b000000000001000111000;
    W_in[11][62] = 21'b000000000001100000011;
    W_in[11][63] = 21'b111111111111000010100;
    W_in[12][0] = 21'b111111111111100011101;
    W_in[12][1] = 21'b000000000000001111100;
    W_in[12][2] = 21'b111111111111110011000;
    W_in[12][3] = 21'b000000000000100011100;
    W_in[12][4] = 21'b111111111111110110010;
    W_in[12][5] = 21'b111111111111101110011;
    W_in[12][6] = 21'b111111111111001000000;
    W_in[12][7] = 21'b111111111111100001101;
    W_in[12][8] = 21'b111111111111101110101;
    W_in[12][9] = 21'b000000000000100101101;
    W_in[12][10] = 21'b000000000000010001011;
    W_in[12][11] = 21'b000000000000110111100;
    W_in[12][12] = 21'b111111111111110001000;
    W_in[12][13] = 21'b000000000000011100110;
    W_in[12][14] = 21'b000000000000011100100;
    W_in[12][15] = 21'b000000000000001100001;
    W_in[12][16] = 21'b111111111111110101101;
    W_in[12][17] = 21'b000000000000101011101;
    W_in[12][18] = 21'b000000000000111111110;
    W_in[12][19] = 21'b000000000000100011100;
    W_in[12][20] = 21'b111111111111111001101;
    W_in[12][21] = 21'b000000000000001011110;
    W_in[12][22] = 21'b000000000000101100011;
    W_in[12][23] = 21'b000000000000001010000;
    W_in[12][24] = 21'b000000000000000011111;
    W_in[12][25] = 21'b111111111111110101001;
    W_in[12][26] = 21'b111111111111000100110;
    W_in[12][27] = 21'b000000000000001101100;
    W_in[12][28] = 21'b000000000000011111010;
    W_in[12][29] = 21'b000000000000000010110;
    W_in[12][30] = 21'b000000000000100111101;
    W_in[12][31] = 21'b000000000000100001111;
    W_in[12][32] = 21'b111111111111110110110;
    W_in[12][33] = 21'b111111111111011011111;
    W_in[12][34] = 21'b111111111111001110000;
    W_in[12][35] = 21'b111111111111100111011;
    W_in[12][36] = 21'b111111111111100100010;
    W_in[12][37] = 21'b111111111110101101001;
    W_in[12][38] = 21'b000000000000001110010;
    W_in[12][39] = 21'b111111111111111011100;
    W_in[12][40] = 21'b111111111111110100110;
    W_in[12][41] = 21'b000000000000110110110;
    W_in[12][42] = 21'b111111111111010101110;
    W_in[12][43] = 21'b000000000000100010110;
    W_in[12][44] = 21'b000000000000000000011;
    W_in[12][45] = 21'b111111111111100000100;
    W_in[12][46] = 21'b111111111111011010101;
    W_in[12][47] = 21'b000000000000101010111;
    W_in[12][48] = 21'b000000000000010001101;
    W_in[12][49] = 21'b000000000001001011101;
    W_in[12][50] = 21'b111111111111111111110;
    W_in[12][51] = 21'b000000000000001111011;
    W_in[12][52] = 21'b111111111111101101010;
    W_in[12][53] = 21'b111111111111010001111;
    W_in[12][54] = 21'b111111111111001011001;
    W_in[12][55] = 21'b111111111111100101110;
    W_in[12][56] = 21'b000000000000111011000;
    W_in[12][57] = 21'b111111111111101101010;
    W_in[12][58] = 21'b000000000000111100111;
    W_in[12][59] = 21'b111111111111110010001;
    W_in[12][60] = 21'b111111111110111010001;
    W_in[12][61] = 21'b111111111110010010000;
    W_in[12][62] = 21'b111111111110000000111;
    W_in[12][63] = 21'b000000000000011011111;
    W_in[13][0] = 21'b000000000000110010110;
    W_in[13][1] = 21'b000000000000010001101;
    W_in[13][2] = 21'b000000000000001011011;
    W_in[13][3] = 21'b000000000000000000110;
    W_in[13][4] = 21'b000000000000000111110;
    W_in[13][5] = 21'b000000000000100110100;
    W_in[13][6] = 21'b111111111111001101001;
    W_in[13][7] = 21'b111111111111010110100;
    W_in[13][8] = 21'b000000000000000001010;
    W_in[13][9] = 21'b000000000001000000100;
    W_in[13][10] = 21'b000000000000100001010;
    W_in[13][11] = 21'b111111111110111100101;
    W_in[13][12] = 21'b111111111111010111000;
    W_in[13][13] = 21'b000000000000101011100;
    W_in[13][14] = 21'b111111111111110010110;
    W_in[13][15] = 21'b000000000000110011010;
    W_in[13][16] = 21'b111111111111000011100;
    W_in[13][17] = 21'b000000000000011101101;
    W_in[13][18] = 21'b000000000001001000100;
    W_in[13][19] = 21'b111111111111010100010;
    W_in[13][20] = 21'b111111111111011001101;
    W_in[13][21] = 21'b111111111111000100001;
    W_in[13][22] = 21'b000000000000100011011;
    W_in[13][23] = 21'b000000000001010011111;
    W_in[13][24] = 21'b000000000000011111000;
    W_in[13][25] = 21'b111111111111100001011;
    W_in[13][26] = 21'b111111111111100110000;
    W_in[13][27] = 21'b111111111111011110110;
    W_in[13][28] = 21'b111111111111101010100;
    W_in[13][29] = 21'b111111111111001101100;
    W_in[13][30] = 21'b111111111111110001111;
    W_in[13][31] = 21'b111111111111001100111;
    W_in[13][32] = 21'b000000000000100111010;
    W_in[13][33] = 21'b111111111111101111101;
    W_in[13][34] = 21'b111111111111011111100;
    W_in[13][35] = 21'b000000000000101001011;
    W_in[13][36] = 21'b111111111110110110111;
    W_in[13][37] = 21'b000000000000001010100;
    W_in[13][38] = 21'b111111111111111110010;
    W_in[13][39] = 21'b111111111111011111100;
    W_in[13][40] = 21'b000000000000101101101;
    W_in[13][41] = 21'b000000000000010111000;
    W_in[13][42] = 21'b000000000000111011111;
    W_in[13][43] = 21'b000000000000110011011;
    W_in[13][44] = 21'b000000000000000011001;
    W_in[13][45] = 21'b000000000000111010101;
    W_in[13][46] = 21'b000000000000010000011;
    W_in[13][47] = 21'b111111111111110010011;
    W_in[13][48] = 21'b111111111111010001010;
    W_in[13][49] = 21'b111111111111110110110;
    W_in[13][50] = 21'b111111111111100101001;
    W_in[13][51] = 21'b000000000000011101001;
    W_in[13][52] = 21'b000000000000101011100;
    W_in[13][53] = 21'b000000000000011000100;
    W_in[13][54] = 21'b111111111111000011000;
    W_in[13][55] = 21'b000000000001001100110;
    W_in[13][56] = 21'b000000000000100110100;
    W_in[13][57] = 21'b111111111111110000101;
    W_in[13][58] = 21'b111111111111111011100;
    W_in[13][59] = 21'b000000000000110111110;
    W_in[13][60] = 21'b111111111110111011100;
    W_in[13][61] = 21'b111111111111111100110;
    W_in[13][62] = 21'b111111111111100100100;
    W_in[13][63] = 21'b111111111111101000000;
    W_in[14][0] = 21'b000000000000010110111;
    W_in[14][1] = 21'b000000000000011111101;
    W_in[14][2] = 21'b111111111111110100001;
    W_in[14][3] = 21'b000000000000001100011;
    W_in[14][4] = 21'b000000000000110011010;
    W_in[14][5] = 21'b000000000000010110010;
    W_in[14][6] = 21'b111111111110110110100;
    W_in[14][7] = 21'b000000000000010111001;
    W_in[14][8] = 21'b111111111110100000110;
    W_in[14][9] = 21'b111111111111110011010;
    W_in[14][10] = 21'b111111111111111110111;
    W_in[14][11] = 21'b111111111111100011111;
    W_in[14][12] = 21'b111111111111001000100;
    W_in[14][13] = 21'b000000000000011001010;
    W_in[14][14] = 21'b111111111111111100100;
    W_in[14][15] = 21'b111111111110101001101;
    W_in[14][16] = 21'b000000000000100001001;
    W_in[14][17] = 21'b000000000000100101001;
    W_in[14][18] = 21'b111111111110100001000;
    W_in[14][19] = 21'b111111111110111100111;
    W_in[14][20] = 21'b000000000000110100111;
    W_in[14][21] = 21'b111111111111001101111;
    W_in[14][22] = 21'b000000000000010101101;
    W_in[14][23] = 21'b111111111111010000011;
    W_in[14][24] = 21'b000000000000011001011;
    W_in[14][25] = 21'b111111111111010100111;
    W_in[14][26] = 21'b000000000001001010111;
    W_in[14][27] = 21'b111111111111110011111;
    W_in[14][28] = 21'b000000000000101101000;
    W_in[14][29] = 21'b000000000001000110111;
    W_in[14][30] = 21'b111111111111110110001;
    W_in[14][31] = 21'b000000000000000000010;
    W_in[14][32] = 21'b000000000001010111000;
    W_in[14][33] = 21'b111111111110111110100;
    W_in[14][34] = 21'b111111111111000010111;
    W_in[14][35] = 21'b111111111111100010110;
    W_in[14][36] = 21'b000000000001010000110;
    W_in[14][37] = 21'b000000000001000010111;
    W_in[14][38] = 21'b111111111111010110100;
    W_in[14][39] = 21'b111111111110101011101;
    W_in[14][40] = 21'b000000000000100011100;
    W_in[14][41] = 21'b111111111111111011010;
    W_in[14][42] = 21'b111111111111000011101;
    W_in[14][43] = 21'b000000000000001011001;
    W_in[14][44] = 21'b111111111111101011011;
    W_in[14][45] = 21'b000000000000100110100;
    W_in[14][46] = 21'b111111111111110001110;
    W_in[14][47] = 21'b111111111111110001100;
    W_in[14][48] = 21'b111111111111100111111;
    W_in[14][49] = 21'b111111111111111111001;
    W_in[14][50] = 21'b111111111111000011100;
    W_in[14][51] = 21'b111111111111100110101;
    W_in[14][52] = 21'b111111111110111111000;
    W_in[14][53] = 21'b000000000000110110101;
    W_in[14][54] = 21'b111111111111111000000;
    W_in[14][55] = 21'b111111111111100011100;
    W_in[14][56] = 21'b111111111111100100101;
    W_in[14][57] = 21'b000000000000111001101;
    W_in[14][58] = 21'b000000000000111101110;
    W_in[14][59] = 21'b000000000001001101101;
    W_in[14][60] = 21'b000000000001111001011;
    W_in[14][61] = 21'b000000000001010001011;
    W_in[14][62] = 21'b000000000010001011110;
    W_in[14][63] = 21'b000000000001100111101;
    W_in[15][0] = 21'b111111111110100110010;
    W_in[15][1] = 21'b000000000001000001011;
    W_in[15][2] = 21'b000000000000000100111;
    W_in[15][3] = 21'b000000000001000111000;
    W_in[15][4] = 21'b111111111110101110010;
    W_in[15][5] = 21'b000000000000010001101;
    W_in[15][6] = 21'b111111111110111000010;
    W_in[15][7] = 21'b000000000000100111101;
    W_in[15][8] = 21'b111111111110010001110;
    W_in[15][9] = 21'b111111111110100110000;
    W_in[15][10] = 21'b000000000001001010001;
    W_in[15][11] = 21'b111111111110100110001;
    W_in[15][12] = 21'b111111111110101000111;
    W_in[15][13] = 21'b000000000000100101001;
    W_in[15][14] = 21'b000000000000011111101;
    W_in[15][15] = 21'b000000000000011111110;
    W_in[15][16] = 21'b000000000001010101001;
    W_in[15][17] = 21'b111111111111101110010;
    W_in[15][18] = 21'b111111111111111111101;
    W_in[15][19] = 21'b000000000001100101100;
    W_in[15][20] = 21'b111111111111110000100;
    W_in[15][21] = 21'b111111111111000011100;
    W_in[15][22] = 21'b111111111111101001011;
    W_in[15][23] = 21'b111111111111100010111;
    W_in[15][24] = 21'b111111111110110000110;
    W_in[15][25] = 21'b111111111111110001011;
    W_in[15][26] = 21'b111111111110111111011;
    W_in[15][27] = 21'b111111111110101111111;
    W_in[15][28] = 21'b000000000001101001110;
    W_in[15][29] = 21'b000000000000100011011;
    W_in[15][30] = 21'b000000000000000110011;
    W_in[15][31] = 21'b000000000000111010101;
    W_in[15][32] = 21'b000000000000100010100;
    W_in[15][33] = 21'b111111111111110000001;
    W_in[15][34] = 21'b000000000000111001010;
    W_in[15][35] = 21'b000000000000011100110;
    W_in[15][36] = 21'b111111111110111011110;
    W_in[15][37] = 21'b111111111110101101110;
    W_in[15][38] = 21'b000000000000100010011;
    W_in[15][39] = 21'b111111111111111101010;
    W_in[15][40] = 21'b111111111110100000101;
    W_in[15][41] = 21'b111111111110101100110;
    W_in[15][42] = 21'b000000000001000001011;
    W_in[15][43] = 21'b000000000000000101111;
    W_in[15][44] = 21'b000000000000010110001;
    W_in[15][45] = 21'b000000000001100011100;
    W_in[15][46] = 21'b111111111111110111000;
    W_in[15][47] = 21'b000000000001010000001;
    W_in[15][48] = 21'b000000000000001001100;
    W_in[15][49] = 21'b111111111111110110110;
    W_in[15][50] = 21'b111111111111010100111;
    W_in[15][51] = 21'b000000000000101100110;
    W_in[15][52] = 21'b111111111111101100001;
    W_in[15][53] = 21'b111111111110101111001;
    W_in[15][54] = 21'b000000000001100010010;
    W_in[15][55] = 21'b000000000000001111001;
    W_in[15][56] = 21'b111111111111010001101;
    W_in[15][57] = 21'b000000000000101101100;
    W_in[15][58] = 21'b111111111111011001111;
    W_in[15][59] = 21'b000000000001011000101;
    W_in[15][60] = 21'b000000000001010111010;
    W_in[15][61] = 21'b000000000000010100110;
    W_in[15][62] = 21'b000000000000000111001;
    W_in[15][63] = 21'b000000000001001011111;

    // Initialize W_hr weights
    W_hr[0][0] = 21'b000000000000000011100;
    W_hr[0][1] = 21'b000000000000001001101;
    W_hr[0][2] = 21'b000000000000001111101;
    W_hr[0][3] = 21'b111111111111010111001;
    W_hr[0][4] = 21'b000000000001000110001;
    W_hr[0][5] = 21'b000000000001001011011;
    W_hr[0][6] = 21'b000000000001001010110;
    W_hr[0][7] = 21'b111111111110110110001;
    W_hr[0][8] = 21'b000000000000111111100;
    W_hr[0][9] = 21'b000000000001000111111;
    W_hr[0][10] = 21'b111111111111011111011;
    W_hr[0][11] = 21'b111111111111011000111;
    W_hr[0][12] = 21'b000000000000011111010;
    W_hr[0][13] = 21'b000000000000101000000;
    W_hr[0][14] = 21'b000000000001011010000;
    W_hr[0][15] = 21'b111111111111000011010;
    W_hr[1][0] = 21'b000000000000110111000;
    W_hr[1][1] = 21'b000000000000011100101;
    W_hr[1][2] = 21'b111111111111101011000;
    W_hr[1][3] = 21'b000000000000100000101;
    W_hr[1][4] = 21'b000000000001101000010;
    W_hr[1][5] = 21'b111111111110011110010;
    W_hr[1][6] = 21'b000000000000000001101;
    W_hr[1][7] = 21'b000000000001000111110;
    W_hr[1][8] = 21'b000000000000110110011;
    W_hr[1][9] = 21'b000000000000000001011;
    W_hr[1][10] = 21'b111111111110000010100;
    W_hr[1][11] = 21'b000000000001110001111;
    W_hr[1][12] = 21'b000000000001011111110;
    W_hr[1][13] = 21'b000000000000100010111;
    W_hr[1][14] = 21'b111111111110110100110;
    W_hr[1][15] = 21'b000000000010100101111;
    W_hr[2][0] = 21'b111111111111110101110;
    W_hr[2][1] = 21'b111111111111101100110;
    W_hr[2][2] = 21'b000000000000100100011;
    W_hr[2][3] = 21'b111111111111001100011;
    W_hr[2][4] = 21'b111111111111010010111;
    W_hr[2][5] = 21'b111111111111111001111;
    W_hr[2][6] = 21'b000000000010111011100;
    W_hr[2][7] = 21'b111111111110100010001;
    W_hr[2][8] = 21'b111111111111110101110;
    W_hr[2][9] = 21'b000000000001101100111;
    W_hr[2][10] = 21'b000000000010011111001;
    W_hr[2][11] = 21'b111111111110010000010;
    W_hr[2][12] = 21'b111111111111010110011;
    W_hr[2][13] = 21'b111111111110110011001;
    W_hr[2][14] = 21'b111111111111001011100;
    W_hr[2][15] = 21'b000000000001001110101;
    W_hr[3][0] = 21'b000000000000000011100;
    W_hr[3][1] = 21'b000000000000001001101;
    W_hr[3][2] = 21'b000000000000001111101;
    W_hr[3][3] = 21'b111111111111010111001;
    W_hr[3][4] = 21'b000000000001000110001;
    W_hr[3][5] = 21'b000000000001001011011;
    W_hr[3][6] = 21'b000000000001001010110;
    W_hr[3][7] = 21'b111111111110110110001;
    W_hr[3][8] = 21'b000000000000111111100;
    W_hr[3][9] = 21'b000000000001000111111;
    W_hr[3][10] = 21'b111111111111011111011;
    W_hr[3][11] = 21'b111111111111011000111;
    W_hr[3][12] = 21'b000000000000011111010;
    W_hr[3][13] = 21'b000000000000101000000;
    W_hr[3][14] = 21'b000000000001011010000;
    W_hr[3][15] = 21'b111111111111000011010;
    W_hr[4][0] = 21'b000000000000110111000;
    W_hr[4][1] = 21'b000000000000011100101;
    W_hr[4][2] = 21'b111111111111101011000;
    W_hr[4][3] = 21'b000000000000100000101;
    W_hr[4][4] = 21'b000000000001101000010;
    W_hr[4][5] = 21'b111111111110011110010;
    W_hr[4][6] = 21'b000000000000000001101;
    W_hr[4][7] = 21'b000000000001000111110;
    W_hr[4][8] = 21'b000000000000110110011;
    W_hr[4][9] = 21'b000000000000000001011;
    W_hr[4][10] = 21'b111111111110000010100;
    W_hr[4][11] = 21'b000000000001110001111;
    W_hr[4][12] = 21'b000000000001011111110;
    W_hr[4][13] = 21'b000000000000100010111;
    W_hr[4][14] = 21'b111111111110110100110;
    W_hr[4][15] = 21'b000000000010100101111;
    W_hr[5][0] = 21'b111111111111110101110;
    W_hr[5][1] = 21'b111111111111101100110;
    W_hr[5][2] = 21'b000000000000100100011;
    W_hr[5][3] = 21'b111111111111001100011;
    W_hr[5][4] = 21'b111111111111010010111;
    W_hr[5][5] = 21'b111111111111111001111;
    W_hr[5][6] = 21'b000000000010111011100;
    W_hr[5][7] = 21'b111111111110100010001;
    W_hr[5][8] = 21'b111111111111110101110;
    W_hr[5][9] = 21'b000000000001101100111;
    W_hr[5][10] = 21'b000000000010011111001;
    W_hr[5][11] = 21'b111111111110010000010;
    W_hr[5][12] = 21'b111111111111010110011;
    W_hr[5][13] = 21'b111111111110110011001;
    W_hr[5][14] = 21'b111111111111001011100;
    W_hr[5][15] = 21'b000000000001001110101;
    W_hr[6][0] = 21'b000000000000000011100;
    W_hr[6][1] = 21'b000000000000001001101;
    W_hr[6][2] = 21'b000000000000001111101;
    W_hr[6][3] = 21'b111111111111010111001;
    W_hr[6][4] = 21'b000000000001000110001;
    W_hr[6][5] = 21'b000000000001001011011;
    W_hr[6][6] = 21'b000000000001001010110;
    W_hr[6][7] = 21'b111111111110110110001;
    W_hr[6][8] = 21'b000000000000111111100;
    W_hr[6][9] = 21'b000000000001000111111;
    W_hr[6][10] = 21'b111111111111011111011;
    W_hr[6][11] = 21'b111111111111011000111;
    W_hr[6][12] = 21'b000000000000011111010;
    W_hr[6][13] = 21'b000000000000101000000;
    W_hr[6][14] = 21'b000000000001011010000;
    W_hr[6][15] = 21'b111111111111000011010;
    W_hr[7][0] = 21'b000000000000110111000;
    W_hr[7][1] = 21'b000000000000011100101;
    W_hr[7][2] = 21'b111111111111101011000;
    W_hr[7][3] = 21'b000000000000100000101;
    W_hr[7][4] = 21'b000000000001101000010;
    W_hr[7][5] = 21'b111111111110011110010;
    W_hr[7][6] = 21'b000000000000000001101;
    W_hr[7][7] = 21'b000000000001000111110;
    W_hr[7][8] = 21'b000000000000110110011;
    W_hr[7][9] = 21'b000000000000000001011;
    W_hr[7][10] = 21'b111111111110000010100;
    W_hr[7][11] = 21'b000000000001110001111;
    W_hr[7][12] = 21'b000000000001011111110;
    W_hr[7][13] = 21'b000000000000100010111;
    W_hr[7][14] = 21'b111111111110110100110;
    W_hr[7][15] = 21'b000000000010100101111;
    W_hr[8][0] = 21'b111111111111110101110;
    W_hr[8][1] = 21'b111111111111101100110;
    W_hr[8][2] = 21'b000000000000100100011;
    W_hr[8][3] = 21'b111111111111001100011;
    W_hr[8][4] = 21'b111111111111010010111;
    W_hr[8][5] = 21'b111111111111111001111;
    W_hr[8][6] = 21'b000000000010111011100;
    W_hr[8][7] = 21'b111111111110100010001;
    W_hr[8][8] = 21'b111111111111110101110;
    W_hr[8][9] = 21'b000000000001101100111;
    W_hr[8][10] = 21'b000000000010011111001;
    W_hr[8][11] = 21'b111111111110010000010;
    W_hr[8][12] = 21'b111111111111010110011;
    W_hr[8][13] = 21'b111111111110110011001;
    W_hr[8][14] = 21'b111111111111001011100;
    W_hr[8][15] = 21'b000000000001001110101;
    W_hr[9][0] = 21'b000000000000000011100;
    W_hr[9][1] = 21'b000000000000001001101;
    W_hr[9][2] = 21'b000000000000001111101;
    W_hr[9][3] = 21'b111111111111010111001;
    W_hr[9][4] = 21'b000000000001000110001;
    W_hr[9][5] = 21'b000000000001001011011;
    W_hr[9][6] = 21'b000000000001001010110;
    W_hr[9][7] = 21'b111111111110110110001;
    W_hr[9][8] = 21'b000000000000111111100;
    W_hr[9][9] = 21'b000000000001000111111;
    W_hr[9][10] = 21'b111111111111011111011;
    W_hr[9][11] = 21'b111111111111011000111;
    W_hr[9][12] = 21'b000000000000011111010;
    W_hr[9][13] = 21'b000000000000101000000;
    W_hr[9][14] = 21'b000000000001011010000;
    W_hr[9][15] = 21'b111111111111000011010;
    W_hr[10][0] = 21'b000000000000110111000;
    W_hr[10][1] = 21'b000000000000011100101;
    W_hr[10][2] = 21'b111111111111101011000;
    W_hr[10][3] = 21'b000000000000100000101;
    W_hr[10][4] = 21'b000000000001101000010;
    W_hr[10][5] = 21'b111111111110011110010;
    W_hr[10][6] = 21'b000000000000000001101;
    W_hr[10][7] = 21'b000000000001000111110;
    W_hr[10][8] = 21'b000000000000110110011;
    W_hr[10][9] = 21'b000000000000000001011;
    W_hr[10][10] = 21'b111111111110000010100;
    W_hr[10][11] = 21'b000000000001110001111;
    W_hr[10][12] = 21'b000000000001011111110;
    W_hr[10][13] = 21'b000000000000100010111;
    W_hr[10][14] = 21'b111111111110110100110;
    W_hr[10][15] = 21'b000000000010100101111;
    W_hr[11][0] = 21'b111111111111110101110;
    W_hr[11][1] = 21'b111111111111101100110;
    W_hr[11][2] = 21'b000000000000100100011;
    W_hr[11][3] = 21'b111111111111001100011;
    W_hr[11][4] = 21'b111111111111010010111;
    W_hr[11][5] = 21'b111111111111111001111;
    W_hr[11][6] = 21'b000000000010111011100;
    W_hr[11][7] = 21'b111111111110100010001;
    W_hr[11][8] = 21'b111111111111110101110;
    W_hr[11][9] = 21'b000000000001101100111;
    W_hr[11][10] = 21'b000000000010011111001;
    W_hr[11][11] = 21'b111111111110010000010;
    W_hr[11][12] = 21'b111111111111010110011;
    W_hr[11][13] = 21'b111111111110110011001;
    W_hr[11][14] = 21'b111111111111001011100;
    W_hr[11][15] = 21'b000000000001001110101;
    W_hr[12][0] = 21'b000000000000000011100;
    W_hr[12][1] = 21'b000000000000001001101;
    W_hr[12][2] = 21'b000000000000001111101;
    W_hr[12][3] = 21'b111111111111010111001;
    W_hr[12][4] = 21'b000000000001000110001;
    W_hr[12][5] = 21'b000000000001001011011;
    W_hr[12][6] = 21'b000000000001001010110;
    W_hr[12][7] = 21'b111111111110110110001;
    W_hr[12][8] = 21'b000000000000111111100;
    W_hr[12][9] = 21'b000000000001000111111;
    W_hr[12][10] = 21'b111111111111011111011;
    W_hr[12][11] = 21'b111111111111011000111;
    W_hr[12][12] = 21'b000000000000011111010;
    W_hr[12][13] = 21'b000000000000101000000;
    W_hr[12][14] = 21'b000000000001011010000;
    W_hr[12][15] = 21'b111111111111000011010;
    W_hr[13][0] = 21'b000000000000110111000;
    W_hr[13][1] = 21'b000000000000011100101;
    W_hr[13][2] = 21'b111111111111101011000;
    W_hr[13][3] = 21'b000000000000100000101;
    W_hr[13][4] = 21'b000000000001101000010;
    W_hr[13][5] = 21'b111111111110011110010;
    W_hr[13][6] = 21'b000000000000000001101;
    W_hr[13][7] = 21'b000000000001000111110;
    W_hr[13][8] = 21'b000000000000110110011;
    W_hr[13][9] = 21'b000000000000000001011;
    W_hr[13][10] = 21'b111111111110000010100;
    W_hr[13][11] = 21'b000000000001110001111;
    W_hr[13][12] = 21'b000000000001011111110;
    W_hr[13][13] = 21'b000000000000100010111;
    W_hr[13][14] = 21'b111111111110110100110;
    W_hr[13][15] = 21'b000000000010100101111;
    W_hr[14][0] = 21'b111111111111110101110;
    W_hr[14][1] = 21'b111111111111101100110;
    W_hr[14][2] = 21'b000000000000100100011;
    W_hr[14][3] = 21'b111111111111001100011;
    W_hr[14][4] = 21'b111111111111010010111;
    W_hr[14][5] = 21'b111111111111111001111;
    W_hr[14][6] = 21'b000000000010111011100;
    W_hr[14][7] = 21'b111111111110100010001;
    W_hr[14][8] = 21'b111111111111110101110;
    W_hr[14][9] = 21'b000000000001101100111;
    W_hr[14][10] = 21'b000000000010011111001;
    W_hr[14][11] = 21'b111111111110010000010;
    W_hr[14][12] = 21'b111111111111010110011;
    W_hr[14][13] = 21'b111111111110110011001;
    W_hr[14][14] = 21'b111111111111001011100;
    W_hr[14][15] = 21'b000000000001001110101;
    W_hr[15][0] = 21'b000000000000000011100;
    W_hr[15][1] = 21'b000000000000001001101;
    W_hr[15][2] = 21'b000000000000001111101;
    W_hr[15][3] = 21'b111111111111010111001;
    W_hr[15][4] = 21'b000000000001000110001;
    W_hr[15][5] = 21'b000000000001001011011;
    W_hr[15][6] = 21'b000000000001001010110;
    W_hr[15][7] = 21'b111111111110110110001;
    W_hr[15][8] = 21'b000000000000111111100;
    W_hr[15][9] = 21'b000000000001000111111;
    W_hr[15][10] = 21'b111111111111011111011;
    W_hr[15][11] = 21'b111111111111011000111;
    W_hr[15][12] = 21'b000000000000011111010;
    W_hr[15][13] = 21'b000000000000101000000;
    W_hr[15][14] = 21'b000000000001011010000;
    W_hr[15][15] = 21'b111111111111000011010;

    // Initialize W_hz weights
    W_hz[0][0] = 21'b000000000000110111000;
    W_hz[0][1] = 21'b000000000000011100101;
    W_hz[0][2] = 21'b111111111111101011000;
    W_hz[0][3] = 21'b000000000000100000101;
    W_hz[0][4] = 21'b000000000001101000010;
    W_hz[0][5] = 21'b111111111110011110010;
    W_hz[0][6] = 21'b000000000000000001101;
    W_hz[0][7] = 21'b000000000001000111110;
    W_hz[0][8] = 21'b000000000000110110011;
    W_hz[0][9] = 21'b000000000000000001011;
    W_hz[0][10] = 21'b111111111110000010100;
    W_hz[0][11] = 21'b000000000001110001111;
    W_hz[0][12] = 21'b000000000001011111110;
    W_hz[0][13] = 21'b000000000000100010111;
    W_hz[0][14] = 21'b111111111110110100110;
    W_hz[0][15] = 21'b000000000010100101111;
    W_hz[1][0] = 21'b111111111111110101110;
    W_hz[1][1] = 21'b111111111111101100110;
    W_hz[1][2] = 21'b000000000000100100011;
    W_hz[1][3] = 21'b111111111111001100011;
    W_hz[1][4] = 21'b111111111111010010111;
    W_hz[1][5] = 21'b111111111111111001111;
    W_hz[1][6] = 21'b000000000010111011100;
    W_hz[1][7] = 21'b111111111110100010001;
    W_hz[1][8] = 21'b111111111111110101110;
    W_hz[1][9] = 21'b000000000001101100111;
    W_hz[1][10] = 21'b000000000010011111001;
    W_hz[1][11] = 21'b111111111110010000010;
    W_hz[1][12] = 21'b111111111111010110011;
    W_hz[1][13] = 21'b111111111110110011001;
    W_hz[1][14] = 21'b111111111111001011100;
    W_hz[1][15] = 21'b000000000001001110101;
    W_hz[2][0] = 21'b000000000000000011100;
    W_hz[2][1] = 21'b000000000000001001101;
    W_hz[2][2] = 21'b000000000000001111101;
    W_hz[2][3] = 21'b111111111111010111001;
    W_hz[2][4] = 21'b000000000001000110001;
    W_hz[2][5] = 21'b000000000001001011011;
    W_hz[2][6] = 21'b000000000001001010110;
    W_hz[2][7] = 21'b111111111110110110001;
    W_hz[2][8] = 21'b000000000000111111100;
    W_hz[2][9] = 21'b000000000001000111111;
    W_hz[2][10] = 21'b111111111111011111011;
    W_hz[2][11] = 21'b111111111111011000111;
    W_hz[2][12] = 21'b000000000000011111010;
    W_hz[2][13] = 21'b000000000000101000000;
    W_hz[2][14] = 21'b000000000001011010000;
    W_hz[2][15] = 21'b111111111111000011010;
    W_hz[3][0] = 21'b000000000000110111000;
    W_hz[3][1] = 21'b000000000000011100101;
    W_hz[3][2] = 21'b111111111111101011000;
    W_hz[3][3] = 21'b000000000000100000101;
    W_hz[3][4] = 21'b000000000001101000010;
    W_hz[3][5] = 21'b111111111110011110010;
    W_hz[3][6] = 21'b000000000000000001101;
    W_hz[3][7] = 21'b000000000001000111110;
    W_hz[3][8] = 21'b000000000000110110011;
    W_hz[3][9] = 21'b000000000000000001011;
    W_hz[3][10] = 21'b111111111110000010100;
    W_hz[3][11] = 21'b000000000001110001111;
    W_hz[3][12] = 21'b000000000001011111110;
    W_hz[3][13] = 21'b000000000000100010111;
    W_hz[3][14] = 21'b111111111110110100110;
    W_hz[3][15] = 21'b000000000010100101111;
    W_hz[4][0] = 21'b111111111111110101110;
    W_hz[4][1] = 21'b111111111111101100110;
    W_hz[4][2] = 21'b000000000000100100011;
    W_hz[4][3] = 21'b111111111111001100011;
    W_hz[4][4] = 21'b111111111111010010111;
    W_hz[4][5] = 21'b111111111111111001111;
    W_hz[4][6] = 21'b000000000010111011100;
    W_hz[4][7] = 21'b111111111110100010001;
    W_hz[4][8] = 21'b111111111111110101110;
    W_hz[4][9] = 21'b000000000001101100111;
    W_hz[4][10] = 21'b000000000010011111001;
    W_hz[4][11] = 21'b111111111110010000010;
    W_hz[4][12] = 21'b111111111111010110011;
    W_hz[4][13] = 21'b111111111110110011001;
    W_hz[4][14] = 21'b111111111111001011100;
    W_hz[4][15] = 21'b000000000001001110101;
    W_hz[5][0] = 21'b000000000000000011100;
    W_hz[5][1] = 21'b000000000000001001101;
    W_hz[5][2] = 21'b000000000000001111101;
    W_hz[5][3] = 21'b111111111111010111001;
    W_hz[5][4] = 21'b000000000001000110001;
    W_hz[5][5] = 21'b000000000001001011011;
    W_hz[5][6] = 21'b000000000001001010110;
    W_hz[5][7] = 21'b111111111110110110001;
    W_hz[5][8] = 21'b000000000000111111100;
    W_hz[5][9] = 21'b000000000001000111111;
    W_hz[5][10] = 21'b111111111111011111011;
    W_hz[5][11] = 21'b111111111111011000111;
    W_hz[5][12] = 21'b000000000000011111010;
    W_hz[5][13] = 21'b000000000000101000000;
    W_hz[5][14] = 21'b000000000001011010000;
    W_hz[5][15] = 21'b111111111111000011010;
    W_hz[6][0] = 21'b000000000000110111000;
    W_hz[6][1] = 21'b000000000000011100101;
    W_hz[6][2] = 21'b111111111111101011000;
    W_hz[6][3] = 21'b000000000000100000101;
    W_hz[6][4] = 21'b000000000001101000010;
    W_hz[6][5] = 21'b111111111110011110010;
    W_hz[6][6] = 21'b000000000000000001101;
    W_hz[6][7] = 21'b000000000001000111110;
    W_hz[6][8] = 21'b000000000000110110011;
    W_hz[6][9] = 21'b000000000000000001011;
    W_hz[6][10] = 21'b111111111110000010100;
    W_hz[6][11] = 21'b000000000001110001111;
    W_hz[6][12] = 21'b000000000001011111110;
    W_hz[6][13] = 21'b000000000000100010111;
    W_hz[6][14] = 21'b111111111110110100110;
    W_hz[6][15] = 21'b000000000010100101111;
    W_hz[7][0] = 21'b111111111111110101110;
    W_hz[7][1] = 21'b111111111111101100110;
    W_hz[7][2] = 21'b000000000000100100011;
    W_hz[7][3] = 21'b111111111111001100011;
    W_hz[7][4] = 21'b111111111111010010111;
    W_hz[7][5] = 21'b111111111111111001111;
    W_hz[7][6] = 21'b000000000010111011100;
    W_hz[7][7] = 21'b111111111110100010001;
    W_hz[7][8] = 21'b111111111111110101110;
    W_hz[7][9] = 21'b000000000001101100111;
    W_hz[7][10] = 21'b000000000010011111001;
    W_hz[7][11] = 21'b111111111110010000010;
    W_hz[7][12] = 21'b111111111111010110011;
    W_hz[7][13] = 21'b111111111110110011001;
    W_hz[7][14] = 21'b111111111111001011100;
    W_hz[7][15] = 21'b000000000001001110101;
    W_hz[8][0] = 21'b000000000000000011100;
    W_hz[8][1] = 21'b000000000000001001101;
    W_hz[8][2] = 21'b000000000000001111101;
    W_hz[8][3] = 21'b111111111111010111001;
    W_hz[8][4] = 21'b000000000001000110001;
    W_hz[8][5] = 21'b000000000001001011011;
    W_hz[8][6] = 21'b000000000001001010110;
    W_hz[8][7] = 21'b111111111110110110001;
    W_hz[8][8] = 21'b000000000000111111100;
    W_hz[8][9] = 21'b000000000001000111111;
    W_hz[8][10] = 21'b111111111111011111011;
    W_hz[8][11] = 21'b111111111111011000111;
    W_hz[8][12] = 21'b000000000000011111010;
    W_hz[8][13] = 21'b000000000000101000000;
    W_hz[8][14] = 21'b000000000001011010000;
    W_hz[8][15] = 21'b111111111111000011010;
    W_hz[9][0] = 21'b000000000000110111000;
    W_hz[9][1] = 21'b000000000000011100101;
    W_hz[9][2] = 21'b111111111111101011000;
    W_hz[9][3] = 21'b000000000000100000101;
    W_hz[9][4] = 21'b000000000001101000010;
    W_hz[9][5] = 21'b111111111110011110010;
    W_hz[9][6] = 21'b000000000000000001101;
    W_hz[9][7] = 21'b000000000001000111110;
    W_hz[9][8] = 21'b000000000000110110011;
    W_hz[9][9] = 21'b000000000000000001011;
    W_hz[9][10] = 21'b111111111110000010100;
    W_hz[9][11] = 21'b000000000001110001111;
    W_hz[9][12] = 21'b000000000001011111110;
    W_hz[9][13] = 21'b000000000000100010111;
    W_hz[9][14] = 21'b111111111110110100110;
    W_hz[9][15] = 21'b000000000010100101111;
    W_hz[10][0] = 21'b111111111111110101110;
    W_hz[10][1] = 21'b111111111111101100110;
    W_hz[10][2] = 21'b000000000000100100011;
    W_hz[10][3] = 21'b111111111111001100011;
    W_hz[10][4] = 21'b111111111111010010111;
    W_hz[10][5] = 21'b111111111111111001111;
    W_hz[10][6] = 21'b000000000010111011100;
    W_hz[10][7] = 21'b111111111110100010001;
    W_hz[10][8] = 21'b111111111111110101110;
    W_hz[10][9] = 21'b000000000001101100111;
    W_hz[10][10] = 21'b000000000010011111001;
    W_hz[10][11] = 21'b111111111110010000010;
    W_hz[10][12] = 21'b111111111111010110011;
    W_hz[10][13] = 21'b111111111110110011001;
    W_hz[10][14] = 21'b111111111111001011100;
    W_hz[10][15] = 21'b000000000001001110101;
    W_hz[11][0] = 21'b000000000000000011100;
    W_hz[11][1] = 21'b000000000000001001101;
    W_hz[11][2] = 21'b000000000000001111101;
    W_hz[11][3] = 21'b111111111111010111001;
    W_hz[11][4] = 21'b000000000001000110001;
    W_hz[11][5] = 21'b000000000001001011011;
    W_hz[11][6] = 21'b000000000001001010110;
    W_hz[11][7] = 21'b111111111110110110001;
    W_hz[11][8] = 21'b000000000000111111100;
    W_hz[11][9] = 21'b000000000001000111111;
    W_hz[11][10] = 21'b111111111111011111011;
    W_hz[11][11] = 21'b111111111111011000111;
    W_hz[11][12] = 21'b000000000000011111010;
    W_hz[11][13] = 21'b000000000000101000000;
    W_hz[11][14] = 21'b000000000001011010000;
    W_hz[11][15] = 21'b111111111111000011010;
    W_hz[12][0] = 21'b000000000000110111000;
    W_hz[12][1] = 21'b000000000000011100101;
    W_hz[12][2] = 21'b111111111111101011000;
    W_hz[12][3] = 21'b000000000000100000101;
    W_hz[12][4] = 21'b000000000001101000010;
    W_hz[12][5] = 21'b111111111110011110010;
    W_hz[12][6] = 21'b000000000000000001101;
    W_hz[12][7] = 21'b000000000001000111110;
    W_hz[12][8] = 21'b000000000000110110011;
    W_hz[12][9] = 21'b000000000000000001011;
    W_hz[12][10] = 21'b111111111110000010100;
    W_hz[12][11] = 21'b000000000001110001111;
    W_hz[12][12] = 21'b000000000001011111110;
    W_hz[12][13] = 21'b000000000000100010111;
    W_hz[12][14] = 21'b111111111110110100110;
    W_hz[12][15] = 21'b000000000010100101111;
    W_hz[13][0] = 21'b111111111111110101110;
    W_hz[13][1] = 21'b111111111111101100110;
    W_hz[13][2] = 21'b000000000000100100011;
    W_hz[13][3] = 21'b111111111111001100011;
    W_hz[13][4] = 21'b111111111111010010111;
    W_hz[13][5] = 21'b111111111111111001111;
    W_hz[13][6] = 21'b000000000010111011100;
    W_hz[13][7] = 21'b111111111110100010001;
    W_hz[13][8] = 21'b111111111111110101110;
    W_hz[13][9] = 21'b000000000001101100111;
    W_hz[13][10] = 21'b000000000010011111001;
    W_hz[13][11] = 21'b111111111110010000010;
    W_hz[13][12] = 21'b111111111111010110011;
    W_hz[13][13] = 21'b111111111110110011001;
    W_hz[13][14] = 21'b111111111111001011100;
    W_hz[13][15] = 21'b000000000001001110101;
    W_hz[14][0] = 21'b000000000000000011100;
    W_hz[14][1] = 21'b000000000000001001101;
    W_hz[14][2] = 21'b000000000000001111101;
    W_hz[14][3] = 21'b111111111111010111001;
    W_hz[14][4] = 21'b000000000001000110001;
    W_hz[14][5] = 21'b000000000001001011011;
    W_hz[14][6] = 21'b000000000001001010110;
    W_hz[14][7] = 21'b111111111110110110001;
    W_hz[14][8] = 21'b000000000000111111100;
    W_hz[14][9] = 21'b000000000001000111111;
    W_hz[14][10] = 21'b111111111111011111011;
    W_hz[14][11] = 21'b111111111111011000111;
    W_hz[14][12] = 21'b000000000000011111010;
    W_hz[14][13] = 21'b000000000000101000000;
    W_hz[14][14] = 21'b000000000001011010000;
    W_hz[14][15] = 21'b111111111111000011010;
    W_hz[15][0] = 21'b000000000000110111000;
    W_hz[15][1] = 21'b000000000000011100101;
    W_hz[15][2] = 21'b111111111111101011000;
    W_hz[15][3] = 21'b000000000000100000101;
    W_hz[15][4] = 21'b000000000001101000010;
    W_hz[15][5] = 21'b111111111110011110010;
    W_hz[15][6] = 21'b000000000000000001101;
    W_hz[15][7] = 21'b000000000001000111110;
    W_hz[15][8] = 21'b000000000000110110011;
    W_hz[15][9] = 21'b000000000000000001011;
    W_hz[15][10] = 21'b111111111110000010100;
    W_hz[15][11] = 21'b000000000001110001111;
    W_hz[15][12] = 21'b000000000001011111110;
    W_hz[15][13] = 21'b000000000000100010111;
    W_hz[15][14] = 21'b111111111110110100110;
    W_hz[15][15] = 21'b000000000010100101111;

    // Initialize W_hn weights
    W_hn[0][0] = 21'b111111111111110101110;
    W_hn[0][1] = 21'b111111111111101100110;
    W_hn[0][2] = 21'b000000000000100100011;
    W_hn[0][3] = 21'b111111111111001100011;
    W_hn[0][4] = 21'b111111111111010010111;
    W_hn[0][5] = 21'b111111111111111001111;
    W_hn[0][6] = 21'b000000000010111011100;
    W_hn[0][7] = 21'b111111111110100010001;
    W_hn[0][8] = 21'b111111111111110101110;
    W_hn[0][9] = 21'b000000000001101100111;
    W_hn[0][10] = 21'b000000000010011111001;
    W_hn[0][11] = 21'b111111111110010000010;
    W_hn[0][12] = 21'b111111111111010110011;
    W_hn[0][13] = 21'b111111111110110011001;
    W_hn[0][14] = 21'b111111111111001011100;
    W_hn[0][15] = 21'b000000000001001110101;
    W_hn[1][0] = 21'b000000000000000011100;
    W_hn[1][1] = 21'b000000000000001001101;
    W_hn[1][2] = 21'b000000000000001111101;
    W_hn[1][3] = 21'b111111111111010111001;
    W_hn[1][4] = 21'b000000000001000110001;
    W_hn[1][5] = 21'b000000000001001011011;
    W_hn[1][6] = 21'b000000000001001010110;
    W_hn[1][7] = 21'b111111111110110110001;
    W_hn[1][8] = 21'b000000000000111111100;
    W_hn[1][9] = 21'b000000000001000111111;
    W_hn[1][10] = 21'b111111111111011111011;
    W_hn[1][11] = 21'b111111111111011000111;
    W_hn[1][12] = 21'b000000000000011111010;
    W_hn[1][13] = 21'b000000000000101000000;
    W_hn[1][14] = 21'b000000000001011010000;
    W_hn[1][15] = 21'b111111111111000011010;
    W_hn[2][0] = 21'b000000000000110111000;
    W_hn[2][1] = 21'b000000000000011100101;
    W_hn[2][2] = 21'b111111111111101011000;
    W_hn[2][3] = 21'b000000000000100000101;
    W_hn[2][4] = 21'b000000000001101000010;
    W_hn[2][5] = 21'b111111111110011110010;
    W_hn[2][6] = 21'b000000000000000001101;
    W_hn[2][7] = 21'b000000000001000111110;
    W_hn[2][8] = 21'b000000000000110110011;
    W_hn[2][9] = 21'b000000000000000001011;
    W_hn[2][10] = 21'b111111111110000010100;
    W_hn[2][11] = 21'b000000000001110001111;
    W_hn[2][12] = 21'b000000000001011111110;
    W_hn[2][13] = 21'b000000000000100010111;
    W_hn[2][14] = 21'b111111111110110100110;
    W_hn[2][15] = 21'b000000000010100101111;
    W_hn[3][0] = 21'b111111111111110101110;
    W_hn[3][1] = 21'b111111111111101100110;
    W_hn[3][2] = 21'b000000000000100100011;
    W_hn[3][3] = 21'b111111111111001100011;
    W_hn[3][4] = 21'b111111111111010010111;
    W_hn[3][5] = 21'b111111111111111001111;
    W_hn[3][6] = 21'b000000000010111011100;
    W_hn[3][7] = 21'b111111111110100010001;
    W_hn[3][8] = 21'b111111111111110101110;
    W_hn[3][9] = 21'b000000000001101100111;
    W_hn[3][10] = 21'b000000000010011111001;
    W_hn[3][11] = 21'b111111111110010000010;
    W_hn[3][12] = 21'b111111111111010110011;
    W_hn[3][13] = 21'b111111111110110011001;
    W_hn[3][14] = 21'b111111111111001011100;
    W_hn[3][15] = 21'b000000000001001110101;
    W_hn[4][0] = 21'b000000000000000011100;
    W_hn[4][1] = 21'b000000000000001001101;
    W_hn[4][2] = 21'b000000000000001111101;
    W_hn[4][3] = 21'b111111111111010111001;
    W_hn[4][4] = 21'b000000000001000110001;
    W_hn[4][5] = 21'b000000000001001011011;
    W_hn[4][6] = 21'b000000000001001010110;
    W_hn[4][7] = 21'b111111111110110110001;
    W_hn[4][8] = 21'b000000000000111111100;
    W_hn[4][9] = 21'b000000000001000111111;
    W_hn[4][10] = 21'b111111111111011111011;
    W_hn[4][11] = 21'b111111111111011000111;
    W_hn[4][12] = 21'b000000000000011111010;
    W_hn[4][13] = 21'b000000000000101000000;
    W_hn[4][14] = 21'b000000000001011010000;
    W_hn[4][15] = 21'b111111111111000011010;
    W_hn[5][0] = 21'b000000000000110111000;
    W_hn[5][1] = 21'b000000000000011100101;
    W_hn[5][2] = 21'b111111111111101011000;
    W_hn[5][3] = 21'b000000000000100000101;
    W_hn[5][4] = 21'b000000000001101000010;
    W_hn[5][5] = 21'b111111111110011110010;
    W_hn[5][6] = 21'b000000000000000001101;
    W_hn[5][7] = 21'b000000000001000111110;
    W_hn[5][8] = 21'b000000000000110110011;
    W_hn[5][9] = 21'b000000000000000001011;
    W_hn[5][10] = 21'b111111111110000010100;
    W_hn[5][11] = 21'b000000000001110001111;
    W_hn[5][12] = 21'b000000000001011111110;
    W_hn[5][13] = 21'b000000000000100010111;
    W_hn[5][14] = 21'b111111111110110100110;
    W_hn[5][15] = 21'b000000000010100101111;
    W_hn[6][0] = 21'b111111111111110101110;
    W_hn[6][1] = 21'b111111111111101100110;
    W_hn[6][2] = 21'b000000000000100100011;
    W_hn[6][3] = 21'b111111111111001100011;
    W_hn[6][4] = 21'b111111111111010010111;
    W_hn[6][5] = 21'b111111111111111001111;
    W_hn[6][6] = 21'b000000000010111011100;
    W_hn[6][7] = 21'b111111111110100010001;
    W_hn[6][8] = 21'b111111111111110101110;
    W_hn[6][9] = 21'b000000000001101100111;
    W_hn[6][10] = 21'b000000000010011111001;
    W_hn[6][11] = 21'b111111111110010000010;
    W_hn[6][12] = 21'b111111111111010110011;
    W_hn[6][13] = 21'b111111111110110011001;
    W_hn[6][14] = 21'b111111111111001011100;
    W_hn[6][15] = 21'b000000000001001110101;
    W_hn[7][0] = 21'b000000000000000011100;
    W_hn[7][1] = 21'b000000000000001001101;
    W_hn[7][2] = 21'b000000000000001111101;
    W_hn[7][3] = 21'b111111111111010111001;
    W_hn[7][4] = 21'b000000000001000110001;
    W_hn[7][5] = 21'b000000000001001011011;
    W_hn[7][6] = 21'b000000000001001010110;
    W_hn[7][7] = 21'b111111111110110110001;
    W_hn[7][8] = 21'b000000000000111111100;
    W_hn[7][9] = 21'b000000000001000111111;
    W_hn[7][10] = 21'b111111111111011111011;
    W_hn[7][11] = 21'b111111111111011000111;
    W_hn[7][12] = 21'b000000000000011111010;
    W_hn[7][13] = 21'b000000000000101000000;
    W_hn[7][14] = 21'b000000000001011010000;
    W_hn[7][15] = 21'b111111111111000011010;
    W_hn[8][0] = 21'b000000000000110111000;
    W_hn[8][1] = 21'b000000000000011100101;
    W_hn[8][2] = 21'b111111111111101011000;
    W_hn[8][3] = 21'b000000000000100000101;
    W_hn[8][4] = 21'b000000000001101000010;
    W_hn[8][5] = 21'b111111111110011110010;
    W_hn[8][6] = 21'b000000000000000001101;
    W_hn[8][7] = 21'b000000000001000111110;
    W_hn[8][8] = 21'b000000000000110110011;
    W_hn[8][9] = 21'b000000000000000001011;
    W_hn[8][10] = 21'b111111111110000010100;
    W_hn[8][11] = 21'b000000000001110001111;
    W_hn[8][12] = 21'b000000000001011111110;
    W_hn[8][13] = 21'b000000000000100010111;
    W_hn[8][14] = 21'b111111111110110100110;
    W_hn[8][15] = 21'b000000000010100101111;
    W_hn[9][0] = 21'b111111111111110101110;
    W_hn[9][1] = 21'b111111111111101100110;
    W_hn[9][2] = 21'b000000000000100100011;
    W_hn[9][3] = 21'b111111111111001100011;
    W_hn[9][4] = 21'b111111111111010010111;
    W_hn[9][5] = 21'b111111111111111001111;
    W_hn[9][6] = 21'b000000000010111011100;
    W_hn[9][7] = 21'b111111111110100010001;
    W_hn[9][8] = 21'b111111111111110101110;
    W_hn[9][9] = 21'b000000000001101100111;
    W_hn[9][10] = 21'b000000000010011111001;
    W_hn[9][11] = 21'b111111111110010000010;
    W_hn[9][12] = 21'b111111111111010110011;
    W_hn[9][13] = 21'b111111111110110011001;
    W_hn[9][14] = 21'b111111111111001011100;
    W_hn[9][15] = 21'b000000000001001110101;
    W_hn[10][0] = 21'b000000000000000011100;
    W_hn[10][1] = 21'b000000000000001001101;
    W_hn[10][2] = 21'b000000000000001111101;
    W_hn[10][3] = 21'b111111111111010111001;
    W_hn[10][4] = 21'b000000000001000110001;
    W_hn[10][5] = 21'b000000000001001011011;
    W_hn[10][6] = 21'b000000000001001010110;
    W_hn[10][7] = 21'b111111111110110110001;
    W_hn[10][8] = 21'b000000000000111111100;
    W_hn[10][9] = 21'b000000000001000111111;
    W_hn[10][10] = 21'b111111111111011111011;
    W_hn[10][11] = 21'b111111111111011000111;
    W_hn[10][12] = 21'b000000000000011111010;
    W_hn[10][13] = 21'b000000000000101000000;
    W_hn[10][14] = 21'b000000000001011010000;
    W_hn[10][15] = 21'b111111111111000011010;
    W_hn[11][0] = 21'b000000000000110111000;
    W_hn[11][1] = 21'b000000000000011100101;
    W_hn[11][2] = 21'b111111111111101011000;
    W_hn[11][3] = 21'b000000000000100000101;
    W_hn[11][4] = 21'b000000000001101000010;
    W_hn[11][5] = 21'b111111111110011110010;
    W_hn[11][6] = 21'b000000000000000001101;
    W_hn[11][7] = 21'b000000000001000111110;
    W_hn[11][8] = 21'b000000000000110110011;
    W_hn[11][9] = 21'b000000000000000001011;
    W_hn[11][10] = 21'b111111111110000010100;
    W_hn[11][11] = 21'b000000000001110001111;
    W_hn[11][12] = 21'b000000000001011111110;
    W_hn[11][13] = 21'b000000000000100010111;
    W_hn[11][14] = 21'b111111111110110100110;
    W_hn[11][15] = 21'b000000000010100101111;
    W_hn[12][0] = 21'b111111111111110101110;
    W_hn[12][1] = 21'b111111111111101100110;
    W_hn[12][2] = 21'b000000000000100100011;
    W_hn[12][3] = 21'b111111111111001100011;
    W_hn[12][4] = 21'b111111111111010010111;
    W_hn[12][5] = 21'b111111111111111001111;
    W_hn[12][6] = 21'b000000000010111011100;
    W_hn[12][7] = 21'b111111111110100010001;
    W_hn[12][8] = 21'b111111111111110101110;
    W_hn[12][9] = 21'b000000000001101100111;
    W_hn[12][10] = 21'b000000000010011111001;
    W_hn[12][11] = 21'b111111111110010000010;
    W_hn[12][12] = 21'b111111111111010110011;
    W_hn[12][13] = 21'b111111111110110011001;
    W_hn[12][14] = 21'b111111111111001011100;
    W_hn[12][15] = 21'b000000000001001110101;
    W_hn[13][0] = 21'b000000000000000011100;
    W_hn[13][1] = 21'b000000000000001001101;
    W_hn[13][2] = 21'b000000000000001111101;
    W_hn[13][3] = 21'b111111111111010111001;
    W_hn[13][4] = 21'b000000000001000110001;
    W_hn[13][5] = 21'b000000000001001011011;
    W_hn[13][6] = 21'b000000000001001010110;
    W_hn[13][7] = 21'b111111111110110110001;
    W_hn[13][8] = 21'b000000000000111111100;
    W_hn[13][9] = 21'b000000000001000111111;
    W_hn[13][10] = 21'b111111111111011111011;
    W_hn[13][11] = 21'b111111111111011000111;
    W_hn[13][12] = 21'b000000000000011111010;
    W_hn[13][13] = 21'b000000000000101000000;
    W_hn[13][14] = 21'b000000000001011010000;
    W_hn[13][15] = 21'b111111111111000011010;
    W_hn[14][0] = 21'b000000000000110111000;
    W_hn[14][1] = 21'b000000000000011100101;
    W_hn[14][2] = 21'b111111111111101011000;
    W_hn[14][3] = 21'b000000000000100000101;
    W_hn[14][4] = 21'b000000000001101000010;
    W_hn[14][5] = 21'b111111111110011110010;
    W_hn[14][6] = 21'b000000000000000001101;
    W_hn[14][7] = 21'b000000000001000111110;
    W_hn[14][8] = 21'b000000000000110110011;
    W_hn[14][9] = 21'b000000000000000001011;
    W_hn[14][10] = 21'b111111111110000010100;
    W_hn[14][11] = 21'b000000000001110001111;
    W_hn[14][12] = 21'b000000000001011111110;
    W_hn[14][13] = 21'b000000000000100010111;
    W_hn[14][14] = 21'b111111111110110100110;
    W_hn[14][15] = 21'b000000000010100101111;
    W_hn[15][0] = 21'b111111111111110101110;
    W_hn[15][1] = 21'b111111111111101100110;
    W_hn[15][2] = 21'b000000000000100100011;
    W_hn[15][3] = 21'b111111111111001100011;
    W_hn[15][4] = 21'b111111111111010010111;
    W_hn[15][5] = 21'b111111111111111001111;
    W_hn[15][6] = 21'b000000000010111011100;
    W_hn[15][7] = 21'b111111111110100010001;
    W_hn[15][8] = 21'b111111111111110101110;
    W_hn[15][9] = 21'b000000000001101100111;
    W_hn[15][10] = 21'b000000000010011111001;
    W_hn[15][11] = 21'b111111111110010000010;
    W_hn[15][12] = 21'b111111111111010110011;
    W_hn[15][13] = 21'b111111111110110011001;
    W_hn[15][14] = 21'b111111111111001011100;
    W_hn[15][15] = 21'b000000000001001110101;

    // Initialize biases

    // Initialize b_ir biases
    b_ir[0] = 21'b000000000000000101110;
    b_ir[1] = 21'b000000000001000010110;
    b_ir[2] = 21'b000000000001110110110;
    b_ir[3] = 21'b000000000000101000111;
    b_ir[4] = 21'b000000000000110000101;
    b_ir[5] = 21'b000000000000100010011;
    b_ir[6] = 21'b000000000001111110001;
    b_ir[7] = 21'b111111111111111101000;
    b_ir[8] = 21'b000000000001010101000;
    b_ir[9] = 21'b000000000000001110100;
    b_ir[10] = 21'b000000000001110000100;
    b_ir[11] = 21'b000000000000010011000;
    b_ir[12] = 21'b000000000000010010010;
    b_ir[13] = 21'b000000000001001110010;
    b_ir[14] = 21'b000000000000110111000;
    b_ir[15] = 21'b000000000001101000110;

    // Initialize b_iz biases
    b_iz[0] = 21'b000000000000110100010;
    b_iz[1] = 21'b000000000001001001010;
    b_iz[2] = 21'b000000000000100111111;
    b_iz[3] = 21'b000000000011001110110;
    b_iz[4] = 21'b000000000000011000010;
    b_iz[5] = 21'b000000000010010111111;
    b_iz[6] = 21'b000000000000111010100;
    b_iz[7] = 21'b111111111110000100001;
    b_iz[8] = 21'b000000000000000101110;
    b_iz[9] = 21'b000000000001000010110;
    b_iz[10] = 21'b000000000001110110110;
    b_iz[11] = 21'b000000000000101000111;
    b_iz[12] = 21'b000000000000110000101;
    b_iz[13] = 21'b000000000000100010011;
    b_iz[14] = 21'b000000000001111110001;
    b_iz[15] = 21'b111111111111111101000;

    // Initialize b_in biases
    b_in[0] = 21'b000000000001010101000;
    b_in[1] = 21'b000000000000001110100;
    b_in[2] = 21'b000000000001110000100;
    b_in[3] = 21'b000000000000010011000;
    b_in[4] = 21'b000000000000010010010;
    b_in[5] = 21'b000000000001001110010;
    b_in[6] = 21'b000000000000110111000;
    b_in[7] = 21'b000000000001101000110;
    b_in[8] = 21'b000000000000110100010;
    b_in[9] = 21'b000000000001001001010;
    b_in[10] = 21'b000000000000100111111;
    b_in[11] = 21'b000000000011001110110;
    b_in[12] = 21'b000000000000011000010;
    b_in[13] = 21'b000000000010010111111;
    b_in[14] = 21'b000000000000111010100;
    b_in[15] = 21'b111111111110000100001;

    // Initialize b_hr biases
    b_hr[0] = 21'b000000000000000101110;
    b_hr[1] = 21'b000000000001000010110;
    b_hr[2] = 21'b000000000001110110110;
    b_hr[3] = 21'b000000000000101000111;
    b_hr[4] = 21'b000000000000110000101;
    b_hr[5] = 21'b000000000000100010011;
    b_hr[6] = 21'b000000000001111110001;
    b_hr[7] = 21'b111111111111111101000;
    b_hr[8] = 21'b000000000001010101000;
    b_hr[9] = 21'b000000000000001110100;
    b_hr[10] = 21'b000000000001110000100;
    b_hr[11] = 21'b000000000000010011000;
    b_hr[12] = 21'b000000000000010010010;
    b_hr[13] = 21'b000000000001001110010;
    b_hr[14] = 21'b000000000000110111000;
    b_hr[15] = 21'b000000000001101000110;

    // Initialize b_hz biases
    b_hz[0] = 21'b000000000000110100010;
    b_hz[1] = 21'b000000000001001001010;
    b_hz[2] = 21'b000000000000100111111;
    b_hz[3] = 21'b000000000011001110110;
    b_hz[4] = 21'b000000000000011000010;
    b_hz[5] = 21'b000000000010010111111;
    b_hz[6] = 21'b000000000000111010100;
    b_hz[7] = 21'b111111111110000100001;
    b_hz[8] = 21'b000000000000000101110;
    b_hz[9] = 21'b000000000001000010110;
    b_hz[10] = 21'b000000000001110110110;
    b_hz[11] = 21'b000000000000101000111;
    b_hz[12] = 21'b000000000000110000101;
    b_hz[13] = 21'b000000000000100010011;
    b_hz[14] = 21'b000000000001111110001;
    b_hz[15] = 21'b111111111111111101000;

    // Initialize b_hn biases
    b_hn[0] = 21'b000000000001010101000;
    b_hn[1] = 21'b000000000000001110100;
    b_hn[2] = 21'b000000000001110000100;
    b_hn[3] = 21'b000000000000010011000;
    b_hn[4] = 21'b000000000000010010010;
    b_hn[5] = 21'b000000000001001110010;
    b_hn[6] = 21'b000000000000110111000;
    b_hn[7] = 21'b000000000001101000110;
    b_hn[8] = 21'b000000000000110100010;
    b_hn[9] = 21'b000000000001001001010;
    b_hn[10] = 21'b000000000000100111111;
    b_hn[11] = 21'b000000000011001110110;
    b_hn[12] = 21'b000000000000011000010;
    b_hn[13] = 21'b000000000010010111111;
    b_hn[14] = 21'b000000000000111010100;
    b_hn[15] = 21'b111111111110000100001;

    // Reset sequence
    rst_n = 0;
    start = 0;
    test_start_cycle = 0;
    test_cycles = 0;
    total_cycles = 0;
    test_timeout = 0;
    repeat(10) @(posedge clk);
    rst_n = 1;
    repeat(5) @(posedge clk);

    // Test Vector 1
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000100100010010;
        x_t[1] = 21'b000000000110110110001;
        x_t[2] = 21'b000000001000001001010;
        x_t[3] = 21'b000000001001000110100;
        x_t[4] = 21'b000000000111010100111;
        x_t[5] = 21'b000000000110101110001;
        x_t[6] = 21'b000000000100111010001;
        x_t[7] = 21'b000000000100100111110;
        x_t[8] = 21'b000000000111100001010;
        x_t[9] = 21'b000000001001000010001;
        x_t[10] = 21'b000000001001011010011;
        x_t[11] = 21'b000000001001001001001;
        x_t[12] = 21'b000000001000111011000;
        x_t[13] = 21'b000000000101100100011;
        x_t[14] = 21'b000000000111010101111;
        x_t[15] = 21'b000000001000110010000;
        x_t[16] = 21'b000000001001001111010;
        x_t[17] = 21'b000000001001100111110;
        x_t[18] = 21'b000000001001111011011;
        x_t[19] = 21'b000000001001101100010;
        x_t[20] = 21'b000000000110110111110;
        x_t[21] = 21'b000000000010000100100;
        x_t[22] = 21'b000000000010011110110;
        x_t[23] = 21'b000000000010111011101;
        x_t[24] = 21'b000000000001011101010;
        x_t[25] = 21'b000000000001110011010;
        x_t[26] = 21'b000000000101000100101;
        x_t[27] = 21'b000000000011011101110;
        x_t[28] = 21'b000000000011101111101;
        x_t[29] = 21'b000000000001011100010;
        x_t[30] = 21'b000000000010111101001;
        x_t[31] = 21'b000000000110001110100;
        x_t[32] = 21'b000000000111101101010;
        x_t[33] = 21'b000000000111110000011;
        x_t[34] = 21'b000000000110111110010;
        x_t[35] = 21'b000000000101111010000;
        x_t[36] = 21'b000000000100111100101;
        x_t[37] = 21'b000000000010100100000;
        x_t[38] = 21'b000000000010111001111;
        x_t[39] = 21'b000000000100011100111;
        x_t[40] = 21'b000000000101010011111;
        x_t[41] = 21'b000000000110100011010;
        x_t[42] = 21'b000000000100000011010;
        x_t[43] = 21'b000000000011011000000;
        x_t[44] = 21'b000000000110000101010;
        x_t[45] = 21'b000000000010111001010;
        x_t[46] = 21'b000000000111010100010;
        x_t[47] = 21'b000000001000010110000;
        x_t[48] = 21'b000000000111111011111;
        x_t[49] = 21'b000000001000101100010;
        x_t[50] = 21'b000000001010001001011;
        x_t[51] = 21'b000000001010101011010;
        x_t[52] = 21'b000000001010000110111;
        x_t[53] = 21'b000000001000110000110;
        x_t[54] = 21'b000000000110110100100;
        x_t[55] = 21'b000000000110110101100;
        x_t[56] = 21'b000000001000010110000;
        x_t[57] = 21'b000000001000110000100;
        x_t[58] = 21'b000000001001000111111;
        x_t[59] = 21'b000000000101110110010;
        x_t[60] = 21'b000000000101111110100;
        x_t[61] = 21'b000000000110011001001;
        x_t[62] = 21'b000000000100101011000;
        x_t[63] = 21'b000000000101111111001;
        
        h_t_prev[0] = 21'b000000000100100010010;
        h_t_prev[1] = 21'b000000000110110110001;
        h_t_prev[2] = 21'b000000001000001001010;
        h_t_prev[3] = 21'b000000001001000110100;
        h_t_prev[4] = 21'b000000000111010100111;
        h_t_prev[5] = 21'b000000000110101110001;
        h_t_prev[6] = 21'b000000000100111010001;
        h_t_prev[7] = 21'b000000000100100111110;
        h_t_prev[8] = 21'b000000000111100001010;
        h_t_prev[9] = 21'b000000001001000010001;
        h_t_prev[10] = 21'b000000001001011010011;
        h_t_prev[11] = 21'b000000001001001001001;
        h_t_prev[12] = 21'b000000001000111011000;
        h_t_prev[13] = 21'b000000000101100100011;
        h_t_prev[14] = 21'b000000000111010101111;
        h_t_prev[15] = 21'b000000001000110010000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 1 timeout!");
                $fdisplay(fd_cycles, "Test Vector   1: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   1: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 1");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 2
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000101110001010;
        x_t[1] = 21'b000000001001001001000;
        x_t[2] = 21'b000000001010001100011;
        x_t[3] = 21'b000000001010101100000;
        x_t[4] = 21'b000000001001111011101;
        x_t[5] = 21'b000000001001011111101;
        x_t[6] = 21'b000000000111111011001;
        x_t[7] = 21'b000000000110110110010;
        x_t[8] = 21'b000000001010001011100;
        x_t[9] = 21'b000000001011001110011;
        x_t[10] = 21'b000000001011010100101;
        x_t[11] = 21'b000000001011110110011;
        x_t[12] = 21'b000000001011010011010;
        x_t[13] = 21'b000000001000000001001;
        x_t[14] = 21'b000000001001101001100;
        x_t[15] = 21'b000000001010110110010;
        x_t[16] = 21'b000000001011000001010;
        x_t[17] = 21'b000000001011101000001;
        x_t[18] = 21'b000000001011101111011;
        x_t[19] = 21'b000000001011100101001;
        x_t[20] = 21'b000000001000011011111;
        x_t[21] = 21'b000000000010010101000;
        x_t[22] = 21'b000000000010011110110;
        x_t[23] = 21'b000000000010110010111;
        x_t[24] = 21'b000000000011000001110;
        x_t[25] = 21'b000000000011001101011;
        x_t[26] = 21'b000000000101100110100;
        x_t[27] = 21'b000000000100001001000;
        x_t[28] = 21'b000000000011010011011;
        x_t[29] = 21'b000000000100010111100;
        x_t[30] = 21'b000000000101001101100;
        x_t[31] = 21'b000000000111000011110;
        x_t[32] = 21'b000000001000010001100;
        x_t[33] = 21'b000000000111111110010;
        x_t[34] = 21'b000000000111001100101;
        x_t[35] = 21'b000000000110100110100;
        x_t[36] = 21'b000000000101001011101;
        x_t[37] = 21'b000000000011001000101;
        x_t[38] = 21'b000000000110100110111;
        x_t[39] = 21'b000000000010101110101;
        x_t[40] = 21'b000000001000010010001;
        x_t[41] = 21'b111111111111100110001;
        x_t[42] = 21'b000000000111010010110;
        x_t[43] = 21'b000000000100100100110;
        x_t[44] = 21'b000000001000111101101;
        x_t[45] = 21'b000000000000100110010;
        x_t[46] = 21'b000000001001000110001;
        x_t[47] = 21'b000000001001000111101;
        x_t[48] = 21'b000000001000000000101;
        x_t[49] = 21'b000000001000000111010;
        x_t[50] = 21'b000000001001101100111;
        x_t[51] = 21'b000000001010001110011;
        x_t[52] = 21'b000000001001001001100;
        x_t[53] = 21'b000000000111011101010;
        x_t[54] = 21'b000000000101001110101;
        x_t[55] = 21'b000000000110100100010;
        x_t[56] = 21'b000000000111101111010;
        x_t[57] = 21'b000000000111110000101;
        x_t[58] = 21'b000000001000010011100;
        x_t[59] = 21'b000000000101000110111;
        x_t[60] = 21'b000000000101110011000;
        x_t[61] = 21'b000000000110011101010;
        x_t[62] = 21'b000000000100110010011;
        x_t[63] = 21'b000000000101101001001;
        
        h_t_prev[0] = 21'b000000000101110001010;
        h_t_prev[1] = 21'b000000001001001001000;
        h_t_prev[2] = 21'b000000001010001100011;
        h_t_prev[3] = 21'b000000001010101100000;
        h_t_prev[4] = 21'b000000001001111011101;
        h_t_prev[5] = 21'b000000001001011111101;
        h_t_prev[6] = 21'b000000000111111011001;
        h_t_prev[7] = 21'b000000000110110110010;
        h_t_prev[8] = 21'b000000001010001011100;
        h_t_prev[9] = 21'b000000001011001110011;
        h_t_prev[10] = 21'b000000001011010100101;
        h_t_prev[11] = 21'b000000001011110110011;
        h_t_prev[12] = 21'b000000001011010011010;
        h_t_prev[13] = 21'b000000001000000001001;
        h_t_prev[14] = 21'b000000001001101001100;
        h_t_prev[15] = 21'b000000001010110110010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 2 timeout!");
                $fdisplay(fd_cycles, "Test Vector   2: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   2: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 2");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 3
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000111111011011;
        x_t[1] = 21'b000000001000011000000;
        x_t[2] = 21'b000000001000000100011;
        x_t[3] = 21'b000000000111111110000;
        x_t[4] = 21'b000000000110110110100;
        x_t[5] = 21'b000000000101100110000;
        x_t[6] = 21'b000000000011101111100;
        x_t[7] = 21'b000000000110001101100;
        x_t[8] = 21'b000000001000001111101;
        x_t[9] = 21'b000000001000001011000;
        x_t[10] = 21'b000000001000000010010;
        x_t[11] = 21'b000000001000011011011;
        x_t[12] = 21'b000000000110100010111;
        x_t[13] = 21'b000000000001101111001;
        x_t[14] = 21'b000000001000000101011;
        x_t[15] = 21'b000000001000010011100;
        x_t[16] = 21'b000000001000000100111;
        x_t[17] = 21'b000000001000011000111;
        x_t[18] = 21'b000000001000000111100;
        x_t[19] = 21'b000000000111011101100;
        x_t[20] = 21'b000000000011101001010;
        x_t[21] = 21'b000000000100001001001;
        x_t[22] = 21'b000000000011001110011;
        x_t[23] = 21'b000000000010111011101;
        x_t[24] = 21'b000000000101100000000;
        x_t[25] = 21'b000000000101101000110;
        x_t[26] = 21'b000000000100011110101;
        x_t[27] = 21'b000000000011011101110;
        x_t[28] = 21'b000000000010111101010;
        x_t[29] = 21'b000000000111011011000;
        x_t[30] = 21'b000000000101011001001;
        x_t[31] = 21'b000000000101000111100;
        x_t[32] = 21'b000000000110011011011;
        x_t[33] = 21'b000000000101101110111;
        x_t[34] = 21'b000000000100110100001;
        x_t[35] = 21'b000000000100001101100;
        x_t[36] = 21'b000000000011001010011;
        x_t[37] = 21'b000000000010010011101;
        x_t[38] = 21'b000000000110011100110;
        x_t[39] = 21'b000000000000001101000;
        x_t[40] = 21'b000000000111000000101;
        x_t[41] = 21'b000000000000001000111;
        x_t[42] = 21'b000000000110101111010;
        x_t[43] = 21'b000000000100001110110;
        x_t[44] = 21'b000000000111011110101;
        x_t[45] = 21'b000000000000011110100;
        x_t[46] = 21'b000000000111001111000;
        x_t[47] = 21'b000000000110110111100;
        x_t[48] = 21'b000000000101011001111;
        x_t[49] = 21'b000000000101100000011;
        x_t[50] = 21'b000000000111000001111;
        x_t[51] = 21'b000000000111011011101;
        x_t[52] = 21'b000000000110011011101;
        x_t[53] = 21'b000000000101010111101;
        x_t[54] = 21'b000000000100001100110;
        x_t[55] = 21'b000000000100101011011;
        x_t[56] = 21'b000000000101111111101;
        x_t[57] = 21'b000000000101110000101;
        x_t[58] = 21'b000000000110101010110;
        x_t[59] = 21'b000000000100101011010;
        x_t[60] = 21'b000000000100110001111;
        x_t[61] = 21'b000000000101110011111;
        x_t[62] = 21'b000000000100010001001;
        x_t[63] = 21'b000000000101110001111;
        
        h_t_prev[0] = 21'b000000000111111011011;
        h_t_prev[1] = 21'b000000001000011000000;
        h_t_prev[2] = 21'b000000001000000100011;
        h_t_prev[3] = 21'b000000000111111110000;
        h_t_prev[4] = 21'b000000000110110110100;
        h_t_prev[5] = 21'b000000000101100110000;
        h_t_prev[6] = 21'b000000000011101111100;
        h_t_prev[7] = 21'b000000000110001101100;
        h_t_prev[8] = 21'b000000001000001111101;
        h_t_prev[9] = 21'b000000001000001011000;
        h_t_prev[10] = 21'b000000001000000010010;
        h_t_prev[11] = 21'b000000001000011011011;
        h_t_prev[12] = 21'b000000000110100010111;
        h_t_prev[13] = 21'b000000000001101111001;
        h_t_prev[14] = 21'b000000001000000101011;
        h_t_prev[15] = 21'b000000001000010011100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 3 timeout!");
                $fdisplay(fd_cycles, "Test Vector   3: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   3: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 3");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 4
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000101100111011;
        x_t[1] = 21'b000000000101111011011;
        x_t[2] = 21'b000000000110100011010;
        x_t[3] = 21'b000000000111001101101;
        x_t[4] = 21'b000000000110000100000;
        x_t[5] = 21'b000000000100100011011;
        x_t[6] = 21'b000000000011011100111;
        x_t[7] = 21'b000000000011110100111;
        x_t[8] = 21'b000000000110000100011;
        x_t[9] = 21'b000000000110101011110;
        x_t[10] = 21'b000000000110111101110;
        x_t[11] = 21'b000000000111011110001;
        x_t[12] = 21'b000000000101010110110;
        x_t[13] = 21'b000000000010001010011;
        x_t[14] = 21'b000000000101110001101;
        x_t[15] = 21'b000000000110101101111;
        x_t[16] = 21'b000000000110100110110;
        x_t[17] = 21'b000000000110110001010;
        x_t[18] = 21'b000000000110111000011;
        x_t[19] = 21'b000000000110010000101;
        x_t[20] = 21'b000000000011011100110;
        x_t[21] = 21'b000000000011011010001;
        x_t[22] = 21'b000000000011001011001;
        x_t[23] = 21'b000000000011110101101;
        x_t[24] = 21'b000000000100000001101;
        x_t[25] = 21'b000000000100010001110;
        x_t[26] = 21'b000000000100110011110;
        x_t[27] = 21'b000000000100010000110;
        x_t[28] = 21'b000000000100011110111;
        x_t[29] = 21'b000000000100001011000;
        x_t[30] = 21'b000000000011111011100;
        x_t[31] = 21'b000000000101000011001;
        x_t[32] = 21'b000000000110000100110;
        x_t[33] = 21'b000000000110000001011;
        x_t[34] = 21'b000000000101011111000;
        x_t[35] = 21'b000000000100100110001;
        x_t[36] = 21'b000000000100011001111;
        x_t[37] = 21'b000000000011011001000;
        x_t[38] = 21'b000000000011100010010;
        x_t[39] = 21'b000000000011100010001;
        x_t[40] = 21'b000000000110000100111;
        x_t[41] = 21'b000000000101100100101;
        x_t[42] = 21'b000000000100001001010;
        x_t[43] = 21'b000000000001101010010;
        x_t[44] = 21'b000000000100010000000;
        x_t[45] = 21'b000000000001111011011;
        x_t[46] = 21'b000000000100011001110;
        x_t[47] = 21'b000000000101000101001;
        x_t[48] = 21'b000000000100010111001;
        x_t[49] = 21'b000000000100011111100;
        x_t[50] = 21'b000000000101100010111;
        x_t[51] = 21'b000000000101110001011;
        x_t[52] = 21'b000000000100111010011;
        x_t[53] = 21'b000000000100011111111;
        x_t[54] = 21'b000000000011111010110;
        x_t[55] = 21'b000000000011101010101;
        x_t[56] = 21'b000000000100111010111;
        x_t[57] = 21'b000000000100111001010;
        x_t[58] = 21'b000000000101100000101;
        x_t[59] = 21'b000000000100001011101;
        x_t[60] = 21'b000000000011101001000;
        x_t[61] = 21'b000000000100110101110;
        x_t[62] = 21'b000000000011010010010;
        x_t[63] = 21'b000000000101101101100;
        
        h_t_prev[0] = 21'b000000000101100111011;
        h_t_prev[1] = 21'b000000000101111011011;
        h_t_prev[2] = 21'b000000000110100011010;
        h_t_prev[3] = 21'b000000000111001101101;
        h_t_prev[4] = 21'b000000000110000100000;
        h_t_prev[5] = 21'b000000000100100011011;
        h_t_prev[6] = 21'b000000000011011100111;
        h_t_prev[7] = 21'b000000000011110100111;
        h_t_prev[8] = 21'b000000000110000100011;
        h_t_prev[9] = 21'b000000000110101011110;
        h_t_prev[10] = 21'b000000000110111101110;
        h_t_prev[11] = 21'b000000000111011110001;
        h_t_prev[12] = 21'b000000000101010110110;
        h_t_prev[13] = 21'b000000000010001010011;
        h_t_prev[14] = 21'b000000000101110001101;
        h_t_prev[15] = 21'b000000000110101101111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 4 timeout!");
                $fdisplay(fd_cycles, "Test Vector   4: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   4: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 4");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 5
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000011100010001;
        x_t[1] = 21'b000000000100101101001;
        x_t[2] = 21'b000000000101001011111;
        x_t[3] = 21'b000000000110001001111;
        x_t[4] = 21'b000000000101100000101;
        x_t[5] = 21'b000000000100000010001;
        x_t[6] = 21'b000000000011101001010;
        x_t[7] = 21'b000000000010100011011;
        x_t[8] = 21'b000000000100001000101;
        x_t[9] = 21'b000000000100111000100;
        x_t[10] = 21'b000000000101010010001;
        x_t[11] = 21'b000000000110000010100;
        x_t[12] = 21'b000000000100000100110;
        x_t[13] = 21'b000000000001111100110;
        x_t[14] = 21'b000000000100010010110;
        x_t[15] = 21'b000000000101000011000;
        x_t[16] = 21'b000000000100111110101;
        x_t[17] = 21'b000000000100111111110;
        x_t[18] = 21'b000000000100111001111;
        x_t[19] = 21'b000000000100001100110;
        x_t[20] = 21'b000000000010010001101;
        x_t[21] = 21'b000000000011110101110;
        x_t[22] = 21'b000000000010101000010;
        x_t[23] = 21'b000000000011011000101;
        x_t[24] = 21'b000000000010101100011;
        x_t[25] = 21'b000000000010110100100;
        x_t[26] = 21'b000000000100000001001;
        x_t[27] = 21'b000000000011101001100;
        x_t[28] = 21'b000000000011111001001;
        x_t[29] = 21'b000000000001110001001;
        x_t[30] = 21'b000000000011001000110;
        x_t[31] = 21'b000000000100001001100;
        x_t[32] = 21'b000000000100111100000;
        x_t[33] = 21'b000000000100110010110;
        x_t[34] = 21'b000000000100100101111;
        x_t[35] = 21'b000000000011010111010;
        x_t[36] = 21'b000000000011001111011;
        x_t[37] = 21'b000000000010011111111;
        x_t[38] = 21'b000000000001011111001;
        x_t[39] = 21'b000000000001101100100;
        x_t[40] = 21'b000000000000110011111;
        x_t[41] = 21'b000000000001100011010;
        x_t[42] = 21'b000000000000011100000;
        x_t[43] = 21'b111111111111011011101;
        x_t[44] = 21'b000000000010001001111;
        x_t[45] = 21'b000000000000011110100;
        x_t[46] = 21'b000000000011101011001;
        x_t[47] = 21'b000000000100100010010;
        x_t[48] = 21'b000000000011100111100;
        x_t[49] = 21'b000000000011110101111;
        x_t[50] = 21'b000000000100100101000;
        x_t[51] = 21'b000000000100101000111;
        x_t[52] = 21'b000000000011101000100;
        x_t[53] = 21'b000000000011010010000;
        x_t[54] = 21'b000000000010011010111;
        x_t[55] = 21'b000000000011010000110;
        x_t[56] = 21'b000000000100011100110;
        x_t[57] = 21'b000000000100011011011;
        x_t[58] = 21'b000000000100101000000;
        x_t[59] = 21'b000000000011001100100;
        x_t[60] = 21'b000000000011000010101;
        x_t[61] = 21'b000000000100000100001;
        x_t[62] = 21'b000000000010010011011;
        x_t[63] = 21'b000000000101010011001;
        
        h_t_prev[0] = 21'b000000000011100010001;
        h_t_prev[1] = 21'b000000000100101101001;
        h_t_prev[2] = 21'b000000000101001011111;
        h_t_prev[3] = 21'b000000000110001001111;
        h_t_prev[4] = 21'b000000000101100000101;
        h_t_prev[5] = 21'b000000000100000010001;
        h_t_prev[6] = 21'b000000000011101001010;
        h_t_prev[7] = 21'b000000000010100011011;
        h_t_prev[8] = 21'b000000000100001000101;
        h_t_prev[9] = 21'b000000000100111000100;
        h_t_prev[10] = 21'b000000000101010010001;
        h_t_prev[11] = 21'b000000000110000010100;
        h_t_prev[12] = 21'b000000000100000100110;
        h_t_prev[13] = 21'b000000000001111100110;
        h_t_prev[14] = 21'b000000000100010010110;
        h_t_prev[15] = 21'b000000000101000011000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 5 timeout!");
                $fdisplay(fd_cycles, "Test Vector   5: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   5: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 5");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 6
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000010011000010;
        x_t[1] = 21'b000000000011110111010;
        x_t[2] = 21'b000000000100100000001;
        x_t[3] = 21'b000000000101011110011;
        x_t[4] = 21'b000000000100101001001;
        x_t[5] = 21'b000000000010110100100;
        x_t[6] = 21'b000000000010100100111;
        x_t[7] = 21'b000000000001010111001;
        x_t[8] = 21'b000000000011100100100;
        x_t[9] = 21'b000000000100101001100;
        x_t[10] = 21'b000000000101000011100;
        x_t[11] = 21'b000000000101111000010;
        x_t[12] = 21'b000000000011110011010;
        x_t[13] = 21'b000000000001101000010;
        x_t[14] = 21'b000000000011111101101;
        x_t[15] = 21'b000000000100111000111;
        x_t[16] = 21'b000000000100111001110;
        x_t[17] = 21'b000000000101001001101;
        x_t[18] = 21'b000000000100110100101;
        x_t[19] = 21'b000000000100100010110;
        x_t[20] = 21'b000000000010100100100;
        x_t[21] = 21'b000000000010011010100;
        x_t[22] = 21'b000000000010000010001;
        x_t[23] = 21'b000000000010010000001;
        x_t[24] = 21'b000000000010010001000;
        x_t[25] = 21'b000000000010010101011;
        x_t[26] = 21'b000000000011001110011;
        x_t[27] = 21'b000000000010011010111;
        x_t[28] = 21'b000000000010010111100;
        x_t[29] = 21'b000000000001100000011;
        x_t[30] = 21'b000000000011101011111;
        x_t[31] = 21'b000000000011101110111;
        x_t[32] = 21'b000000000100111100000;
        x_t[33] = 21'b000000000100100100111;
        x_t[34] = 21'b000000000100000100100;
        x_t[35] = 21'b000000000011001101011;
        x_t[36] = 21'b000000000010011101101;
        x_t[37] = 21'b000000000001100110110;
        x_t[38] = 21'b000000000001010101000;
        x_t[39] = 21'b000000000001000111110;
        x_t[40] = 21'b000000000010001010111;
        x_t[41] = 21'b000000000000101011101;
        x_t[42] = 21'b000000000010101010011;
        x_t[43] = 21'b000000000011011000000;
        x_t[44] = 21'b000000000011001101000;
        x_t[45] = 21'b000000000001001100111;
        x_t[46] = 21'b000000000011001100000;
        x_t[47] = 21'b000000000011101011100;
        x_t[48] = 21'b000000000010101001101;
        x_t[49] = 21'b000000000011011110101;
        x_t[50] = 21'b000000000100100101000;
        x_t[51] = 21'b000000000101000101111;
        x_t[52] = 21'b000000000100100000110;
        x_t[53] = 21'b000000000100101011000;
        x_t[54] = 21'b000000000011010110110;
        x_t[55] = 21'b000000000010001011110;
        x_t[56] = 21'b000000000011011100010;
        x_t[57] = 21'b000000000011111001010;
        x_t[58] = 21'b000000000100110101000;
        x_t[59] = 21'b000000000011001000100;
        x_t[60] = 21'b000000000010100000001;
        x_t[61] = 21'b000000000011010110101;
        x_t[62] = 21'b000000000001011000001;
        x_t[63] = 21'b000000000100010101100;
        
        h_t_prev[0] = 21'b000000000010011000010;
        h_t_prev[1] = 21'b000000000011110111010;
        h_t_prev[2] = 21'b000000000100100000001;
        h_t_prev[3] = 21'b000000000101011110011;
        h_t_prev[4] = 21'b000000000100101001001;
        h_t_prev[5] = 21'b000000000010110100100;
        h_t_prev[6] = 21'b000000000010100100111;
        h_t_prev[7] = 21'b000000000001010111001;
        h_t_prev[8] = 21'b000000000011100100100;
        h_t_prev[9] = 21'b000000000100101001100;
        h_t_prev[10] = 21'b000000000101000011100;
        h_t_prev[11] = 21'b000000000101111000010;
        h_t_prev[12] = 21'b000000000011110011010;
        h_t_prev[13] = 21'b000000000001101000010;
        h_t_prev[14] = 21'b000000000011111101101;
        h_t_prev[15] = 21'b000000000100111000111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 6 timeout!");
                $fdisplay(fd_cycles, "Test Vector   6: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   6: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 6");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 7
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000011000100101;
        x_t[1] = 21'b000000000100101000010;
        x_t[2] = 21'b000000000101011111010;
        x_t[3] = 21'b000000000110100111000;
        x_t[4] = 21'b000000000101110100111;
        x_t[5] = 21'b000000000100010010110;
        x_t[6] = 21'b000000000011100011000;
        x_t[7] = 21'b000000000000110011100;
        x_t[8] = 21'b000000000100000011100;
        x_t[9] = 21'b000000000101010110101;
        x_t[10] = 21'b000000000110001000000;
        x_t[11] = 21'b000000000111010100000;
        x_t[12] = 21'b000000000101110100000;
        x_t[13] = 21'b000000000011100010111;
        x_t[14] = 21'b000000000010011001100;
        x_t[15] = 21'b000000000100100100100;
        x_t[16] = 21'b000000000101000011101;
        x_t[17] = 21'b000000000101010011100;
        x_t[18] = 21'b000000000101101110101;
        x_t[19] = 21'b000000000110010000101;
        x_t[20] = 21'b000000000101000111001;
        x_t[21] = 21'b000000000010000100100;
        x_t[22] = 21'b000000000001110101100;
        x_t[23] = 21'b000000000001111000111;
        x_t[24] = 21'b000000000010110010100;
        x_t[25] = 21'b000000000010110111101;
        x_t[26] = 21'b000000000011101100000;
        x_t[27] = 21'b000000000010110010100;
        x_t[28] = 21'b000000000010010001010;
        x_t[29] = 21'b000000000010001010000;
        x_t[30] = 21'b000000000100011110101;
        x_t[31] = 21'b000000000100010110110;
        x_t[32] = 21'b000000000101010010110;
        x_t[33] = 21'b000000000101001110100;
        x_t[34] = 21'b000000000100101111011;
        x_t[35] = 21'b000000000100000011101;
        x_t[36] = 21'b000000000011101000010;
        x_t[37] = 21'b000000000010011111111;
        x_t[38] = 21'b000000000010011011101;
        x_t[39] = 21'b000000000010011000101;
        x_t[40] = 21'b000000000100000010011;
        x_t[41] = 21'b000000000010011011000;
        x_t[42] = 21'b000000000010101010011;
        x_t[43] = 21'b000000001001001101000;
        x_t[44] = 21'b000000000011000111011;
        x_t[45] = 21'b000000000100000110101;
        x_t[46] = 21'b000000000010011000001;
        x_t[47] = 21'b000000000010101010111;
        x_t[48] = 21'b000000000001101011101;
        x_t[49] = 21'b000000000010100010100;
        x_t[50] = 21'b000000000100010110110;
        x_t[51] = 21'b000000000101100111110;
        x_t[52] = 21'b000000000101110111110;
        x_t[53] = 21'b000000000110011010011;
        x_t[54] = 21'b000000000101111000101;
        x_t[55] = 21'b000000000001000110101;
        x_t[56] = 21'b000000000010100100100;
        x_t[57] = 21'b000000000011010111010;
        x_t[58] = 21'b000000000101100101000;
        x_t[59] = 21'b000000000011111111111;
        x_t[60] = 21'b000000000001101110011;
        x_t[61] = 21'b000000000010011100101;
        x_t[62] = 21'b000000000000110110111;
        x_t[63] = 21'b000000000010111101100;
        
        h_t_prev[0] = 21'b000000000011000100101;
        h_t_prev[1] = 21'b000000000100101000010;
        h_t_prev[2] = 21'b000000000101011111010;
        h_t_prev[3] = 21'b000000000110100111000;
        h_t_prev[4] = 21'b000000000101110100111;
        h_t_prev[5] = 21'b000000000100010010110;
        h_t_prev[6] = 21'b000000000011100011000;
        h_t_prev[7] = 21'b000000000000110011100;
        h_t_prev[8] = 21'b000000000100000011100;
        h_t_prev[9] = 21'b000000000101010110101;
        h_t_prev[10] = 21'b000000000110001000000;
        h_t_prev[11] = 21'b000000000111010100000;
        h_t_prev[12] = 21'b000000000101110100000;
        h_t_prev[13] = 21'b000000000011100010111;
        h_t_prev[14] = 21'b000000000010011001100;
        h_t_prev[15] = 21'b000000000100100100100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 7 timeout!");
                $fdisplay(fd_cycles, "Test Vector   7: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   7: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 7");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 8
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000011000100101;
        x_t[1] = 21'b000000000100010100101;
        x_t[2] = 21'b000000000101001011111;
        x_t[3] = 21'b000000000110101011110;
        x_t[4] = 21'b000000000110001001001;
        x_t[5] = 21'b000000000100111001101;
        x_t[6] = 21'b000000000100101101110;
        x_t[7] = 21'b000000000001000111111;
        x_t[8] = 21'b000000000011011111011;
        x_t[9] = 21'b000000000100100100100;
        x_t[10] = 21'b000000000101101111100;
        x_t[11] = 21'b000000000111010100000;
        x_t[12] = 21'b000000000110010111001;
        x_t[13] = 21'b000000000100110100110;
        x_t[14] = 21'b000000000010010100001;
        x_t[15] = 21'b000000000100000000111;
        x_t[16] = 21'b000000000100010010000;
        x_t[17] = 21'b000000000100110000111;
        x_t[18] = 21'b000000000101101110101;
        x_t[19] = 21'b000000000110100001001;
        x_t[20] = 21'b000000000101111111100;
        x_t[21] = 21'b000000000010110011011;
        x_t[22] = 21'b000000000010001110111;
        x_t[23] = 21'b000000000010100111010;
        x_t[24] = 21'b000000000010110010100;
        x_t[25] = 21'b000000000010111101111;
        x_t[26] = 21'b000000000100000101011;
        x_t[27] = 21'b000000000011011001110;
        x_t[28] = 21'b000000000011000000100;
        x_t[29] = 21'b000000000010001010000;
        x_t[30] = 21'b000000000100001011001;
        x_t[31] = 21'b000000000100110001011;
        x_t[32] = 21'b000000000101010111010;
        x_t[33] = 21'b000000000101001001111;
        x_t[34] = 21'b000000000100110100001;
        x_t[35] = 21'b000000000100001000100;
        x_t[36] = 21'b000000000100010100111;
        x_t[37] = 21'b000000000011011101000;
        x_t[38] = 21'b000000000001100100001;
        x_t[39] = 21'b000000000010111101011;
        x_t[40] = 21'b000000000011000001001;
        x_t[41] = 21'b000000000011000100101;
        x_t[42] = 21'b000000000001101111000;
        x_t[43] = 21'b000000000101010000101;
        x_t[44] = 21'b000000000001101110000;
        x_t[45] = 21'b000000000100011101111;
        x_t[46] = 21'b000000000001101001100;
        x_t[47] = 21'b000000000010010010000;
        x_t[48] = 21'b000000000001011000101;
        x_t[49] = 21'b000000000010010100100;
        x_t[50] = 21'b000000000100001000100;
        x_t[51] = 21'b000000000101011110000;
        x_t[52] = 21'b000000000101011001001;
        x_t[53] = 21'b000000000110000100001;
        x_t[54] = 21'b000000000101001110101;
        x_t[55] = 21'b000000000001001011000;
        x_t[56] = 21'b000000000010100000001;
        x_t[57] = 21'b000000000011010011000;
        x_t[58] = 21'b000000000100111101110;
        x_t[59] = 21'b000000000010111000110;
        x_t[60] = 21'b000000000001001000000;
        x_t[61] = 21'b000000000001101111001;
        x_t[62] = 21'b000000000000011001010;
        x_t[63] = 21'b000000000001011100101;
        
        h_t_prev[0] = 21'b000000000011000100101;
        h_t_prev[1] = 21'b000000000100010100101;
        h_t_prev[2] = 21'b000000000101001011111;
        h_t_prev[3] = 21'b000000000110101011110;
        h_t_prev[4] = 21'b000000000110001001001;
        h_t_prev[5] = 21'b000000000100111001101;
        h_t_prev[6] = 21'b000000000100101101110;
        h_t_prev[7] = 21'b000000000001000111111;
        h_t_prev[8] = 21'b000000000011011111011;
        h_t_prev[9] = 21'b000000000100100100100;
        h_t_prev[10] = 21'b000000000101101111100;
        h_t_prev[11] = 21'b000000000111010100000;
        h_t_prev[12] = 21'b000000000110010111001;
        h_t_prev[13] = 21'b000000000100110100110;
        h_t_prev[14] = 21'b000000000010010100001;
        h_t_prev[15] = 21'b000000000100000000111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 8 timeout!");
                $fdisplay(fd_cycles, "Test Vector   8: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   8: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 8");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 9
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000010111010110;
        x_t[1] = 21'b000000000011101101100;
        x_t[2] = 21'b000000000100101110110;
        x_t[3] = 21'b000000000101111011011;
        x_t[4] = 21'b000000000101011011101;
        x_t[5] = 21'b000000000100011101111;
        x_t[6] = 21'b000000000100101101110;
        x_t[7] = 21'b000000000000101110011;
        x_t[8] = 21'b000000000010100110101;
        x_t[9] = 21'b000000000011101000011;
        x_t[10] = 21'b000000000100101011000;
        x_t[11] = 21'b000000000110100001000;
        x_t[12] = 21'b000000000101100010100;
        x_t[13] = 21'b000000000101001001001;
        x_t[14] = 21'b000000000001101111010;
        x_t[15] = 21'b000000000011000011111;
        x_t[16] = 21'b000000000011011011100;
        x_t[17] = 21'b000000000100001001011;
        x_t[18] = 21'b000000000100110100101;
        x_t[19] = 21'b000000000101011111001;
        x_t[20] = 21'b000000000101000000111;
        x_t[21] = 21'b000000000011010111011;
        x_t[22] = 21'b000000000010010101010;
        x_t[23] = 21'b000000000010110010111;
        x_t[24] = 21'b000000000011001010111;
        x_t[25] = 21'b000000000011011001110;
        x_t[26] = 21'b000000000100001001100;
        x_t[27] = 21'b000000000011001110000;
        x_t[28] = 21'b000000000010001110001;
        x_t[29] = 21'b000000000010010110100;
        x_t[30] = 21'b000000000100001011001;
        x_t[31] = 21'b000000000100010010011;
        x_t[32] = 21'b000000000101001001101;
        x_t[33] = 21'b000000000100101110001;
        x_t[34] = 21'b000000000100010111101;
        x_t[35] = 21'b000000000011110100110;
        x_t[36] = 21'b000000000011000101011;
        x_t[37] = 21'b000000000010110100010;
        x_t[38] = 21'b000000000010000010011;
        x_t[39] = 21'b000000000001101100100;
        x_t[40] = 21'b000000000010110110011;
        x_t[41] = 21'b000000000001101010010;
        x_t[42] = 21'b000000000001101111000;
        x_t[43] = 21'b000000000100100100110;
        x_t[44] = 21'b000000000000011010010;
        x_t[45] = 21'b000000000010000011001;
        x_t[46] = 21'b000000000010001101111;
        x_t[47] = 21'b000000000010101111111;
        x_t[48] = 21'b000000000001100010001;
        x_t[49] = 21'b000000000010100111001;
        x_t[50] = 21'b000000000011110000110;
        x_t[51] = 21'b000000000100110010101;
        x_t[52] = 21'b000000000100001100011;
        x_t[53] = 21'b000000000100011010011;
        x_t[54] = 21'b000000000011110100110;
        x_t[55] = 21'b000000000010101001111;
        x_t[56] = 21'b000000000011100100111;
        x_t[57] = 21'b000000000011110000110;
        x_t[58] = 21'b000000000100010110100;
        x_t[59] = 21'b000000000010001101011;
        x_t[60] = 21'b000000000001100110101;
        x_t[61] = 21'b000000000001110011010;
        x_t[62] = 21'b000000000000001010100;
        x_t[63] = 21'b000000000001011000010;
        
        h_t_prev[0] = 21'b000000000010111010110;
        h_t_prev[1] = 21'b000000000011101101100;
        h_t_prev[2] = 21'b000000000100101110110;
        h_t_prev[3] = 21'b000000000101111011011;
        h_t_prev[4] = 21'b000000000101011011101;
        h_t_prev[5] = 21'b000000000100011101111;
        h_t_prev[6] = 21'b000000000100101101110;
        h_t_prev[7] = 21'b000000000000101110011;
        h_t_prev[8] = 21'b000000000010100110101;
        h_t_prev[9] = 21'b000000000011101000011;
        h_t_prev[10] = 21'b000000000100101011000;
        h_t_prev[11] = 21'b000000000110100001000;
        h_t_prev[12] = 21'b000000000101100010100;
        h_t_prev[13] = 21'b000000000101001001001;
        h_t_prev[14] = 21'b000000000001101111010;
        h_t_prev[15] = 21'b000000000011000011111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 9 timeout!");
                $fdisplay(fd_cycles, "Test Vector   9: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   9: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 9");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 10
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000010001001011;
        x_t[1] = 21'b000000000010011010010;
        x_t[2] = 21'b000000000011001101101;
        x_t[3] = 21'b000000000100010001001;
        x_t[4] = 21'b000000000011110110101;
        x_t[5] = 21'b000000000010011000110;
        x_t[6] = 21'b000000000001110011000;
        x_t[7] = 21'b000000000001000010110;
        x_t[8] = 21'b000000000001111101011;
        x_t[9] = 21'b000000000010100010010;
        x_t[10] = 21'b000000000011010011000;
        x_t[11] = 21'b000000000100100110110;
        x_t[12] = 21'b000000000011010000001;
        x_t[13] = 21'b000000000001000110010;
        x_t[14] = 21'b000000000010010100001;
        x_t[15] = 21'b000000000011001110000;
        x_t[16] = 21'b000000000011000111110;
        x_t[17] = 21'b000000000011010011001;
        x_t[18] = 21'b000000000011010101110;
        x_t[19] = 21'b000000000011100000111;
        x_t[20] = 21'b000000000010011000000;
        x_t[21] = 21'b000000000010100000001;
        x_t[22] = 21'b000000000001011111010;
        x_t[23] = 21'b000000000001110110000;
        x_t[24] = 21'b000000000001100110011;
        x_t[25] = 21'b000000000001110110011;
        x_t[26] = 21'b000000000010011011110;
        x_t[27] = 21'b000000000001101011110;
        x_t[28] = 21'b000000000010000100101;
        x_t[29] = 21'b000000000000111011000;
        x_t[30] = 21'b000000000010010110000;
        x_t[31] = 21'b000000000001111011100;
        x_t[32] = 21'b000000000010101111010;
        x_t[33] = 21'b000000000010011010001;
        x_t[34] = 21'b000000000010000100000;
        x_t[35] = 21'b000000000001001000001;
        x_t[36] = 21'b000000000000001101100;
        x_t[37] = 21'b000000000001001010010;
        x_t[38] = 21'b000000000000111011111;
        x_t[39] = 21'b111111111111010010001;
        x_t[40] = 21'b000000000001001001101;
        x_t[41] = 21'b111111111111100110001;
        x_t[42] = 21'b000000000001100011001;
        x_t[43] = 21'b000000000100011001110;
        x_t[44] = 21'b000000000011000001110;
        x_t[45] = 21'b000000000010011010010;
        x_t[46] = 21'b000000000101010010101;
        x_t[47] = 21'b000000000100010011011;
        x_t[48] = 21'b000000000010010110100;
        x_t[49] = 21'b000000000011011010000;
        x_t[50] = 21'b000000000011100111010;
        x_t[51] = 21'b000000000011111000101;
        x_t[52] = 21'b000000000011001001111;
        x_t[53] = 21'b000000000011011101001;
        x_t[54] = 21'b000000000011011100110;
        x_t[55] = 21'b000000000100010101110;
        x_t[56] = 21'b000000000101010000011;
        x_t[57] = 21'b000000000100010010111;
        x_t[58] = 21'b000000000100000101000;
        x_t[59] = 21'b000000000010101001000;
        x_t[60] = 21'b000000000011000010101;
        x_t[61] = 21'b000000000011000110000;
        x_t[62] = 21'b000000000000110011010;
        x_t[63] = 21'b000000000011000110010;
        
        h_t_prev[0] = 21'b000000000010001001011;
        h_t_prev[1] = 21'b000000000010011010010;
        h_t_prev[2] = 21'b000000000011001101101;
        h_t_prev[3] = 21'b000000000100010001001;
        h_t_prev[4] = 21'b000000000011110110101;
        h_t_prev[5] = 21'b000000000010011000110;
        h_t_prev[6] = 21'b000000000001110011000;
        h_t_prev[7] = 21'b000000000001000010110;
        h_t_prev[8] = 21'b000000000001111101011;
        h_t_prev[9] = 21'b000000000010100010010;
        h_t_prev[10] = 21'b000000000011010011000;
        h_t_prev[11] = 21'b000000000100100110110;
        h_t_prev[12] = 21'b000000000011010000001;
        h_t_prev[13] = 21'b000000000001000110010;
        h_t_prev[14] = 21'b000000000010010100001;
        h_t_prev[15] = 21'b000000000011001110000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 10 timeout!");
                $fdisplay(fd_cycles, "Test Vector  10: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  10: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 10");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 11
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000000110000101;
        x_t[1] = 21'b000000000000111000011;
        x_t[2] = 21'b000000000001010100010;
        x_t[3] = 21'b000000000010000100111;
        x_t[4] = 21'b000000000001101001001;
        x_t[5] = 21'b111111111111111101011;
        x_t[6] = 21'b111111111111011101101;
        x_t[7] = 21'b111111111111111011100;
        x_t[8] = 21'b000000000001100011101;
        x_t[9] = 21'b000000000001110101001;
        x_t[10] = 21'b000000000010001001101;
        x_t[11] = 21'b000000000010001101111;
        x_t[12] = 21'b000000000001011011000;
        x_t[13] = 21'b111111111111100000000;
        x_t[14] = 21'b000000000011000011101;
        x_t[15] = 21'b000000000011100010011;
        x_t[16] = 21'b000000000011000010110;
        x_t[17] = 21'b000000000010110101100;
        x_t[18] = 21'b000000000010001011111;
        x_t[19] = 21'b000000000010001001000;
        x_t[20] = 21'b000000000001011001011;
        x_t[21] = 21'b000000000000111001111;
        x_t[22] = 21'b000000000000010011001;
        x_t[23] = 21'b000000000000110000011;
        x_t[24] = 21'b000000000000111000110;
        x_t[25] = 21'b000000000001000001100;
        x_t[26] = 21'b000000000000100001010;
        x_t[27] = 21'b111111111111101110000;
        x_t[28] = 21'b000000000000111001000;
        x_t[29] = 21'b000000000000010101100;
        x_t[30] = 21'b000000000001110110111;
        x_t[31] = 21'b000000000000110000001;
        x_t[32] = 21'b000000000001100110100;
        x_t[33] = 21'b000000000001000010010;
        x_t[34] = 21'b000000000000011011001;
        x_t[35] = 21'b111111111111101111010;
        x_t[36] = 21'b111111111110101111001;
        x_t[37] = 21'b111111111111111100110;
        x_t[38] = 21'b000000000001101110010;
        x_t[39] = 21'b111111111110010111011;
        x_t[40] = 21'b000000000011101100101;
        x_t[41] = 21'b000000000010001101000;
        x_t[42] = 21'b000000000100001001010;
        x_t[43] = 21'b000000000000110011011;
        x_t[44] = 21'b000000000100110111001;
        x_t[45] = 21'b000000000001111011011;
        x_t[46] = 21'b000000000101100111011;
        x_t[47] = 21'b000000000101000101001;
        x_t[48] = 21'b000000000010110111111;
        x_t[49] = 21'b000000000011110101111;
        x_t[50] = 21'b000000000011011101110;
        x_t[51] = 21'b000000000011010110111;
        x_t[52] = 21'b000000000010100000111;
        x_t[53] = 21'b000000000011000001010;
        x_t[54] = 21'b000000000011010000110;
        x_t[55] = 21'b000000000101011010111;
        x_t[56] = 21'b000000000110000011111;
        x_t[57] = 21'b000000000100101100100;
        x_t[58] = 21'b000000000011110011101;
        x_t[59] = 21'b000000000010101100111;
        x_t[60] = 21'b000000000100101110000;
        x_t[61] = 21'b000000000100100101010;
        x_t[62] = 21'b000000000001100011010;
        x_t[63] = 21'b000000000101010011001;
        
        h_t_prev[0] = 21'b000000000000110000101;
        h_t_prev[1] = 21'b000000000000111000011;
        h_t_prev[2] = 21'b000000000001010100010;
        h_t_prev[3] = 21'b000000000010000100111;
        h_t_prev[4] = 21'b000000000001101001001;
        h_t_prev[5] = 21'b111111111111111101011;
        h_t_prev[6] = 21'b111111111111011101101;
        h_t_prev[7] = 21'b111111111111111011100;
        h_t_prev[8] = 21'b000000000001100011101;
        h_t_prev[9] = 21'b000000000001110101001;
        h_t_prev[10] = 21'b000000000010001001101;
        h_t_prev[11] = 21'b000000000010001101111;
        h_t_prev[12] = 21'b000000000001011011000;
        h_t_prev[13] = 21'b111111111111100000000;
        h_t_prev[14] = 21'b000000000011000011101;
        h_t_prev[15] = 21'b000000000011100010011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 11 timeout!");
                $fdisplay(fd_cycles, "Test Vector  11: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  11: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 11");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 12
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000010100111000;
        x_t[1] = 21'b000000000010000001110;
        x_t[2] = 21'b000000000001111111111;
        x_t[3] = 21'b000000000010000100111;
        x_t[4] = 21'b000000000001100100001;
        x_t[5] = 21'b111111111111100111010;
        x_t[6] = 21'b111111111111010111100;
        x_t[7] = 21'b000000000001101011100;
        x_t[8] = 21'b000000000010011100011;
        x_t[9] = 21'b000000000010001001001;
        x_t[10] = 21'b000000000001110001001;
        x_t[11] = 21'b000000000001111001100;
        x_t[12] = 21'b000000000000110010001;
        x_t[13] = 21'b111111111111011001001;
        x_t[14] = 21'b000000000100000010111;
        x_t[15] = 21'b000000000011111011111;
        x_t[16] = 21'b000000000010111101110;
        x_t[17] = 21'b000000000010001001001;
        x_t[18] = 21'b000000000001010111010;
        x_t[19] = 21'b000000000001100010100;
        x_t[20] = 21'b000000000000101101101;
        x_t[21] = 21'b000000000001011000010;
        x_t[22] = 21'b000000000000011111110;
        x_t[23] = 21'b000000000000011100000;
        x_t[24] = 21'b000000000001100011011;
        x_t[25] = 21'b000000000001101001111;
        x_t[26] = 21'b000000000000110010001;
        x_t[27] = 21'b111111111111110101111;
        x_t[28] = 21'b000000000000100011000;
        x_t[29] = 21'b000000000001111101100;
        x_t[30] = 21'b000000000010001010011;
        x_t[31] = 21'b000000000000110100100;
        x_t[32] = 21'b000000000010001111011;
        x_t[33] = 21'b000000000001110000100;
        x_t[34] = 21'b000000000000111100100;
        x_t[35] = 21'b000000000000010110110;
        x_t[36] = 21'b111111111111000011000;
        x_t[37] = 21'b000000000000001101001;
        x_t[38] = 21'b000000000010010110101;
        x_t[39] = 21'b111111111101110010101;
        x_t[40] = 21'b000000000100110011011;
        x_t[41] = 21'b111111111111000011011;
        x_t[42] = 21'b000000000101101000000;
        x_t[43] = 21'b111111111101001101000;
        x_t[44] = 21'b000000000100111100101;
        x_t[45] = 21'b111111111111111111100;
        x_t[46] = 21'b000000000101001101100;
        x_t[47] = 21'b000000000101000101001;
        x_t[48] = 21'b000000000010110111111;
        x_t[49] = 21'b000000000011011010000;
        x_t[50] = 21'b000000000010110011000;
        x_t[51] = 21'b000000000010100001110;
        x_t[52] = 21'b000000000001010100001;
        x_t[53] = 21'b000000000001101101110;
        x_t[54] = 21'b000000000001011110111;
        x_t[55] = 21'b000000000101010010010;
        x_t[56] = 21'b000000000101110010110;
        x_t[57] = 21'b000000000100011011011;
        x_t[58] = 21'b000000000010110010001;
        x_t[59] = 21'b000000000001010010001;
        x_t[60] = 21'b000000000101010100011;
        x_t[61] = 21'b000000000101000010001;
        x_t[62] = 21'b000000000001011111101;
        x_t[63] = 21'b000000000101111010110;
        
        h_t_prev[0] = 21'b000000000010100111000;
        h_t_prev[1] = 21'b000000000010000001110;
        h_t_prev[2] = 21'b000000000001111111111;
        h_t_prev[3] = 21'b000000000010000100111;
        h_t_prev[4] = 21'b000000000001100100001;
        h_t_prev[5] = 21'b111111111111100111010;
        h_t_prev[6] = 21'b111111111111010111100;
        h_t_prev[7] = 21'b000000000001101011100;
        h_t_prev[8] = 21'b000000000010011100011;
        h_t_prev[9] = 21'b000000000010001001001;
        h_t_prev[10] = 21'b000000000001110001001;
        h_t_prev[11] = 21'b000000000001111001100;
        h_t_prev[12] = 21'b000000000000110010001;
        h_t_prev[13] = 21'b111111111111011001001;
        h_t_prev[14] = 21'b000000000100000010111;
        h_t_prev[15] = 21'b000000000011111011111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 12 timeout!");
                $fdisplay(fd_cycles, "Test Vector  12: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  12: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 12");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 13
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000010101011111;
        x_t[1] = 21'b000000000010010000100;
        x_t[2] = 21'b000000000010001001101;
        x_t[3] = 21'b000000000010001110101;
        x_t[4] = 21'b000000000001001111111;
        x_t[5] = 21'b111111111111000101111;
        x_t[6] = 21'b111111111110111110100;
        x_t[7] = 21'b000000000001111111110;
        x_t[8] = 21'b000000000010010010000;
        x_t[9] = 21'b000000000001110000001;
        x_t[10] = 21'b000000000001100111011;
        x_t[11] = 21'b000000000001100101001;
        x_t[12] = 21'b111111111111111101011;
        x_t[13] = 21'b111111111110001110010;
        x_t[14] = 21'b000000000011111101101;
        x_t[15] = 21'b000000000011011101011;
        x_t[16] = 21'b000000000010100000000;
        x_t[17] = 21'b000000000001100001101;
        x_t[18] = 21'b000000000001000111011;
        x_t[19] = 21'b000000000001000111001;
        x_t[20] = 21'b000000000000000001110;
        x_t[21] = 21'b000000000001100000100;
        x_t[22] = 21'b000000000000000110011;
        x_t[23] = 21'b000000000000010000100;
        x_t[24] = 21'b000000000001111000101;
        x_t[25] = 21'b000000000010000010110;
        x_t[26] = 21'b000000000000011101000;
        x_t[27] = 21'b111111111111110001111;
        x_t[28] = 21'b000000000000011111111;
        x_t[29] = 21'b000000000010101111100;
        x_t[30] = 21'b000000000001011011100;
        x_t[31] = 21'b000000000000110000001;
        x_t[32] = 21'b000000000001111000101;
        x_t[33] = 21'b000000000001001011100;
        x_t[34] = 21'b000000000000011011001;
        x_t[35] = 21'b111111111111100000100;
        x_t[36] = 21'b111111111110110100000;
        x_t[37] = 21'b000000000000010001010;
        x_t[38] = 21'b000000000011000100000;
        x_t[39] = 21'b111111111100110111111;
        x_t[40] = 21'b000000000101011001011;
        x_t[41] = 21'b111111111100001110100;
        x_t[42] = 21'b000000000100101100110;
        x_t[43] = 21'b000000000101111100100;
        x_t[44] = 21'b000000000100110111001;
        x_t[45] = 21'b111111111111101000011;
        x_t[46] = 21'b000000000100101001010;
        x_t[47] = 21'b000000000100001110011;
        x_t[48] = 21'b000000000010001101000;
        x_t[49] = 21'b000000000011000010111;
        x_t[50] = 21'b000000000010101001100;
        x_t[51] = 21'b000000000010011000000;
        x_t[52] = 21'b000000000001001111001;
        x_t[53] = 21'b000000000001010111100;
        x_t[54] = 21'b000000000000100011000;
        x_t[55] = 21'b000000000011101010101;
        x_t[56] = 21'b000000000100100001000;
        x_t[57] = 21'b000000000011100100000;
        x_t[58] = 21'b000000000010000010010;
        x_t[59] = 21'b000000000000001111000;
        x_t[60] = 21'b000000000100100010100;
        x_t[61] = 21'b000000000100000100001;
        x_t[62] = 21'b000000000000011101000;
        x_t[63] = 21'b000000000011111111100;
        
        h_t_prev[0] = 21'b000000000010101011111;
        h_t_prev[1] = 21'b000000000010010000100;
        h_t_prev[2] = 21'b000000000010001001101;
        h_t_prev[3] = 21'b000000000010001110101;
        h_t_prev[4] = 21'b000000000001001111111;
        h_t_prev[5] = 21'b111111111111000101111;
        h_t_prev[6] = 21'b111111111110111110100;
        h_t_prev[7] = 21'b000000000001111111110;
        h_t_prev[8] = 21'b000000000010010010000;
        h_t_prev[9] = 21'b000000000001110000001;
        h_t_prev[10] = 21'b000000000001100111011;
        h_t_prev[11] = 21'b000000000001100101001;
        h_t_prev[12] = 21'b111111111111111101011;
        h_t_prev[13] = 21'b111111111110001110010;
        h_t_prev[14] = 21'b000000000011111101101;
        h_t_prev[15] = 21'b000000000011011101011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 13 timeout!");
                $fdisplay(fd_cycles, "Test Vector  13: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  13: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 13");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 14
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000001111010101;
        x_t[1] = 21'b000000000000101110101;
        x_t[2] = 21'b000000000001000000110;
        x_t[3] = 21'b000000000001100111111;
        x_t[4] = 21'b111111111111101111111;
        x_t[5] = 21'b111111111101100111101;
        x_t[6] = 21'b111111111101101101101;
        x_t[7] = 21'b000000000000000101101;
        x_t[8] = 21'b000000000000110101010;
        x_t[9] = 21'b000000000000110100000;
        x_t[10] = 21'b000000000001000000001;
        x_t[11] = 21'b000000000000011101110;
        x_t[12] = 21'b111111111110101011100;
        x_t[13] = 21'b111111111101011110100;
        x_t[14] = 21'b000000000001111001111;
        x_t[15] = 21'b000000000001110111101;
        x_t[16] = 21'b000000000001000110111;
        x_t[17] = 21'b000000000000100110011;
        x_t[18] = 21'b000000000000010010110;
        x_t[19] = 21'b000000000000000101010;
        x_t[20] = 21'b111111111110110110110;
        x_t[21] = 21'b000000000000110100011;
        x_t[22] = 21'b111111111110100111010;
        x_t[23] = 21'b111111111110110110100;
        x_t[24] = 21'b000000000001011010010;
        x_t[25] = 21'b000000000001100011110;
        x_t[26] = 21'b111111111110011110010;
        x_t[27] = 21'b111111111101110000001;
        x_t[28] = 21'b111111111110111000000;
        x_t[29] = 21'b000000000001110001001;
        x_t[30] = 21'b000000000000101000110;
        x_t[31] = 21'b111111111111000101101;
        x_t[32] = 21'b000000000000011101111;
        x_t[33] = 21'b111111111111001010000;
        x_t[34] = 21'b111111111110010001000;
        x_t[35] = 21'b111111111101111000111;
        x_t[36] = 21'b111111111100101000111;
        x_t[37] = 21'b111111111110100111010;
        x_t[38] = 21'b000000000010101111110;
        x_t[39] = 21'b111111111011010000111;
        x_t[40] = 21'b000000000100100011000;
        x_t[41] = 21'b111111111101000110001;
        x_t[42] = 21'b000000000001011101010;
        x_t[43] = 21'b000000000101011011101;
        x_t[44] = 21'b000000000001111110110;
        x_t[45] = 21'b111111111011001010000;
        x_t[46] = 21'b000000000001110011111;
        x_t[47] = 21'b000000000001111001001;
        x_t[48] = 21'b000000000000010001001;
        x_t[49] = 21'b000000000001000101110;
        x_t[50] = 21'b000000000000110111100;
        x_t[51] = 21'b000000000000101001000;
        x_t[52] = 21'b111111111111011001011;
        x_t[53] = 21'b111111111111000001001;
        x_t[54] = 21'b111111111101010111010;
        x_t[55] = 21'b000000000001011100010;
        x_t[56] = 21'b000000000010011011111;
        x_t[57] = 21'b000000000001110101001;
        x_t[58] = 21'b000000000000001100011;
        x_t[59] = 21'b111111111110101100011;
        x_t[60] = 21'b000000000010100111111;
        x_t[61] = 21'b000000000010000011110;
        x_t[62] = 21'b111111111110100011000;
        x_t[63] = 21'b000000000001000010010;
        
        h_t_prev[0] = 21'b000000000001111010101;
        h_t_prev[1] = 21'b000000000000101110101;
        h_t_prev[2] = 21'b000000000001000000110;
        h_t_prev[3] = 21'b000000000001100111111;
        h_t_prev[4] = 21'b111111111111101111111;
        h_t_prev[5] = 21'b111111111101100111101;
        h_t_prev[6] = 21'b111111111101101101101;
        h_t_prev[7] = 21'b000000000000000101101;
        h_t_prev[8] = 21'b000000000000110101010;
        h_t_prev[9] = 21'b000000000000110100000;
        h_t_prev[10] = 21'b000000000001000000001;
        h_t_prev[11] = 21'b000000000000011101110;
        h_t_prev[12] = 21'b111111111110101011100;
        h_t_prev[13] = 21'b111111111101011110100;
        h_t_prev[14] = 21'b000000000001111001111;
        h_t_prev[15] = 21'b000000000001110111101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 14 timeout!");
                $fdisplay(fd_cycles, "Test Vector  14: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  14: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 14");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 15
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000010011101001;
        x_t[1] = 21'b000000000001011010101;
        x_t[2] = 21'b000000000001011001000;
        x_t[3] = 21'b000000000001101100110;
        x_t[4] = 21'b000000000000001001001;
        x_t[5] = 21'b111111111101110010110;
        x_t[6] = 21'b111111111100111011111;
        x_t[7] = 21'b000000000001101011100;
        x_t[8] = 21'b000000000001111101011;
        x_t[9] = 21'b000000000010000100001;
        x_t[10] = 21'b000000000010011000010;
        x_t[11] = 21'b000000000010001000110;
        x_t[12] = 21'b111111111111100110000;
        x_t[13] = 21'b111111111110000000101;
        x_t[14] = 21'b000000000010101001010;
        x_t[15] = 21'b000000000011001001000;
        x_t[16] = 21'b000000000010011011001;
        x_t[17] = 21'b000000000010001001001;
        x_t[18] = 21'b000000000001111100001;
        x_t[19] = 21'b000000000001101101100;
        x_t[20] = 21'b111111111111111011100;
        x_t[21] = 21'b000000000000011000110;
        x_t[22] = 21'b111111111110111010010;
        x_t[23] = 21'b111111111111010110100;
        x_t[24] = 21'b000000000001000100111;
        x_t[25] = 21'b000000000001010111010;
        x_t[26] = 21'b111111111111100110001;
        x_t[27] = 21'b111111111110011011011;
        x_t[28] = 21'b111111111111011010101;
        x_t[29] = 21'b000000000001111001011;
        x_t[30] = 21'b000000000000111000011;
        x_t[31] = 21'b000000000000100010110;
        x_t[32] = 21'b000000000010010011111;
        x_t[33] = 21'b000000000001010100110;
        x_t[34] = 21'b000000000000010001101;
        x_t[35] = 21'b111111111111101111010;
        x_t[36] = 21'b111111111110001100010;
        x_t[37] = 21'b000000000000110001110;
        x_t[38] = 21'b000000000011100010010;
        x_t[39] = 21'b111111111110000001010;
        x_t[40] = 21'b000000000100000010011;
        x_t[41] = 21'b000000000001011100011;
        x_t[42] = 21'b000000000011001000000;
        x_t[43] = 21'b000000000011011000000;
        x_t[44] = 21'b000000000010110110101;
        x_t[45] = 21'b000000000001011100011;
        x_t[46] = 21'b000000000011001100000;
        x_t[47] = 21'b000000000011100110101;
        x_t[48] = 21'b000000000010001000010;
        x_t[49] = 21'b000000000011010000110;
        x_t[50] = 21'b000000000011010100010;
        x_t[51] = 21'b000000000011001000011;
        x_t[52] = 21'b000000000010000111011;
        x_t[53] = 21'b000000000001111110100;
        x_t[54] = 21'b000000000001100100111;
        x_t[55] = 21'b000000000010111111100;
        x_t[56] = 21'b000000000100000111010;
        x_t[57] = 21'b000000000011101000010;
        x_t[58] = 21'b000000000010001111010;
        x_t[59] = 21'b000000000000100110110;
        x_t[60] = 21'b000000000010000101011;
        x_t[61] = 21'b000000000001110111011;
        x_t[62] = 21'b111111111110010111111;
        x_t[63] = 21'b000000000001000010010;
        
        h_t_prev[0] = 21'b000000000010011101001;
        h_t_prev[1] = 21'b000000000001011010101;
        h_t_prev[2] = 21'b000000000001011001000;
        h_t_prev[3] = 21'b000000000001101100110;
        h_t_prev[4] = 21'b000000000000001001001;
        h_t_prev[5] = 21'b111111111101110010110;
        h_t_prev[6] = 21'b111111111100111011111;
        h_t_prev[7] = 21'b000000000001101011100;
        h_t_prev[8] = 21'b000000000001111101011;
        h_t_prev[9] = 21'b000000000010000100001;
        h_t_prev[10] = 21'b000000000010011000010;
        h_t_prev[11] = 21'b000000000010001000110;
        h_t_prev[12] = 21'b111111111111100110000;
        h_t_prev[13] = 21'b111111111110000000101;
        h_t_prev[14] = 21'b000000000010101001010;
        h_t_prev[15] = 21'b000000000011001001000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 15 timeout!");
                $fdisplay(fd_cycles, "Test Vector  15: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  15: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 15");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 16
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000011010011011;
        x_t[1] = 21'b000000000011001011010;
        x_t[2] = 21'b000000000011011100001;
        x_t[3] = 21'b000000000011111101110;
        x_t[4] = 21'b000000000011000100001;
        x_t[5] = 21'b000000000000100100010;
        x_t[6] = 21'b111111111111101010001;
        x_t[7] = 21'b000000000010110111110;
        x_t[8] = 21'b000000000011101001110;
        x_t[9] = 21'b000000000011110010011;
        x_t[10] = 21'b000000000100010111100;
        x_t[11] = 21'b000000000100100001101;
        x_t[12] = 21'b000000000010111000110;
        x_t[13] = 21'b000000000001000110010;
        x_t[14] = 21'b000000000100100111111;
        x_t[15] = 21'b000000000100011111011;
        x_t[16] = 21'b000000000100010111000;
        x_t[17] = 21'b000000000100000100100;
        x_t[18] = 21'b000000000100000101001;
        x_t[19] = 21'b000000000011111100011;
        x_t[20] = 21'b000000000010011000000;
        x_t[21] = 21'b000000000000111111011;
        x_t[22] = 21'b000000000000000110011;
        x_t[23] = 21'b000000000000010011011;
        x_t[24] = 21'b000000000001001011000;
        x_t[25] = 21'b000000000001100011110;
        x_t[26] = 21'b000000000000111110110;
        x_t[27] = 21'b111111111111011110010;
        x_t[28] = 21'b000000000000000011100;
        x_t[29] = 21'b000000000001101100111;
        x_t[30] = 21'b000000000000110100100;
        x_t[31] = 21'b000000000001011000000;
        x_t[32] = 21'b000000000010101111010;
        x_t[33] = 21'b000000000010000011000;
        x_t[34] = 21'b000000000001001111100;
        x_t[35] = 21'b000000000000001100111;
        x_t[36] = 21'b111111111111000011000;
        x_t[37] = 21'b000000000001011010101;
        x_t[38] = 21'b000000000001101001010;
        x_t[39] = 21'b111111111111000011100;
        x_t[40] = 21'b000000000001111010100;
        x_t[41] = 21'b000000000001011100011;
        x_t[42] = 21'b000000000011001000000;
        x_t[43] = 21'b000000000011101101111;
        x_t[44] = 21'b000000000010101011100;
        x_t[45] = 21'b000000000010101001110;
        x_t[46] = 21'b000000000011110101011;
        x_t[47] = 21'b000000000100001110011;
        x_t[48] = 21'b000000000010001101000;
        x_t[49] = 21'b000000000011101100101;
        x_t[50] = 21'b000000000011110000110;
        x_t[51] = 21'b000000000011101010001;
        x_t[52] = 21'b000000000010110101011;
        x_t[53] = 21'b000000000010010100110;
        x_t[54] = 21'b000000000001010011000;
        x_t[55] = 21'b000000000011101010101;
        x_t[56] = 21'b000000000100100101011;
        x_t[57] = 21'b000000000100000001111;
        x_t[58] = 21'b000000000010110010001;
        x_t[59] = 21'b000000000000101110101;
        x_t[60] = 21'b000000000011001010011;
        x_t[61] = 21'b000000000011000110000;
        x_t[62] = 21'b111111111111110100011;
        x_t[63] = 21'b000000000010100111100;
        
        h_t_prev[0] = 21'b000000000011010011011;
        h_t_prev[1] = 21'b000000000011001011010;
        h_t_prev[2] = 21'b000000000011011100001;
        h_t_prev[3] = 21'b000000000011111101110;
        h_t_prev[4] = 21'b000000000011000100001;
        h_t_prev[5] = 21'b000000000000100100010;
        h_t_prev[6] = 21'b111111111111101010001;
        h_t_prev[7] = 21'b000000000010110111110;
        h_t_prev[8] = 21'b000000000011101001110;
        h_t_prev[9] = 21'b000000000011110010011;
        h_t_prev[10] = 21'b000000000100010111100;
        h_t_prev[11] = 21'b000000000100100001101;
        h_t_prev[12] = 21'b000000000010111000110;
        h_t_prev[13] = 21'b000000000001000110010;
        h_t_prev[14] = 21'b000000000100100111111;
        h_t_prev[15] = 21'b000000000100011111011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 16 timeout!");
                $fdisplay(fd_cycles, "Test Vector  16: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  16: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 16");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 17
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000000100110110;
        x_t[1] = 21'b000000000000111000011;
        x_t[2] = 21'b111111111100111111011;
        x_t[3] = 21'b111111111101111111111;
        x_t[4] = 21'b111111111101100111100;
        x_t[5] = 21'b111111111101000110011;
        x_t[6] = 21'b111111111110011111011;
        x_t[7] = 21'b000000000010001010000;
        x_t[8] = 21'b000000000000000110110;
        x_t[9] = 21'b111111111110100010101;
        x_t[10] = 21'b111111111101011111001;
        x_t[11] = 21'b111111111011110110001;
        x_t[12] = 21'b111111111100001101011;
        x_t[13] = 21'b111111111100101110111;
        x_t[14] = 21'b000000000011000011101;
        x_t[15] = 21'b000000000001000100110;
        x_t[16] = 21'b111111111110111100000;
        x_t[17] = 21'b111111111101111110101;
        x_t[18] = 21'b111111111011110110001;
        x_t[19] = 21'b111111111011111101101;
        x_t[20] = 21'b111111111101001100011;
        x_t[21] = 21'b111111111111110111100;
        x_t[22] = 21'b000000000000111100011;
        x_t[23] = 21'b000000000001010000010;
        x_t[24] = 21'b000000000000101100100;
        x_t[25] = 21'b000000000000100101100;
        x_t[26] = 21'b111111111110001001001;
        x_t[27] = 21'b111111111110111110110;
        x_t[28] = 21'b000000000001111000000;
        x_t[29] = 21'b000000000000011001110;
        x_t[30] = 21'b000000000010001110010;
        x_t[31] = 21'b111111111111101101101;
        x_t[32] = 21'b111111111111000111100;
        x_t[33] = 21'b111111111110101001101;
        x_t[34] = 21'b111111111110010101110;
        x_t[35] = 21'b111111111101101111000;
        x_t[36] = 21'b111111111111101111110;
        x_t[37] = 21'b111111111011000111000;
        x_t[38] = 21'b000000000001000101111;
        x_t[39] = 21'b000000000000100011000;
        x_t[40] = 21'b000000000010001010111;
        x_t[41] = 21'b000000000000111001101;
        x_t[42] = 21'b000000000011000010000;
        x_t[43] = 21'b111111111111110001100;
        x_t[44] = 21'b000000000011011101110;
        x_t[45] = 21'b111111111111111111100;
        x_t[46] = 21'b000000000011011011100;
        x_t[47] = 21'b000000000010101111111;
        x_t[48] = 21'b000000000001110000011;
        x_t[49] = 21'b000000000000101010000;
        x_t[50] = 21'b111111111110101001000;
        x_t[51] = 21'b111111111101111011001;
        x_t[52] = 21'b111111111110000111100;
        x_t[53] = 21'b111111111110111011101;
        x_t[54] = 21'b000000000001001101000;
        x_t[55] = 21'b000000000001110001110;
        x_t[56] = 21'b000000000010100100100;
        x_t[57] = 21'b111111111111010011001;
        x_t[58] = 21'b111111111111001011000;
        x_t[59] = 21'b000000000010101001000;
        x_t[60] = 21'b000000000000010110001;
        x_t[61] = 21'b111111111111010001111;
        x_t[62] = 21'b111111111111100101100;
        x_t[63] = 21'b000000000000111101111;
        
        h_t_prev[0] = 21'b000000000000100110110;
        h_t_prev[1] = 21'b000000000000111000011;
        h_t_prev[2] = 21'b111111111100111111011;
        h_t_prev[3] = 21'b111111111101111111111;
        h_t_prev[4] = 21'b111111111101100111100;
        h_t_prev[5] = 21'b111111111101000110011;
        h_t_prev[6] = 21'b111111111110011111011;
        h_t_prev[7] = 21'b000000000010001010000;
        h_t_prev[8] = 21'b000000000000000110110;
        h_t_prev[9] = 21'b111111111110100010101;
        h_t_prev[10] = 21'b111111111101011111001;
        h_t_prev[11] = 21'b111111111011110110001;
        h_t_prev[12] = 21'b111111111100001101011;
        h_t_prev[13] = 21'b111111111100101110111;
        h_t_prev[14] = 21'b000000000011000011101;
        h_t_prev[15] = 21'b000000000001000100110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 17 timeout!");
                $fdisplay(fd_cycles, "Test Vector  17: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  17: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 17");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 18
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000010100111000;
        x_t[1] = 21'b000000000011000001011;
        x_t[2] = 21'b000000000000000001101;
        x_t[3] = 21'b000000000000101001000;
        x_t[4] = 21'b111111111111101010111;
        x_t[5] = 21'b111111111111000101111;
        x_t[6] = 21'b111111111111110000011;
        x_t[7] = 21'b000000000100101100111;
        x_t[8] = 21'b000000000010010010000;
        x_t[9] = 21'b000000000000111001000;
        x_t[10] = 21'b000000000000000000101;
        x_t[11] = 21'b111111111110101101101;
        x_t[12] = 21'b111111111111000010111;
        x_t[13] = 21'b111111111111011001001;
        x_t[14] = 21'b000000000011000011101;
        x_t[15] = 21'b000000000010100000010;
        x_t[16] = 21'b000000000000111100111;
        x_t[17] = 21'b000000000000110000010;
        x_t[18] = 21'b111111111110110011111;
        x_t[19] = 21'b111111111111001110010;
        x_t[20] = 21'b000000000000000001110;
        x_t[21] = 21'b000000000000001010111;
        x_t[22] = 21'b000000000001010010100;
        x_t[23] = 21'b000000000001100100101;
        x_t[24] = 21'b000000000001011010010;
        x_t[25] = 21'b000000000001010111010;
        x_t[26] = 21'b111111111111100001111;
        x_t[27] = 21'b111111111111111001110;
        x_t[28] = 21'b000000000010000001100;
        x_t[29] = 21'b000000000001111001011;
        x_t[30] = 21'b000000000011110011110;
        x_t[31] = 21'b000000000000111101011;
        x_t[32] = 21'b000000000001000110110;
        x_t[33] = 21'b000000000000010100000;
        x_t[34] = 21'b111111111111101011100;
        x_t[35] = 21'b111111111111010110101;
        x_t[36] = 21'b000000000000010010100;
        x_t[37] = 21'b111111111010101010011;
        x_t[38] = 21'b000000000011100111010;
        x_t[39] = 21'b000000000000110001101;
        x_t[40] = 21'b000000000100111000110;
        x_t[41] = 21'b111111111110011001101;
        x_t[42] = 21'b000000000011001000000;
        x_t[43] = 21'b000000000010100001001;
        x_t[44] = 21'b000000000011011101110;
        x_t[45] = 21'b000000000001001100111;
        x_t[46] = 21'b000000000010000011100;
        x_t[47] = 21'b000000000010011100000;
        x_t[48] = 21'b000000000001110000011;
        x_t[49] = 21'b000000000001000101110;
        x_t[50] = 21'b000000000000001100110;
        x_t[51] = 21'b000000000000000111001;
        x_t[52] = 21'b000000000000001100101;
        x_t[53] = 21'b000000000000011111110;
        x_t[54] = 21'b000000000010001110111;
        x_t[55] = 21'b000000000001000110101;
        x_t[56] = 21'b000000000001111001100;
        x_t[57] = 21'b000000000000000010000;
        x_t[58] = 21'b000000000001001101111;
        x_t[59] = 21'b000000000010101100111;
        x_t[60] = 21'b111111111111011100101;
        x_t[61] = 21'b111111111111101010101;
        x_t[62] = 21'b000000000001000101101;
        x_t[63] = 21'b111111111110110101100;
        
        h_t_prev[0] = 21'b000000000010100111000;
        h_t_prev[1] = 21'b000000000011000001011;
        h_t_prev[2] = 21'b000000000000000001101;
        h_t_prev[3] = 21'b000000000000101001000;
        h_t_prev[4] = 21'b111111111111101010111;
        h_t_prev[5] = 21'b111111111111000101111;
        h_t_prev[6] = 21'b111111111111110000011;
        h_t_prev[7] = 21'b000000000100101100111;
        h_t_prev[8] = 21'b000000000010010010000;
        h_t_prev[9] = 21'b000000000000111001000;
        h_t_prev[10] = 21'b000000000000000000101;
        h_t_prev[11] = 21'b111111111110101101101;
        h_t_prev[12] = 21'b111111111111000010111;
        h_t_prev[13] = 21'b111111111111011001001;
        h_t_prev[14] = 21'b000000000011000011101;
        h_t_prev[15] = 21'b000000000010100000010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 18 timeout!");
                $fdisplay(fd_cycles, "Test Vector  18: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  18: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 18");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 19
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000100100111010;
        x_t[1] = 21'b000000000100001010111;
        x_t[2] = 21'b000000000001001111011;
        x_t[3] = 21'b000000000001011001011;
        x_t[4] = 21'b000000000000000100001;
        x_t[5] = 21'b111111111111100111010;
        x_t[6] = 21'b111111111111101010001;
        x_t[7] = 21'b000000000101010000100;
        x_t[8] = 21'b000000000010100001100;
        x_t[9] = 21'b000000000001100001000;
        x_t[10] = 21'b000000000000011101111;
        x_t[11] = 21'b000000000000000100010;
        x_t[12] = 21'b000000000000001111000;
        x_t[13] = 21'b111111111111011001001;
        x_t[14] = 21'b000000000011100011010;
        x_t[15] = 21'b000000000010101111100;
        x_t[16] = 21'b000000000001011010101;
        x_t[17] = 21'b000000000001101011100;
        x_t[18] = 21'b000000000000100111110;
        x_t[19] = 21'b000000000001010111101;
        x_t[20] = 21'b000000000001110010011;
        x_t[21] = 21'b000000000010100010111;
        x_t[22] = 21'b000000000011001000000;
        x_t[23] = 21'b000000000010110000000;
        x_t[24] = 21'b000000000100011101000;
        x_t[25] = 21'b000000000100010001110;
        x_t[26] = 21'b000000000001000011000;
        x_t[27] = 21'b000000000000101100111;
        x_t[28] = 21'b000000000010010100011;
        x_t[29] = 21'b000000000100111100111;
        x_t[30] = 21'b000000000110111010110;
        x_t[31] = 21'b000000000010100111111;
        x_t[32] = 21'b000000000011000001011;
        x_t[33] = 21'b000000000001110101001;
        x_t[34] = 21'b000000000001000110000;
        x_t[35] = 21'b000000000000101111011;
        x_t[36] = 21'b000000000000010111100;
        x_t[37] = 21'b111111111001110001011;
        x_t[38] = 21'b000000000111000101001;
        x_t[39] = 21'b111111111111101111100;
        x_t[40] = 21'b000000000110111011001;
        x_t[41] = 21'b111111111100000111101;
        x_t[42] = 21'b000000000101110011111;
        x_t[43] = 21'b000000000000000111100;
        x_t[44] = 21'b000000000101000111111;
        x_t[45] = 21'b000000000101001100010;
        x_t[46] = 21'b000000000011110000010;
        x_t[47] = 21'b000000000011111111100;
        x_t[48] = 21'b000000000011111111011;
        x_t[49] = 21'b000000000011010101011;
        x_t[50] = 21'b000000000011011101110;
        x_t[51] = 21'b000000000100011010100;
        x_t[52] = 21'b000000000100111111100;
        x_t[53] = 21'b000000000101000110111;
        x_t[54] = 21'b000000000101111110101;
        x_t[55] = 21'b000000000010110110111;
        x_t[56] = 21'b000000000011101001010;
        x_t[57] = 21'b000000000011011111110;
        x_t[58] = 21'b000000000101111111001;
        x_t[59] = 21'b000000000101110010010;
        x_t[60] = 21'b111111111111100000100;
        x_t[61] = 21'b000000000000011100011;
        x_t[62] = 21'b000000000001111101001;
        x_t[63] = 21'b111111111101000011000;
        
        h_t_prev[0] = 21'b000000000100100111010;
        h_t_prev[1] = 21'b000000000100001010111;
        h_t_prev[2] = 21'b000000000001001111011;
        h_t_prev[3] = 21'b000000000001011001011;
        h_t_prev[4] = 21'b000000000000000100001;
        h_t_prev[5] = 21'b111111111111100111010;
        h_t_prev[6] = 21'b111111111111101010001;
        h_t_prev[7] = 21'b000000000101010000100;
        h_t_prev[8] = 21'b000000000010100001100;
        h_t_prev[9] = 21'b000000000001100001000;
        h_t_prev[10] = 21'b000000000000011101111;
        h_t_prev[11] = 21'b000000000000000100010;
        h_t_prev[12] = 21'b000000000000001111000;
        h_t_prev[13] = 21'b111111111111011001001;
        h_t_prev[14] = 21'b000000000011100011010;
        h_t_prev[15] = 21'b000000000010101111100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 19 timeout!");
                $fdisplay(fd_cycles, "Test Vector  19: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  19: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 19");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 20
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000111001010000;
        x_t[1] = 21'b000000000110101100011;
        x_t[2] = 21'b000000000011110100011;
        x_t[3] = 21'b000000000011100000110;
        x_t[4] = 21'b000000000010111010000;
        x_t[5] = 21'b000000000010101110111;
        x_t[6] = 21'b000000000001111111100;
        x_t[7] = 21'b000000000111010100110;
        x_t[8] = 21'b000000000101010000111;
        x_t[9] = 21'b000000000100101001100;
        x_t[10] = 21'b000000000100001000110;
        x_t[11] = 21'b000000000011100100100;
        x_t[12] = 21'b000000000100110011101;
        x_t[13] = 21'b000000000011111110010;
        x_t[14] = 21'b000000000110000110110;
        x_t[15] = 21'b000000000101111011000;
        x_t[16] = 21'b000000000100101010111;
        x_t[17] = 21'b000000000100110101111;
        x_t[18] = 21'b000000000101001111000;
        x_t[19] = 21'b000000000110011011101;
        x_t[20] = 21'b000000000111001010100;
        x_t[21] = 21'b000000000011000100000;
        x_t[22] = 21'b000000000011001011001;
        x_t[23] = 21'b000000000010110010111;
        x_t[24] = 21'b000000000100010111000;
        x_t[25] = 21'b000000000100010100111;
        x_t[26] = 21'b000000000001111110001;
        x_t[27] = 21'b000000000001010100001;
        x_t[28] = 21'b000000000010100001000;
        x_t[29] = 21'b000000000011110110001;
        x_t[30] = 21'b000000000110111110101;
        x_t[31] = 21'b000000000011000110111;
        x_t[32] = 21'b000000000011010011100;
        x_t[33] = 21'b000000000010011110110;
        x_t[34] = 21'b000000000001111010011;
        x_t[35] = 21'b000000000001011011111;
        x_t[36] = 21'b000000000001011000001;
        x_t[37] = 21'b111111111010110010101;
        x_t[38] = 21'b000000000101101010011;
        x_t[39] = 21'b000000000010011000101;
        x_t[40] = 21'b000000000101100100010;
        x_t[41] = 21'b000000000001110001010;
        x_t[42] = 21'b000000000101000100100;
        x_t[43] = 21'b111111111111110001100;
        x_t[44] = 21'b000000000101011110010;
        x_t[45] = 21'b000000001000010101100;
        x_t[46] = 21'b000000000100101110011;
        x_t[47] = 21'b000000000100100010010;
        x_t[48] = 21'b000000000100011011111;
        x_t[49] = 21'b000000000100011010111;
        x_t[50] = 21'b000000000100101110100;
        x_t[51] = 21'b000000000110111110101;
        x_t[52] = 21'b000000000111101000011;
        x_t[53] = 21'b000000000111110011100;
        x_t[54] = 21'b000000001000000010011;
        x_t[55] = 21'b000000000011001000001;
        x_t[56] = 21'b000000000011100000101;
        x_t[57] = 21'b000000000100110101000;
        x_t[58] = 21'b000000001000100000101;
        x_t[59] = 21'b000000000111001101001;
        x_t[60] = 21'b000000000000100001101;
        x_t[61] = 21'b000000000010101001000;
        x_t[62] = 21'b000000000100000110000;
        x_t[63] = 21'b111111111110100011111;
        
        h_t_prev[0] = 21'b000000000111001010000;
        h_t_prev[1] = 21'b000000000110101100011;
        h_t_prev[2] = 21'b000000000011110100011;
        h_t_prev[3] = 21'b000000000011100000110;
        h_t_prev[4] = 21'b000000000010111010000;
        h_t_prev[5] = 21'b000000000010101110111;
        h_t_prev[6] = 21'b000000000001111111100;
        h_t_prev[7] = 21'b000000000111010100110;
        h_t_prev[8] = 21'b000000000101010000111;
        h_t_prev[9] = 21'b000000000100101001100;
        h_t_prev[10] = 21'b000000000100001000110;
        h_t_prev[11] = 21'b000000000011100100100;
        h_t_prev[12] = 21'b000000000100110011101;
        h_t_prev[13] = 21'b000000000011111110010;
        h_t_prev[14] = 21'b000000000110000110110;
        h_t_prev[15] = 21'b000000000101111011000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 20 timeout!");
                $fdisplay(fd_cycles, "Test Vector  20: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  20: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 20");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 21
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000010111010110;
        x_t[1] = 21'b000000000011001011010;
        x_t[2] = 21'b000000000001000000110;
        x_t[3] = 21'b000000000001000110000;
        x_t[4] = 21'b000000000001100100001;
        x_t[5] = 21'b000000000001111101000;
        x_t[6] = 21'b000000000010100100111;
        x_t[7] = 21'b000000000011001100001;
        x_t[8] = 21'b000000000010000010101;
        x_t[9] = 21'b000000000001110000001;
        x_t[10] = 21'b000000000001101100010;
        x_t[11] = 21'b000000000001111110100;
        x_t[12] = 21'b000000000100011100010;
        x_t[13] = 21'b000000000100101101111;
        x_t[14] = 21'b000000000011000011101;
        x_t[15] = 21'b000000000010111001110;
        x_t[16] = 21'b000000000010001100010;
        x_t[17] = 21'b000000000010111010100;
        x_t[18] = 21'b000000000011101010110;
        x_t[19] = 21'b000000000101010100010;
        x_t[20] = 21'b000000000110110001100;
        x_t[21] = 21'b111111111110111010110;
        x_t[22] = 21'b000000000000001001101;
        x_t[23] = 21'b000000000001011001000;
        x_t[24] = 21'b111111111111001110001;
        x_t[25] = 21'b111111111111001110100;
        x_t[26] = 21'b111111111111000100010;
        x_t[27] = 21'b000000000000001001100;
        x_t[28] = 21'b000000000001101011011;
        x_t[29] = 21'b111111111110101101101;
        x_t[30] = 21'b000000000001001000000;
        x_t[31] = 21'b000000000000111001000;
        x_t[32] = 21'b111111111111011001101;
        x_t[33] = 21'b111111111111010111111;
        x_t[34] = 21'b111111111111110000010;
        x_t[35] = 21'b111111111110111001000;
        x_t[36] = 21'b000000000001011000001;
        x_t[37] = 21'b111111111011011111011;
        x_t[38] = 21'b111111111111100110001;
        x_t[39] = 21'b000000000010111101011;
        x_t[40] = 21'b000000000010010101110;
        x_t[41] = 21'b000000000010110110110;
        x_t[42] = 21'b000000000000100010000;
        x_t[43] = 21'b000000000100111010110;
        x_t[44] = 21'b000000000010001001111;
        x_t[45] = 21'b000000000110001010001;
        x_t[46] = 21'b000000000010001101111;
        x_t[47] = 21'b000000000010001101000;
        x_t[48] = 21'b000000000010001000010;
        x_t[49] = 21'b000000000010011001001;
        x_t[50] = 21'b000000000011010100010;
        x_t[51] = 21'b000000000101100111110;
        x_t[52] = 21'b000000000110000010000;
        x_t[53] = 21'b000000000110000100001;
        x_t[54] = 21'b000000000101001110101;
        x_t[55] = 21'b000000000001110110001;
        x_t[56] = 21'b000000000010010111101;
        x_t[57] = 21'b000000000100001010011;
        x_t[58] = 21'b000000000111001001011;
        x_t[59] = 21'b000000000101110010010;
        x_t[60] = 21'b000000000000111000101;
        x_t[61] = 21'b000000000100001100011;
        x_t[62] = 21'b000000000101100110010;
        x_t[63] = 21'b000000000000011010101;
        
        h_t_prev[0] = 21'b000000000010111010110;
        h_t_prev[1] = 21'b000000000011001011010;
        h_t_prev[2] = 21'b000000000001000000110;
        h_t_prev[3] = 21'b000000000001000110000;
        h_t_prev[4] = 21'b000000000001100100001;
        h_t_prev[5] = 21'b000000000001111101000;
        h_t_prev[6] = 21'b000000000010100100111;
        h_t_prev[7] = 21'b000000000011001100001;
        h_t_prev[8] = 21'b000000000010000010101;
        h_t_prev[9] = 21'b000000000001110000001;
        h_t_prev[10] = 21'b000000000001101100010;
        h_t_prev[11] = 21'b000000000001111110100;
        h_t_prev[12] = 21'b000000000100011100010;
        h_t_prev[13] = 21'b000000000100101101111;
        h_t_prev[14] = 21'b000000000011000011101;
        h_t_prev[15] = 21'b000000000010111001110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 21 timeout!");
                $fdisplay(fd_cycles, "Test Vector  21: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  21: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 21");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 22
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000000110000101;
        x_t[1] = 21'b000000000001011010101;
        x_t[2] = 21'b111111111111101001011;
        x_t[3] = 21'b000000000000010000111;
        x_t[4] = 21'b000000000001000101110;
        x_t[5] = 21'b000000000001110001111;
        x_t[6] = 21'b000000000010100100111;
        x_t[7] = 21'b000000000010101101101;
        x_t[8] = 21'b000000000000111010011;
        x_t[9] = 21'b000000000001000011000;
        x_t[10] = 21'b000000000001011000101;
        x_t[11] = 21'b000000000010000011101;
        x_t[12] = 21'b000000000011111001001;
        x_t[13] = 21'b000000000100110100110;
        x_t[14] = 21'b000000000010110011111;
        x_t[15] = 21'b000000000010011011010;
        x_t[16] = 21'b000000000001110011011;
        x_t[17] = 21'b000000000010101011101;
        x_t[18] = 21'b000000000011001011001;
        x_t[19] = 21'b000000000100100010110;
        x_t[20] = 21'b000000000110001100000;
        x_t[21] = 21'b000000000000011000110;
        x_t[22] = 21'b000000000001001100010;
        x_t[23] = 21'b000000000001110000001;
        x_t[24] = 21'b000000000001100110011;
        x_t[25] = 21'b000000000001010111010;
        x_t[26] = 21'b111111111111101110100;
        x_t[27] = 21'b000000000000100001000;
        x_t[28] = 21'b000000000010000100101;
        x_t[29] = 21'b000000000001111101100;
        x_t[30] = 21'b000000000011111011100;
        x_t[31] = 21'b000000000001110010101;
        x_t[32] = 21'b000000000000100110111;
        x_t[33] = 21'b000000000000011101010;
        x_t[34] = 21'b000000000000011011001;
        x_t[35] = 21'b000000000000000011000;
        x_t[36] = 21'b000000000001101100000;
        x_t[37] = 21'b111111111010011110010;
        x_t[38] = 21'b000000000100000101100;
        x_t[39] = 21'b000000000010000010100;
        x_t[40] = 21'b000000000011011100011;
        x_t[41] = 21'b000000000001111111001;
        x_t[42] = 21'b000000000101111001111;
        x_t[43] = 21'b111111111111110001100;
        x_t[44] = 21'b000000000011101110100;
        x_t[45] = 21'b000000000100010110001;
        x_t[46] = 21'b000000000100011110111;
        x_t[47] = 21'b000000000100100010010;
        x_t[48] = 21'b000000000011110101110;
        x_t[49] = 21'b000000000011111010100;
        x_t[50] = 21'b000000000100010010000;
        x_t[51] = 21'b000000000101111011000;
        x_t[52] = 21'b000000000101111100111;
        x_t[53] = 21'b000000000101101000010;
        x_t[54] = 21'b000000000100110110101;
        x_t[55] = 21'b000000000100101011011;
        x_t[56] = 21'b000000000100110110100;
        x_t[57] = 21'b000000000101010111001;
        x_t[58] = 21'b000000000111001101110;
        x_t[59] = 21'b000000000101110010010;
        x_t[60] = 21'b000000000010000101011;
        x_t[61] = 21'b000000000101100011010;
        x_t[62] = 21'b000000000110010010101;
        x_t[63] = 21'b000000000011010011100;
        
        h_t_prev[0] = 21'b000000000000110000101;
        h_t_prev[1] = 21'b000000000001011010101;
        h_t_prev[2] = 21'b111111111111101001011;
        h_t_prev[3] = 21'b000000000000010000111;
        h_t_prev[4] = 21'b000000000001000101110;
        h_t_prev[5] = 21'b000000000001110001111;
        h_t_prev[6] = 21'b000000000010100100111;
        h_t_prev[7] = 21'b000000000010101101101;
        h_t_prev[8] = 21'b000000000000111010011;
        h_t_prev[9] = 21'b000000000001000011000;
        h_t_prev[10] = 21'b000000000001011000101;
        h_t_prev[11] = 21'b000000000010000011101;
        h_t_prev[12] = 21'b000000000011111001001;
        h_t_prev[13] = 21'b000000000100110100110;
        h_t_prev[14] = 21'b000000000010110011111;
        h_t_prev[15] = 21'b000000000010011011010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 22 timeout!");
                $fdisplay(fd_cycles, "Test Vector  22: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  22: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 22");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 23
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000100110001001;
        x_t[1] = 21'b000000000100001010111;
        x_t[2] = 21'b000000000001011001000;
        x_t[3] = 21'b000000000010000100111;
        x_t[4] = 21'b000000000001101001001;
        x_t[5] = 21'b000000000001110001111;
        x_t[6] = 21'b000000000010011110101;
        x_t[7] = 21'b000000000110101100001;
        x_t[8] = 21'b000000000011100100100;
        x_t[9] = 21'b000000000010101100010;
        x_t[10] = 21'b000000000010101011111;
        x_t[11] = 21'b000000000010011000000;
        x_t[12] = 21'b000000000011001010010;
        x_t[13] = 21'b000000000011100010111;
        x_t[14] = 21'b000000000110000110110;
        x_t[15] = 21'b000000000100011111011;
        x_t[16] = 21'b000000000011100000100;
        x_t[17] = 21'b000000000011101011111;
        x_t[18] = 21'b000000000011010101110;
        x_t[19] = 21'b000000000100010010010;
        x_t[20] = 21'b000000000101000111001;
        x_t[21] = 21'b000000000001110011111;
        x_t[22] = 21'b000000000010101011011;
        x_t[23] = 21'b000000000010111011101;
        x_t[24] = 21'b000000000010111011101;
        x_t[25] = 21'b000000000010110111101;
        x_t[26] = 21'b000000000000010100100;
        x_t[27] = 21'b000000000001001100010;
        x_t[28] = 21'b000000000011101100100;
        x_t[29] = 21'b000000000011010000110;
        x_t[30] = 21'b000000000100111010000;
        x_t[31] = 21'b000000000001011100100;
        x_t[32] = 21'b000000000001001011010;
        x_t[33] = 21'b000000000000101111110;
        x_t[34] = 21'b000000000000011011001;
        x_t[35] = 21'b111111111111111001001;
        x_t[36] = 21'b000000000001100010000;
        x_t[37] = 21'b111111111011111100000;
        x_t[38] = 21'b000000000100001010101;
        x_t[39] = 21'b000000000010010001010;
        x_t[40] = 21'b000000000100111000110;
        x_t[41] = 21'b000000000000110010101;
        x_t[42] = 21'b000000000101101110000;
        x_t[43] = 21'b000000000001011111010;
        x_t[44] = 21'b000000000110110010000;
        x_t[45] = 21'b000000000011010000100;
        x_t[46] = 21'b000000000110100000011;
        x_t[47] = 21'b000000000101011001000;
        x_t[48] = 21'b000000000100001101101;
        x_t[49] = 21'b000000000011111010100;
        x_t[50] = 21'b000000000011110101100;
        x_t[51] = 21'b000000000101000101111;
        x_t[52] = 21'b000000000100111010011;
        x_t[53] = 21'b000000000100101011000;
        x_t[54] = 21'b000000000100100100110;
        x_t[55] = 21'b000000000100111000011;
        x_t[56] = 21'b000000000100101001101;
        x_t[57] = 21'b000000000100101000010;
        x_t[58] = 21'b000000000110100010001;
        x_t[59] = 21'b000000000101100010100;
        x_t[60] = 21'b000000000011010101111;
        x_t[61] = 21'b000000000110011001001;
        x_t[62] = 21'b000000000110001110111;
        x_t[63] = 21'b000000000101001110110;
        
        h_t_prev[0] = 21'b000000000100110001001;
        h_t_prev[1] = 21'b000000000100001010111;
        h_t_prev[2] = 21'b000000000001011001000;
        h_t_prev[3] = 21'b000000000010000100111;
        h_t_prev[4] = 21'b000000000001101001001;
        h_t_prev[5] = 21'b000000000001110001111;
        h_t_prev[6] = 21'b000000000010011110101;
        h_t_prev[7] = 21'b000000000110101100001;
        h_t_prev[8] = 21'b000000000011100100100;
        h_t_prev[9] = 21'b000000000010101100010;
        h_t_prev[10] = 21'b000000000010101011111;
        h_t_prev[11] = 21'b000000000010011000000;
        h_t_prev[12] = 21'b000000000011001010010;
        h_t_prev[13] = 21'b000000000011100010111;
        h_t_prev[14] = 21'b000000000110000110110;
        h_t_prev[15] = 21'b000000000100011111011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 23 timeout!");
                $fdisplay(fd_cycles, "Test Vector  23: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  23: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 23");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 24
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000001000100011;
        x_t[1] = 21'b000000000001101110010;
        x_t[2] = 21'b111111111111110111111;
        x_t[3] = 21'b000000000000110111100;
        x_t[4] = 21'b111111111111111010000;
        x_t[5] = 21'b111111111111100001101;
        x_t[6] = 21'b000000000000011011111;
        x_t[7] = 21'b000000000011001100001;
        x_t[8] = 21'b000000000001011001010;
        x_t[9] = 21'b000000000001011100000;
        x_t[10] = 21'b000000000001100010011;
        x_t[11] = 21'b000000000000001001011;
        x_t[12] = 21'b000000000000111101110;
        x_t[13] = 21'b000000000000010110100;
        x_t[14] = 21'b000000000100011101010;
        x_t[15] = 21'b000000000011000011111;
        x_t[16] = 21'b000000000010010001001;
        x_t[17] = 21'b000000000010101011101;
        x_t[18] = 21'b000000000001110110111;
        x_t[19] = 21'b000000000010100100100;
        x_t[20] = 21'b000000000011000011110;
        x_t[21] = 21'b111111111110101010010;
        x_t[22] = 21'b111111111111110011011;
        x_t[23] = 21'b000000000000100111101;
        x_t[24] = 21'b111111111111010001001;
        x_t[25] = 21'b111111111111010001101;
        x_t[26] = 21'b111111111101110100000;
        x_t[27] = 21'b111111111110101011001;
        x_t[28] = 21'b000000000001001111001;
        x_t[29] = 21'b111111111111000010011;
        x_t[30] = 21'b000000000001100111010;
        x_t[31] = 21'b111111111111100000010;
        x_t[32] = 21'b111111111111001100000;
        x_t[33] = 21'b111111111110101110010;
        x_t[34] = 21'b111111111110001100010;
        x_t[35] = 21'b111111111101011011010;
        x_t[36] = 21'b111111111110100000001;
        x_t[37] = 21'b111111111010100110011;
        x_t[38] = 21'b111111111111111010010;
        x_t[39] = 21'b111111111111011001100;
        x_t[40] = 21'b000000000101001110100;
        x_t[41] = 21'b111111111011100100110;
        x_t[42] = 21'b000000000101001010011;
        x_t[43] = 21'b000000000010001011001;
        x_t[44] = 21'b000000000110101100011;
        x_t[45] = 21'b000000000100011101111;
        x_t[46] = 21'b000000000110001011101;
        x_t[47] = 21'b000000000100110110001;
        x_t[48] = 21'b000000000100000100001;
        x_t[49] = 21'b000000000011101100101;
        x_t[50] = 21'b000000000011100010100;
        x_t[51] = 21'b000000000100111100010;
        x_t[52] = 21'b000000000100111010011;
        x_t[53] = 21'b000000000100110000101;
        x_t[54] = 21'b000000000101100110101;
        x_t[55] = 21'b000000000011111011111;
        x_t[56] = 21'b000000000100001011101;
        x_t[57] = 21'b000000000100010111001;
        x_t[58] = 21'b000000000110101111001;
        x_t[59] = 21'b000000000110011001110;
        x_t[60] = 21'b000000000011011001101;
        x_t[61] = 21'b000000000110011001001;
        x_t[62] = 21'b000000000110000000001;
        x_t[63] = 21'b000000000101001010011;
        
        h_t_prev[0] = 21'b000000000001000100011;
        h_t_prev[1] = 21'b000000000001101110010;
        h_t_prev[2] = 21'b111111111111110111111;
        h_t_prev[3] = 21'b000000000000110111100;
        h_t_prev[4] = 21'b111111111111111010000;
        h_t_prev[5] = 21'b111111111111100001101;
        h_t_prev[6] = 21'b000000000000011011111;
        h_t_prev[7] = 21'b000000000011001100001;
        h_t_prev[8] = 21'b000000000001011001010;
        h_t_prev[9] = 21'b000000000001011100000;
        h_t_prev[10] = 21'b000000000001100010011;
        h_t_prev[11] = 21'b000000000000001001011;
        h_t_prev[12] = 21'b000000000000111101110;
        h_t_prev[13] = 21'b000000000000010110100;
        h_t_prev[14] = 21'b000000000100011101010;
        h_t_prev[15] = 21'b000000000011000011111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 24 timeout!");
                $fdisplay(fd_cycles, "Test Vector  24: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  24: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 24");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 25
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000001001001010;
        x_t[1] = 21'b000000000010010000100;
        x_t[2] = 21'b000000000000011110110;
        x_t[3] = 21'b000000000001001111110;
        x_t[4] = 21'b111111111111111111000;
        x_t[5] = 21'b111111111111000101111;
        x_t[6] = 21'b111111111110101011111;
        x_t[7] = 21'b000000000101010000100;
        x_t[8] = 21'b000000000010110001000;
        x_t[9] = 21'b000000000010101100010;
        x_t[10] = 21'b000000000010100010000;
        x_t[11] = 21'b000000000001010000101;
        x_t[12] = 21'b000000000001011011000;
        x_t[13] = 21'b111111111111110100011;
        x_t[14] = 21'b000000000110000110110;
        x_t[15] = 21'b000000000100111000111;
        x_t[16] = 21'b000000000011100000100;
        x_t[17] = 21'b000000000011110101101;
        x_t[18] = 21'b000000000010110000111;
        x_t[19] = 21'b000000000011001010111;
        x_t[20] = 21'b000000000011101001010;
        x_t[21] = 21'b111111111111101111010;
        x_t[22] = 21'b000000000000001001101;
        x_t[23] = 21'b000000000000100111101;
        x_t[24] = 21'b000000000000110101101;
        x_t[25] = 21'b000000000000101000101;
        x_t[26] = 21'b111111111110111011111;
        x_t[27] = 21'b111111111110101111001;
        x_t[28] = 21'b000000000000011111111;
        x_t[29] = 21'b000000000000000000110;
        x_t[30] = 21'b000000000010111101001;
        x_t[31] = 21'b000000000000011110011;
        x_t[32] = 21'b000000000001000010001;
        x_t[33] = 21'b000000000000100001111;
        x_t[34] = 21'b111111111111011000100;
        x_t[35] = 21'b111111111110110100001;
        x_t[36] = 21'b111111111110110100000;
        x_t[37] = 21'b111111111010100010010;
        x_t[38] = 21'b000000000001011010001;
        x_t[39] = 21'b111111111110110100110;
        x_t[40] = 21'b000000000010011011001;
        x_t[41] = 21'b111111111100100011011;
        x_t[42] = 21'b000000000011110001100;
        x_t[43] = 21'b000000000010100001001;
        x_t[44] = 21'b000000000100010101101;
        x_t[45] = 21'b000000000101000100100;
        x_t[46] = 21'b000000000101010111111;
        x_t[47] = 21'b000000000101011001000;
        x_t[48] = 21'b000000000100111000100;
        x_t[49] = 21'b000000000100100100001;
        x_t[50] = 21'b000000000100100000010;
        x_t[51] = 21'b000000000101001111101;
        x_t[52] = 21'b000000000101000100101;
        x_t[53] = 21'b000000000100110110001;
        x_t[54] = 21'b000000000101001110101;
        x_t[55] = 21'b000000000100011010001;
        x_t[56] = 21'b000000000100011000100;
        x_t[57] = 21'b000000000100010111001;
        x_t[58] = 21'b000000000110100010001;
        x_t[59] = 21'b000000000101110010010;
        x_t[60] = 21'b000000000011000110100;
        x_t[61] = 21'b000000000101111100001;
        x_t[62] = 21'b000000000101100010100;
        x_t[63] = 21'b000000000100010101100;
        
        h_t_prev[0] = 21'b000000000001001001010;
        h_t_prev[1] = 21'b000000000010010000100;
        h_t_prev[2] = 21'b000000000000011110110;
        h_t_prev[3] = 21'b000000000001001111110;
        h_t_prev[4] = 21'b111111111111111111000;
        h_t_prev[5] = 21'b111111111111000101111;
        h_t_prev[6] = 21'b111111111110101011111;
        h_t_prev[7] = 21'b000000000101010000100;
        h_t_prev[8] = 21'b000000000010110001000;
        h_t_prev[9] = 21'b000000000010101100010;
        h_t_prev[10] = 21'b000000000010100010000;
        h_t_prev[11] = 21'b000000000001010000101;
        h_t_prev[12] = 21'b000000000001011011000;
        h_t_prev[13] = 21'b111111111111110100011;
        h_t_prev[14] = 21'b000000000110000110110;
        h_t_prev[15] = 21'b000000000100111000111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 25 timeout!");
                $fdisplay(fd_cycles, "Test Vector  25: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  25: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 25");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 26
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000001010011001;
        x_t[1] = 21'b000000000011000110011;
        x_t[2] = 21'b000000000001110001011;
        x_t[3] = 21'b000000000010110000011;
        x_t[4] = 21'b000000000001001111111;
        x_t[5] = 21'b000000000000101111011;
        x_t[6] = 21'b000000000000010101101;
        x_t[7] = 21'b000000000100000100001;
        x_t[8] = 21'b000000000010110110001;
        x_t[9] = 21'b000000000010110110010;
        x_t[10] = 21'b000000000010101011111;
        x_t[11] = 21'b000000000001111001100;
        x_t[12] = 21'b000000000010001001111;
        x_t[13] = 21'b000000000000110001110;
        x_t[14] = 21'b000000000100000010111;
        x_t[15] = 21'b000000000011011000010;
        x_t[16] = 21'b000000000010110011111;
        x_t[17] = 21'b000000000011011101000;
        x_t[18] = 21'b000000000010100001000;
        x_t[19] = 21'b000000000010101111100;
        x_t[20] = 21'b000000000011010000010;
        x_t[21] = 21'b111111111111000011000;
        x_t[22] = 21'b111111111111110110100;
        x_t[23] = 21'b000000000000011111000;
        x_t[24] = 21'b111111111111100000011;
        x_t[25] = 21'b111111111111100111011;
        x_t[26] = 21'b111111111111100001111;
        x_t[27] = 21'b111111111111010010100;
        x_t[28] = 21'b000000000000101111101;
        x_t[29] = 21'b111111111101011010011;
        x_t[30] = 21'b000000000001011111011;
        x_t[31] = 21'b000000000000010101100;
        x_t[32] = 21'b000000000000110000000;
        x_t[33] = 21'b000000000000100001111;
        x_t[34] = 21'b111111111111101011100;
        x_t[35] = 21'b111111111110100101010;
        x_t[36] = 21'b111111111111011011111;
        x_t[37] = 21'b111111111010110110101;
        x_t[38] = 21'b111111111110100100100;
        x_t[39] = 21'b000000000000000101101;
        x_t[40] = 21'b000000000000001000011;
        x_t[41] = 21'b111111111110101110100;
        x_t[42] = 21'b000000000001011101010;
        x_t[43] = 21'b111111111101111000111;
        x_t[44] = 21'b000000000010001111100;
        x_t[45] = 21'b000000000010101001110;
        x_t[46] = 21'b000000000010010011000;
        x_t[47] = 21'b000000000010010010000;
        x_t[48] = 21'b000000000010100100110;
        x_t[49] = 21'b000000000010000110101;
        x_t[50] = 21'b000000000010100100110;
        x_t[51] = 21'b000000000011010010000;
        x_t[52] = 21'b000000000011001001111;
        x_t[53] = 21'b000000000010110110001;
        x_t[54] = 21'b000000000011001010110;
        x_t[55] = 21'b000000000010000011001;
        x_t[56] = 21'b000000000010010011010;
        x_t[57] = 21'b000000000010010011000;
        x_t[58] = 21'b000000000100011111010;
        x_t[59] = 21'b000000000011110111111;
        x_t[60] = 21'b000000000001111001111;
        x_t[61] = 21'b000000000100010100101;
        x_t[62] = 21'b000000000011100100110;
        x_t[63] = 21'b000000000001111111111;
        
        h_t_prev[0] = 21'b000000000001010011001;
        h_t_prev[1] = 21'b000000000011000110011;
        h_t_prev[2] = 21'b000000000001110001011;
        h_t_prev[3] = 21'b000000000010110000011;
        h_t_prev[4] = 21'b000000000001001111111;
        h_t_prev[5] = 21'b000000000000101111011;
        h_t_prev[6] = 21'b000000000000010101101;
        h_t_prev[7] = 21'b000000000100000100001;
        h_t_prev[8] = 21'b000000000010110110001;
        h_t_prev[9] = 21'b000000000010110110010;
        h_t_prev[10] = 21'b000000000010101011111;
        h_t_prev[11] = 21'b000000000001111001100;
        h_t_prev[12] = 21'b000000000010001001111;
        h_t_prev[13] = 21'b000000000000110001110;
        h_t_prev[14] = 21'b000000000100000010111;
        h_t_prev[15] = 21'b000000000011011000010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 26 timeout!");
                $fdisplay(fd_cycles, "Test Vector  26: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  26: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 26");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 27
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111111001110000;
        x_t[1] = 21'b000000000000101110101;
        x_t[2] = 21'b000000000000000110100;
        x_t[3] = 21'b000000000001001010111;
        x_t[4] = 21'b111111111111111111000;
        x_t[5] = 21'b111111111111110010010;
        x_t[6] = 21'b000000000000001001010;
        x_t[7] = 21'b000000000000100100001;
        x_t[8] = 21'b111111111111110111011;
        x_t[9] = 21'b000000000000111110000;
        x_t[10] = 21'b000000000001000101001;
        x_t[11] = 21'b000000000000000100010;
        x_t[12] = 21'b000000000000101100010;
        x_t[13] = 21'b000000000000010110100;
        x_t[14] = 21'b000000000000101010110;
        x_t[15] = 21'b000000000001001001111;
        x_t[16] = 21'b000000000000111100111;
        x_t[17] = 21'b000000000001110101011;
        x_t[18] = 21'b000000000000110010011;
        x_t[19] = 21'b000000000001000111001;
        x_t[20] = 21'b000000000010011000000;
        x_t[21] = 21'b111111111111101100100;
        x_t[22] = 21'b000000000000100011000;
        x_t[23] = 21'b000000000001010011001;
        x_t[24] = 21'b000000000000001011000;
        x_t[25] = 21'b000000000000001001101;
        x_t[26] = 21'b111111111111011001011;
        x_t[27] = 21'b111111111111100110001;
        x_t[28] = 21'b000000000001100010000;
        x_t[29] = 21'b111111111111010111001;
        x_t[30] = 21'b000000000001100011010;
        x_t[31] = 21'b000000000000001100101;
        x_t[32] = 21'b000000000000000010100;
        x_t[33] = 21'b111111111111111100111;
        x_t[34] = 21'b111111111111000101011;
        x_t[35] = 21'b111111111110010001100;
        x_t[36] = 21'b111111111111110100101;
        x_t[37] = 21'b111111111011111100000;
        x_t[38] = 21'b000000000000100010101;
        x_t[39] = 21'b000000000000111001000;
        x_t[40] = 21'b000000000010101011100;
        x_t[41] = 21'b111111111101110110111;
        x_t[42] = 21'b000000000010001100101;
        x_t[43] = 21'b111111111110100100110;
        x_t[44] = 21'b000000000010001001111;
        x_t[45] = 21'b000000000100011101111;
        x_t[46] = 21'b000000000001111110010;
        x_t[47] = 21'b000000000001111110001;
        x_t[48] = 21'b000000000010101001101;
        x_t[49] = 21'b000000000010000010000;
        x_t[50] = 21'b000000000001110101010;
        x_t[51] = 21'b000000000010011000000;
        x_t[52] = 21'b000000000010001100100;
        x_t[53] = 21'b000000000010001111001;
        x_t[54] = 21'b000000000011101110110;
        x_t[55] = 21'b000000000010001011110;
        x_t[56] = 21'b000000000010110101101;
        x_t[57] = 21'b000000000010000110010;
        x_t[58] = 21'b000000000011100110100;
        x_t[59] = 21'b000000000011100000010;
        x_t[60] = 21'b000000000001001011111;
        x_t[61] = 21'b000000000011010010011;
        x_t[62] = 21'b000000000010001100000;
        x_t[63] = 21'b000000000001000010010;
        
        h_t_prev[0] = 21'b111111111111001110000;
        h_t_prev[1] = 21'b000000000000101110101;
        h_t_prev[2] = 21'b000000000000000110100;
        h_t_prev[3] = 21'b000000000001001010111;
        h_t_prev[4] = 21'b111111111111111111000;
        h_t_prev[5] = 21'b111111111111110010010;
        h_t_prev[6] = 21'b000000000000001001010;
        h_t_prev[7] = 21'b000000000000100100001;
        h_t_prev[8] = 21'b111111111111110111011;
        h_t_prev[9] = 21'b000000000000111110000;
        h_t_prev[10] = 21'b000000000001000101001;
        h_t_prev[11] = 21'b000000000000000100010;
        h_t_prev[12] = 21'b000000000000101100010;
        h_t_prev[13] = 21'b000000000000010110100;
        h_t_prev[14] = 21'b000000000000101010110;
        h_t_prev[15] = 21'b000000000001001001111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 27 timeout!");
                $fdisplay(fd_cycles, "Test Vector  27: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  27: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 27");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 28
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000001000100011;
        x_t[1] = 21'b000000000001000111001;
        x_t[2] = 21'b111111111111110011001;
        x_t[3] = 21'b000000000000000111010;
        x_t[4] = 21'b111111111110111101011;
        x_t[5] = 21'b111111111110110101010;
        x_t[6] = 21'b111111111111100011111;
        x_t[7] = 21'b000000000011000010000;
        x_t[8] = 21'b000000000000110000000;
        x_t[9] = 21'b000000000001001000000;
        x_t[10] = 21'b000000000001000101001;
        x_t[11] = 21'b111111111111010110011;
        x_t[12] = 21'b111111111111100110000;
        x_t[13] = 21'b111111111111000100110;
        x_t[14] = 21'b000000000010010100001;
        x_t[15] = 21'b000000000010000110111;
        x_t[16] = 21'b000000000001011111101;
        x_t[17] = 21'b000000000001111010010;
        x_t[18] = 21'b111111111111111101101;
        x_t[19] = 21'b111111111111110100110;
        x_t[20] = 21'b000000000001001100111;
        x_t[21] = 21'b000000000000100110100;
        x_t[22] = 21'b000000000001010010100;
        x_t[23] = 21'b000000000001101101010;
        x_t[24] = 21'b000000000001010100001;
        x_t[25] = 21'b000000000001010100001;
        x_t[26] = 21'b111111111110111011111;
        x_t[27] = 21'b111111111111001110100;
        x_t[28] = 21'b000000000000111100010;
        x_t[29] = 21'b000000000000010001011;
        x_t[30] = 21'b000000000010101001100;
        x_t[31] = 21'b111111111111010011000;
        x_t[32] = 21'b111111111111001100000;
        x_t[33] = 21'b111111111111000101011;
        x_t[34] = 21'b111111111110001100010;
        x_t[35] = 21'b111111111101100000001;
        x_t[36] = 21'b111111111110101111001;
        x_t[37] = 21'b111111111011100011100;
        x_t[38] = 21'b000000000001111101011;
        x_t[39] = 21'b111111111110101101011;
        x_t[40] = 21'b000000000011010001100;
        x_t[41] = 21'b111111111100011100100;
        x_t[42] = 21'b000000000001110101000;
        x_t[43] = 21'b000000000011000010000;
        x_t[44] = 21'b000000000010110001000;
        x_t[45] = 21'b000000000010000011001;
        x_t[46] = 21'b000000000010101100111;
        x_t[47] = 21'b000000000010100001000;
        x_t[48] = 21'b000000000010100100110;
        x_t[49] = 21'b000000000001110100001;
        x_t[50] = 21'b000000000000100100100;
        x_t[51] = 21'b000000000000010101101;
        x_t[52] = 21'b111111111111101101111;
        x_t[53] = 21'b111111111111101000001;
        x_t[54] = 21'b000000000001001101000;
        x_t[55] = 21'b000000000010110010100;
        x_t[56] = 21'b000000000011001011001;
        x_t[57] = 21'b000000000001000110010;
        x_t[58] = 21'b000000000001000101001;
        x_t[59] = 21'b000000000001000010011;
        x_t[60] = 21'b000000000001010011100;
        x_t[61] = 21'b000000000010110001011;
        x_t[62] = 21'b000000000001001101001;
        x_t[63] = 21'b000000000001001011001;
        
        h_t_prev[0] = 21'b000000000001000100011;
        h_t_prev[1] = 21'b000000000001000111001;
        h_t_prev[2] = 21'b111111111111110011001;
        h_t_prev[3] = 21'b000000000000000111010;
        h_t_prev[4] = 21'b111111111110111101011;
        h_t_prev[5] = 21'b111111111110110101010;
        h_t_prev[6] = 21'b111111111111100011111;
        h_t_prev[7] = 21'b000000000011000010000;
        h_t_prev[8] = 21'b000000000000110000000;
        h_t_prev[9] = 21'b000000000001001000000;
        h_t_prev[10] = 21'b000000000001000101001;
        h_t_prev[11] = 21'b111111111111010110011;
        h_t_prev[12] = 21'b111111111111100110000;
        h_t_prev[13] = 21'b111111111111000100110;
        h_t_prev[14] = 21'b000000000010010100001;
        h_t_prev[15] = 21'b000000000010000110111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 28 timeout!");
                $fdisplay(fd_cycles, "Test Vector  28: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  28: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 28");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 29
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000001010011001;
        x_t[1] = 21'b000000000001010000111;
        x_t[2] = 21'b111111111111011010110;
        x_t[3] = 21'b111111111111100101011;
        x_t[4] = 21'b111111111110000000110;
        x_t[5] = 21'b111111111101000110011;
        x_t[6] = 21'b111111111110000000011;
        x_t[7] = 21'b000000000011011011011;
        x_t[8] = 21'b000000000001101000110;
        x_t[9] = 21'b000000000001000011000;
        x_t[10] = 21'b000000000000011001000;
        x_t[11] = 21'b111111111111001100010;
        x_t[12] = 21'b111111111110000010100;
        x_t[13] = 21'b111111111101010000111;
        x_t[14] = 21'b000000000010110011111;
        x_t[15] = 21'b000000000010000001110;
        x_t[16] = 21'b000000000001010101110;
        x_t[17] = 21'b000000000001010010111;
        x_t[18] = 21'b111111111110111001001;
        x_t[19] = 21'b111111111110010001111;
        x_t[20] = 21'b111111111111001001100;
        x_t[21] = 21'b000000000000001010111;
        x_t[22] = 21'b000000000000110110000;
        x_t[23] = 21'b000000000001000100101;
        x_t[24] = 21'b000000000001000100111;
        x_t[25] = 21'b000000000001000100101;
        x_t[26] = 21'b111111111111010001000;
        x_t[27] = 21'b111111111110111110110;
        x_t[28] = 21'b000000000000010110011;
        x_t[29] = 21'b000000000000110110111;
        x_t[30] = 21'b000000000010010110000;
        x_t[31] = 21'b111111111111110110100;
        x_t[32] = 21'b111111111111110100111;
        x_t[33] = 21'b000000000000000001100;
        x_t[34] = 21'b111111111110111011111;
        x_t[35] = 21'b111111111101111000111;
        x_t[36] = 21'b111111111110111110000;
        x_t[37] = 21'b111111111011011111011;
        x_t[38] = 21'b000000000010010110101;
        x_t[39] = 21'b111111111110110100110;
        x_t[40] = 21'b000000000011100111010;
        x_t[41] = 21'b000000000000100100110;
        x_t[42] = 21'b000000000101011100010;
        x_t[43] = 21'b111111111111010000101;
        x_t[44] = 21'b000000000100100110011;
        x_t[45] = 21'b000000000000011110100;
        x_t[46] = 21'b000000000100001111011;
        x_t[47] = 21'b000000000011010111101;
        x_t[48] = 21'b000000000011001111110;
        x_t[49] = 21'b000000000010010100100;
        x_t[50] = 21'b000000000001001111010;
        x_t[51] = 21'b000000000000000010011;
        x_t[52] = 21'b111111111111100011101;
        x_t[53] = 21'b111111111110111011101;
        x_t[54] = 21'b000000000000000101000;
        x_t[55] = 21'b000000000100000100100;
        x_t[56] = 21'b000000000100001011101;
        x_t[57] = 21'b000000000001001110110;
        x_t[58] = 21'b111111111111101101111;
        x_t[59] = 21'b111111111111111111010;
        x_t[60] = 21'b000000000010001101000;
        x_t[61] = 21'b000000000010101101010;
        x_t[62] = 21'b000000000000001010100;
        x_t[63] = 21'b000000000001011100101;
        
        h_t_prev[0] = 21'b000000000001010011001;
        h_t_prev[1] = 21'b000000000001010000111;
        h_t_prev[2] = 21'b111111111111011010110;
        h_t_prev[3] = 21'b111111111111100101011;
        h_t_prev[4] = 21'b111111111110000000110;
        h_t_prev[5] = 21'b111111111101000110011;
        h_t_prev[6] = 21'b111111111110000000011;
        h_t_prev[7] = 21'b000000000011011011011;
        h_t_prev[8] = 21'b000000000001101000110;
        h_t_prev[9] = 21'b000000000001000011000;
        h_t_prev[10] = 21'b000000000000011001000;
        h_t_prev[11] = 21'b111111111111001100010;
        h_t_prev[12] = 21'b111111111110000010100;
        h_t_prev[13] = 21'b111111111101010000111;
        h_t_prev[14] = 21'b000000000010110011111;
        h_t_prev[15] = 21'b000000000010000001110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 29 timeout!");
                $fdisplay(fd_cycles, "Test Vector  29: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  29: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 29");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 30
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000010111111101;
        x_t[1] = 21'b000000000011100011101;
        x_t[2] = 21'b000000000001100111101;
        x_t[3] = 21'b000000000001111011010;
        x_t[4] = 21'b000000000000110110101;
        x_t[5] = 21'b111111111111100111010;
        x_t[6] = 21'b000000000000101110101;
        x_t[7] = 21'b000000000101100100111;
        x_t[8] = 21'b000000000011101001110;
        x_t[9] = 21'b000000000011001010010;
        x_t[10] = 21'b000000000010101011111;
        x_t[11] = 21'b000000000001001011101;
        x_t[12] = 21'b000000000000000011010;
        x_t[13] = 21'b000000000000111000101;
        x_t[14] = 21'b000000000100001000010;
        x_t[15] = 21'b000000000011100010011;
        x_t[16] = 21'b000000000010101110111;
        x_t[17] = 21'b000000000010110101100;
        x_t[18] = 21'b000000000000011101010;
        x_t[19] = 21'b111111111111010011110;
        x_t[20] = 21'b000000000000001110010;
        x_t[21] = 21'b000000000010011010100;
        x_t[22] = 21'b000000000011001000000;
        x_t[23] = 21'b000000000010111110100;
        x_t[24] = 21'b000000000011100011010;
        x_t[25] = 21'b000000000011011100111;
        x_t[26] = 21'b000000000001101101010;
        x_t[27] = 21'b000000000001010100001;
        x_t[28] = 21'b000000000010011101111;
        x_t[29] = 21'b000000000011110010000;
        x_t[30] = 21'b000000000100010110111;
        x_t[31] = 21'b000000000010001000111;
        x_t[32] = 21'b000000000010010011111;
        x_t[33] = 21'b000000000010011110110;
        x_t[34] = 21'b000000000001100010101;
        x_t[35] = 21'b000000000000011011110;
        x_t[36] = 21'b000000000001010011001;
        x_t[37] = 21'b111111111101011001110;
        x_t[38] = 21'b000000000100100011110;
        x_t[39] = 21'b000000000010001001111;
        x_t[40] = 21'b000000000100101000100;
        x_t[41] = 21'b000000000010000110001;
        x_t[42] = 21'b000000000111101010100;
        x_t[43] = 21'b111111111110100100110;
        x_t[44] = 21'b000000000101111010001;
        x_t[45] = 21'b111111111111011000111;
        x_t[46] = 21'b000000000101100010010;
        x_t[47] = 21'b000000000011110101100;
        x_t[48] = 21'b000000000011010100100;
        x_t[49] = 21'b000000000010001111111;
        x_t[50] = 21'b000000000000011111110;
        x_t[51] = 21'b111111111101110001011;
        x_t[52] = 21'b111111111101001111010;
        x_t[53] = 21'b111111111100001001100;
        x_t[54] = 21'b111111111101100011010;
        x_t[55] = 21'b000000000100011110100;
        x_t[56] = 21'b000000000100000011000;
        x_t[57] = 21'b111111111111011011101;
        x_t[58] = 21'b111111111011011011001;
        x_t[59] = 21'b111111111100110010000;
        x_t[60] = 21'b000000000011000010101;
        x_t[61] = 21'b000000000010001100001;
        x_t[62] = 21'b111111111110000001101;
        x_t[63] = 21'b000000000001101001111;
        
        h_t_prev[0] = 21'b000000000010111111101;
        h_t_prev[1] = 21'b000000000011100011101;
        h_t_prev[2] = 21'b000000000001100111101;
        h_t_prev[3] = 21'b000000000001111011010;
        h_t_prev[4] = 21'b000000000000110110101;
        h_t_prev[5] = 21'b111111111111100111010;
        h_t_prev[6] = 21'b000000000000101110101;
        h_t_prev[7] = 21'b000000000101100100111;
        h_t_prev[8] = 21'b000000000011101001110;
        h_t_prev[9] = 21'b000000000011001010010;
        h_t_prev[10] = 21'b000000000010101011111;
        h_t_prev[11] = 21'b000000000001001011101;
        h_t_prev[12] = 21'b000000000000000011010;
        h_t_prev[13] = 21'b000000000000111000101;
        h_t_prev[14] = 21'b000000000100001000010;
        h_t_prev[15] = 21'b000000000011100010011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 30 timeout!");
                $fdisplay(fd_cycles, "Test Vector  30: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  30: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 30");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 31
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000011111010111;
        x_t[1] = 21'b000000000100000001000;
        x_t[2] = 21'b000000000001110001011;
        x_t[3] = 21'b000000000010110101010;
        x_t[4] = 21'b000000000001010100111;
        x_t[5] = 21'b111111111111111101011;
        x_t[6] = 21'b000000000000000011000;
        x_t[7] = 21'b000000000101000110010;
        x_t[8] = 21'b000000000011000101101;
        x_t[9] = 21'b000000000010101100010;
        x_t[10] = 21'b000000000010001110100;
        x_t[11] = 21'b111111111111110101000;
        x_t[12] = 21'b111111111110110111001;
        x_t[13] = 21'b111111111110001110010;
        x_t[14] = 21'b000000000011101101111;
        x_t[15] = 21'b000000000010011011010;
        x_t[16] = 21'b000000000001011111101;
        x_t[17] = 21'b000000000001000100000;
        x_t[18] = 21'b111111111110101001010;
        x_t[19] = 21'b111111111100111111100;
        x_t[20] = 21'b111111111101000110001;
        x_t[21] = 21'b000000000010100010111;
        x_t[22] = 21'b000000000011010001100;
        x_t[23] = 21'b000000000011011000101;
        x_t[24] = 21'b000000000010111011101;
        x_t[25] = 21'b000000000010111101111;
        x_t[26] = 21'b000000000001011100011;
        x_t[27] = 21'b000000000001010000010;
        x_t[28] = 21'b000000000010010111100;
        x_t[29] = 21'b000000000010110111110;
        x_t[30] = 21'b000000000011001000110;
        x_t[31] = 21'b000000000001010011101;
        x_t[32] = 21'b000000000001101011000;
        x_t[33] = 21'b000000000001110000100;
        x_t[34] = 21'b000000000001000001010;
        x_t[35] = 21'b111111111111101111010;
        x_t[36] = 21'b000000000000100001011;
        x_t[37] = 21'b111111111100001100010;
        x_t[38] = 21'b000000000010100000101;
        x_t[39] = 21'b111111111111110110111;
        x_t[40] = 21'b000000000100010010110;
        x_t[41] = 21'b111111111011000010000;
        x_t[42] = 21'b000000000101000100100;
        x_t[43] = 21'b000000000010100001001;
        x_t[44] = 21'b000000000101010011000;
        x_t[45] = 21'b111111111101010101010;
        x_t[46] = 21'b000000000101000011001;
        x_t[47] = 21'b000000000010010010000;
        x_t[48] = 21'b000000000001000000110;
        x_t[49] = 21'b000000000000000100111;
        x_t[50] = 21'b111111111101110100101;
        x_t[51] = 21'b111111111010101011011;
        x_t[52] = 21'b111111111010000010101;
        x_t[53] = 21'b111111111001011100111;
        x_t[54] = 21'b111111111011110111011;
        x_t[55] = 21'b000000000011011001011;
        x_t[56] = 21'b000000000010101000110;
        x_t[57] = 21'b111111111101001111000;
        x_t[58] = 21'b111111111000010110110;
        x_t[59] = 21'b111111111010111111100;
        x_t[60] = 21'b000000000010101011101;
        x_t[61] = 21'b000000000000100100101;
        x_t[62] = 21'b111111111011010000001;
        x_t[63] = 21'b000000000001101001111;
        
        h_t_prev[0] = 21'b000000000011111010111;
        h_t_prev[1] = 21'b000000000100000001000;
        h_t_prev[2] = 21'b000000000001110001011;
        h_t_prev[3] = 21'b000000000010110101010;
        h_t_prev[4] = 21'b000000000001010100111;
        h_t_prev[5] = 21'b111111111111111101011;
        h_t_prev[6] = 21'b000000000000000011000;
        h_t_prev[7] = 21'b000000000101000110010;
        h_t_prev[8] = 21'b000000000011000101101;
        h_t_prev[9] = 21'b000000000010101100010;
        h_t_prev[10] = 21'b000000000010001110100;
        h_t_prev[11] = 21'b111111111111110101000;
        h_t_prev[12] = 21'b111111111110110111001;
        h_t_prev[13] = 21'b111111111110001110010;
        h_t_prev[14] = 21'b000000000011101101111;
        h_t_prev[15] = 21'b000000000010011011010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 31 timeout!");
                $fdisplay(fd_cycles, "Test Vector  31: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  31: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 31");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 32
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000001100001111;
        x_t[1] = 21'b000000000010100100000;
        x_t[2] = 21'b111111111111110011001;
        x_t[3] = 21'b000000000010010011011;
        x_t[4] = 21'b000000000000110001100;
        x_t[5] = 21'b111111111111000000011;
        x_t[6] = 21'b111111111111010111100;
        x_t[7] = 21'b000000000011100101101;
        x_t[8] = 21'b000000000001110011001;
        x_t[9] = 21'b000000000001100110001;
        x_t[10] = 21'b000000000001000101001;
        x_t[11] = 21'b111111111111010110011;
        x_t[12] = 21'b111111111111000010111;
        x_t[13] = 21'b111111111101100101011;
        x_t[14] = 21'b000000000010110011111;
        x_t[15] = 21'b000000000001010100000;
        x_t[16] = 21'b000000000000010000010;
        x_t[17] = 21'b111111111111110101001;
        x_t[18] = 21'b111111111110001001101;
        x_t[19] = 21'b111111111101100000100;
        x_t[20] = 21'b111111111101111000001;
        x_t[21] = 21'b000000000001000010001;
        x_t[22] = 21'b000000000010000010001;
        x_t[23] = 21'b000000000010011011101;
        x_t[24] = 21'b000000000001101100100;
        x_t[25] = 21'b000000000001110000001;
        x_t[26] = 21'b000000000000100101011;
        x_t[27] = 21'b000000000000001101011;
        x_t[28] = 21'b000000000001101000010;
        x_t[29] = 21'b000000000000100110010;
        x_t[30] = 21'b000000000001111010110;
        x_t[31] = 21'b000000000001000001111;
        x_t[32] = 21'b000000000001001111110;
        x_t[33] = 21'b000000000001110000100;
        x_t[34] = 21'b000000000000100100101;
        x_t[35] = 21'b111111111111000010111;
        x_t[36] = 21'b000000000000010111100;
        x_t[37] = 21'b111111111011100011100;
        x_t[38] = 21'b111111111111110101010;
        x_t[39] = 21'b000000000000110001101;
        x_t[40] = 21'b000000000010011011001;
        x_t[41] = 21'b111111111101100010000;
        x_t[42] = 21'b000000000011001101111;
        x_t[43] = 21'b111111111110000011111;
        x_t[44] = 21'b000000000010111100010;
        x_t[45] = 21'b111111111111101000011;
        x_t[46] = 21'b000000000010111100100;
        x_t[47] = 21'b000000000001101010010;
        x_t[48] = 21'b000000000001000000110;
        x_t[49] = 21'b111111111111010010000;
        x_t[50] = 21'b111111111101101111111;
        x_t[51] = 21'b111111111011010110111;
        x_t[52] = 21'b111111111011000101001;
        x_t[53] = 21'b111111111010101010110;
        x_t[54] = 21'b111111111100011011010;
        x_t[55] = 21'b000000000010101110010;
        x_t[56] = 21'b000000000001111001100;
        x_t[57] = 21'b111111111100101000101;
        x_t[58] = 21'b111111111001000110110;
        x_t[59] = 21'b111111111011000111011;
        x_t[60] = 21'b000000000001110110000;
        x_t[61] = 21'b111111111111000001010;
        x_t[62] = 21'b111111111001110000000;
        x_t[63] = 21'b000000000001011000010;
        
        h_t_prev[0] = 21'b000000000001100001111;
        h_t_prev[1] = 21'b000000000010100100000;
        h_t_prev[2] = 21'b111111111111110011001;
        h_t_prev[3] = 21'b000000000010010011011;
        h_t_prev[4] = 21'b000000000000110001100;
        h_t_prev[5] = 21'b111111111111000000011;
        h_t_prev[6] = 21'b111111111111010111100;
        h_t_prev[7] = 21'b000000000011100101101;
        h_t_prev[8] = 21'b000000000001110011001;
        h_t_prev[9] = 21'b000000000001100110001;
        h_t_prev[10] = 21'b000000000001000101001;
        h_t_prev[11] = 21'b111111111111010110011;
        h_t_prev[12] = 21'b111111111111000010111;
        h_t_prev[13] = 21'b111111111101100101011;
        h_t_prev[14] = 21'b000000000010110011111;
        h_t_prev[15] = 21'b000000000001010100000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 32 timeout!");
                $fdisplay(fd_cycles, "Test Vector  32: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  32: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 32");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 33
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111110101011011;
        x_t[1] = 21'b111111111110100101100;
        x_t[2] = 21'b111111111110000011011;
        x_t[3] = 21'b111111111110001001100;
        x_t[4] = 21'b111111111101011101011;
        x_t[5] = 21'b111111111011011101000;
        x_t[6] = 21'b111111111010111111011;
        x_t[7] = 21'b111111111111100111001;
        x_t[8] = 21'b111111111110000101111;
        x_t[9] = 21'b111111111101100110100;
        x_t[10] = 21'b111111111101011111001;
        x_t[11] = 21'b111111111100101001001;
        x_t[12] = 21'b111111111011100100100;
        x_t[13] = 21'b111111111001000000011;
        x_t[14] = 21'b111111111111101011011;
        x_t[15] = 21'b111111111110010111111;
        x_t[16] = 21'b111111111101110001101;
        x_t[17] = 21'b111111111101001000011;
        x_t[18] = 21'b111111111101001010011;
        x_t[19] = 21'b111111111100101001100;
        x_t[20] = 21'b111111111100000111100;
        x_t[21] = 21'b111111111110101111110;
        x_t[22] = 21'b111111111101010001100;
        x_t[23] = 21'b111111111110001011000;
        x_t[24] = 21'b111111111110101001101;
        x_t[25] = 21'b111111111110110010100;
        x_t[26] = 21'b111111111100110000011;
        x_t[27] = 21'b111111111101010000110;
        x_t[28] = 21'b111111111101010011010;
        x_t[29] = 21'b111111111110110101111;
        x_t[30] = 21'b111111111101001010011;
        x_t[31] = 21'b111111111110101111100;
        x_t[32] = 21'b111111111110000111111;
        x_t[33] = 21'b111111111101001000011;
        x_t[34] = 21'b111111111100011010000;
        x_t[35] = 21'b111111111011101110110;
        x_t[36] = 21'b111111111011100011011;
        x_t[37] = 21'b111111111000010111101;
        x_t[38] = 21'b111111111110001011011;
        x_t[39] = 21'b111111111000110110101;
        x_t[40] = 21'b111111111110000000100;
        x_t[41] = 21'b111111111010100110010;
        x_t[42] = 21'b111111111111100000110;
        x_t[43] = 21'b111111111110101111110;
        x_t[44] = 21'b111111111011100001011;
        x_t[45] = 21'b111111111011000010010;
        x_t[46] = 21'b111111111111101101010;
        x_t[47] = 21'b111111111111000001001;
        x_t[48] = 21'b111111111110011010000;
        x_t[49] = 21'b111111111111010010000;
        x_t[50] = 21'b111111111110000111110;
        x_t[51] = 21'b111111111110010011010;
        x_t[52] = 21'b111111111110010001110;
        x_t[53] = 21'b111111111101000001001;
        x_t[54] = 21'b111111111100100001010;
        x_t[55] = 21'b111111111110111100100;
        x_t[56] = 21'b111111111111110000000;
        x_t[57] = 21'b111111111111110001000;
        x_t[58] = 21'b000000000000001100011;
        x_t[59] = 21'b000000000000001011001;
        x_t[60] = 21'b111111111110101110101;
        x_t[61] = 21'b111111111101101110100;
        x_t[62] = 21'b111111111110100011000;
        x_t[63] = 21'b111111111100000101011;
        
        h_t_prev[0] = 21'b111111111110101011011;
        h_t_prev[1] = 21'b111111111110100101100;
        h_t_prev[2] = 21'b111111111110000011011;
        h_t_prev[3] = 21'b111111111110001001100;
        h_t_prev[4] = 21'b111111111101011101011;
        h_t_prev[5] = 21'b111111111011011101000;
        h_t_prev[6] = 21'b111111111010111111011;
        h_t_prev[7] = 21'b111111111111100111001;
        h_t_prev[8] = 21'b111111111110000101111;
        h_t_prev[9] = 21'b111111111101100110100;
        h_t_prev[10] = 21'b111111111101011111001;
        h_t_prev[11] = 21'b111111111100101001001;
        h_t_prev[12] = 21'b111111111011100100100;
        h_t_prev[13] = 21'b111111111001000000011;
        h_t_prev[14] = 21'b111111111111101011011;
        h_t_prev[15] = 21'b111111111110010111111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 33 timeout!");
                $fdisplay(fd_cycles, "Test Vector  33: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  33: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 33");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 34
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111100011100011;
        x_t[1] = 21'b111111111100011100100;
        x_t[2] = 21'b111111111011110110101;
        x_t[3] = 21'b111111111011101010000;
        x_t[4] = 21'b111111111011011010000;
        x_t[5] = 21'b111111111001111001001;
        x_t[6] = 21'b111111111001111010111;
        x_t[7] = 21'b111111111110101010000;
        x_t[8] = 21'b111111111100111101101;
        x_t[9] = 21'b111111111100010001010;
        x_t[10] = 21'b111111111100010000111;
        x_t[11] = 21'b111111111100000000011;
        x_t[12] = 21'b111111111011110000001;
        x_t[13] = 21'b111111111010001011010;
        x_t[14] = 21'b111111111110110001011;
        x_t[15] = 21'b111111111101101111001;
        x_t[16] = 21'b111111111101000101001;
        x_t[17] = 21'b111111111100100101110;
        x_t[18] = 21'b111111111101001111101;
        x_t[19] = 21'b111111111101100101111;
        x_t[20] = 21'b111111111101010010101;
        x_t[21] = 21'b111111111101001111000;
        x_t[22] = 21'b111111111011110101100;
        x_t[23] = 21'b111111111100101110010;
        x_t[24] = 21'b111111111101010100011;
        x_t[25] = 21'b111111111101011000011;
        x_t[26] = 21'b111111111010110001110;
        x_t[27] = 21'b111111111011010110111;
        x_t[28] = 21'b111111111011110001101;
        x_t[29] = 21'b111111111101000001011;
        x_t[30] = 21'b111111111011010001011;
        x_t[31] = 21'b111111111100111100001;
        x_t[32] = 21'b111111111011111111101;
        x_t[33] = 21'b111111111011000010010;
        x_t[34] = 21'b111111111010010100101;
        x_t[35] = 21'b111111111001101001100;
        x_t[36] = 21'b111111111001110110000;
        x_t[37] = 21'b111111111000011111110;
        x_t[38] = 21'b111111111100010111011;
        x_t[39] = 21'b111111111001100010110;
        x_t[40] = 21'b111111111100011110110;
        x_t[41] = 21'b111111111100110001010;
        x_t[42] = 21'b111111111100000101011;
        x_t[43] = 21'b111111111001010000101;
        x_t[44] = 21'b111111111001110111010;
        x_t[45] = 21'b111111111101000101111;
        x_t[46] = 21'b111111111110010000000;
        x_t[47] = 21'b111111111110111100001;
        x_t[48] = 21'b111111111111000100111;
        x_t[49] = 21'b000000000000011100001;
        x_t[50] = 21'b111111111111001010010;
        x_t[51] = 21'b111111111111111000101;
        x_t[52] = 21'b111111111111111101010;
        x_t[53] = 21'b111111111110111011101;
        x_t[54] = 21'b111111111110101011001;
        x_t[55] = 21'b111111111111101100000;
        x_t[56] = 21'b000000000000110000100;
        x_t[57] = 21'b000000000001011011101;
        x_t[58] = 21'b000000000001110101001;
        x_t[59] = 21'b000000000010000001100;
        x_t[60] = 21'b111111111111010001001;
        x_t[61] = 21'b111111111110110100111;
        x_t[62] = 21'b000000000000001010100;
        x_t[63] = 21'b111111111101101010101;
        
        h_t_prev[0] = 21'b111111111100011100011;
        h_t_prev[1] = 21'b111111111100011100100;
        h_t_prev[2] = 21'b111111111011110110101;
        h_t_prev[3] = 21'b111111111011101010000;
        h_t_prev[4] = 21'b111111111011011010000;
        h_t_prev[5] = 21'b111111111001111001001;
        h_t_prev[6] = 21'b111111111001111010111;
        h_t_prev[7] = 21'b111111111110101010000;
        h_t_prev[8] = 21'b111111111100111101101;
        h_t_prev[9] = 21'b111111111100010001010;
        h_t_prev[10] = 21'b111111111100010000111;
        h_t_prev[11] = 21'b111111111100000000011;
        h_t_prev[12] = 21'b111111111011110000001;
        h_t_prev[13] = 21'b111111111010001011010;
        h_t_prev[14] = 21'b111111111110110001011;
        h_t_prev[15] = 21'b111111111101101111001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 34 timeout!");
                $fdisplay(fd_cycles, "Test Vector  34: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  34: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 34");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 35
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111100001101101;
        x_t[1] = 21'b111111111100000100000;
        x_t[2] = 21'b111111111011011001100;
        x_t[3] = 21'b111111111011101010000;
        x_t[4] = 21'b111111111011011010000;
        x_t[5] = 21'b111111111010011010011;
        x_t[6] = 21'b111111111001101110100;
        x_t[7] = 21'b111111111110001011100;
        x_t[8] = 21'b111111111101000010110;
        x_t[9] = 21'b111111111100111001011;
        x_t[10] = 21'b111111111101100100000;
        x_t[11] = 21'b111111111101110101100;
        x_t[12] = 21'b111111111101010011101;
        x_t[13] = 21'b111111111100010011101;
        x_t[14] = 21'b111111111101110010001;
        x_t[15] = 21'b111111111110001000101;
        x_t[16] = 21'b111111111110001010100;
        x_t[17] = 21'b111111111101110100110;
        x_t[18] = 21'b111111111110101001010;
        x_t[19] = 21'b111111111111010011110;
        x_t[20] = 21'b111111111111000011010;
        x_t[21] = 21'b111111111100111011101;
        x_t[22] = 21'b111111111011010101110;
        x_t[23] = 21'b111111111100010100001;
        x_t[24] = 21'b111111111101000010001;
        x_t[25] = 21'b111111111101000101110;
        x_t[26] = 21'b111111111011000010101;
        x_t[27] = 21'b111111111011011010111;
        x_t[28] = 21'b111111111011001011110;
        x_t[29] = 21'b111111111100110101000;
        x_t[30] = 21'b111111111011001101011;
        x_t[31] = 21'b111111111101111010010;
        x_t[32] = 21'b111111111101000011110;
        x_t[33] = 21'b111111111100010000111;
        x_t[34] = 21'b111111111011100000110;
        x_t[35] = 21'b111111111010110011100;
        x_t[36] = 21'b111111111011000000100;
        x_t[37] = 21'b111111111000110000001;
        x_t[38] = 21'b111111111101010011111;
        x_t[39] = 21'b111111111011011000010;
        x_t[40] = 21'b111111111110011011110;
        x_t[41] = 21'b111111111111101101001;
        x_t[42] = 21'b111111111110101011011;
        x_t[43] = 21'b111111110111011000000;
        x_t[44] = 21'b111111111011011011111;
        x_t[45] = 21'b111111111110001011100;
        x_t[46] = 21'b000000000000000001111;
        x_t[47] = 21'b000000000000100100101;
        x_t[48] = 21'b000000000000110111010;
        x_t[49] = 21'b000000000010100111001;
        x_t[50] = 21'b000000000001001010100;
        x_t[51] = 21'b000000000001011001010;
        x_t[52] = 21'b000000000001001111001;
        x_t[53] = 21'b000000000000011010010;
        x_t[54] = 21'b000000000000100011000;
        x_t[55] = 21'b000000000001110110001;
        x_t[56] = 21'b000000000010111110010;
        x_t[57] = 21'b000000000011011011100;
        x_t[58] = 21'b000000000010111010111;
        x_t[59] = 21'b000000000011100000010;
        x_t[60] = 21'b000000000001010011100;
        x_t[61] = 21'b000000000001000001101;
        x_t[62] = 21'b000000000010000100101;
        x_t[63] = 21'b000000000000011010101;
        
        h_t_prev[0] = 21'b111111111100001101101;
        h_t_prev[1] = 21'b111111111100000100000;
        h_t_prev[2] = 21'b111111111011011001100;
        h_t_prev[3] = 21'b111111111011101010000;
        h_t_prev[4] = 21'b111111111011011010000;
        h_t_prev[5] = 21'b111111111010011010011;
        h_t_prev[6] = 21'b111111111001101110100;
        h_t_prev[7] = 21'b111111111110001011100;
        h_t_prev[8] = 21'b111111111101000010110;
        h_t_prev[9] = 21'b111111111100111001011;
        h_t_prev[10] = 21'b111111111101100100000;
        h_t_prev[11] = 21'b111111111101110101100;
        h_t_prev[12] = 21'b111111111101010011101;
        h_t_prev[13] = 21'b111111111100010011101;
        h_t_prev[14] = 21'b111111111101110010001;
        h_t_prev[15] = 21'b111111111110001000101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 35 timeout!");
                $fdisplay(fd_cycles, "Test Vector  35: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  35: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 35");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 36
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111101100110011;
        x_t[1] = 21'b111111111110101010100;
        x_t[2] = 21'b111111111110010110111;
        x_t[3] = 21'b111111111110100001110;
        x_t[4] = 21'b111111111110010101000;
        x_t[5] = 21'b111111111101011100100;
        x_t[6] = 21'b111111111100111011111;
        x_t[7] = 21'b000000000000101001010;
        x_t[8] = 21'b111111111111110010001;
        x_t[9] = 21'b111111111111110010110;
        x_t[10] = 21'b000000000000100010111;
        x_t[11] = 21'b000000000000101101000;
        x_t[12] = 21'b111111111111110111100;
        x_t[13] = 21'b111111111110011011111;
        x_t[14] = 21'b000000000000111111110;
        x_t[15] = 21'b000000000000111111101;
        x_t[16] = 21'b000000000001000001111;
        x_t[17] = 21'b000000000000101011011;
        x_t[18] = 21'b000000000001010010000;
        x_t[19] = 21'b000000000001011101001;
        x_t[20] = 21'b000000000001000110101;
        x_t[21] = 21'b111111111110011001101;
        x_t[22] = 21'b111111111100111011011;
        x_t[23] = 21'b111111111101011100101;
        x_t[24] = 21'b111111111110011010011;
        x_t[25] = 21'b111111111110100011000;
        x_t[26] = 21'b111111111101100011001;
        x_t[27] = 21'b111111111101101000011;
        x_t[28] = 21'b111111111100101101011;
        x_t[29] = 21'b111111111110001100010;
        x_t[30] = 21'b111111111101000010100;
        x_t[31] = 21'b000000000000001100101;
        x_t[32] = 21'b111111111111110100111;
        x_t[33] = 21'b111111111110111100001;
        x_t[34] = 21'b111111111101111110000;
        x_t[35] = 21'b111111111101101111000;
        x_t[36] = 21'b111111111101111000011;
        x_t[37] = 21'b111111111010010110000;
        x_t[38] = 21'b111111111111111010010;
        x_t[39] = 21'b111111111100111111001;
        x_t[40] = 21'b000000000000110011111;
        x_t[41] = 21'b111111111111011111001;
        x_t[42] = 21'b000000000001010001011;
        x_t[43] = 21'b111111111110101111110;
        x_t[44] = 21'b111111111110001110101;
        x_t[45] = 21'b111111111111101000011;
        x_t[46] = 21'b000000000010111100100;
        x_t[47] = 21'b000000000011100110101;
        x_t[48] = 21'b000000000011100010110;
        x_t[49] = 21'b000000000101000100101;
        x_t[50] = 21'b000000000011110101100;
        x_t[51] = 21'b000000000011010110111;
        x_t[52] = 21'b000000000010110101011;
        x_t[53] = 21'b000000000001110011011;
        x_t[54] = 21'b000000000010010100111;
        x_t[55] = 21'b000000000100100010110;
        x_t[56] = 21'b000000000101100001100;
        x_t[57] = 21'b000000000101110101000;
        x_t[58] = 21'b000000000100001101110;
        x_t[59] = 21'b000000000100011011100;
        x_t[60] = 21'b000000000100010111000;
        x_t[61] = 21'b000000000100001000010;
        x_t[62] = 21'b000000000100001001110;
        x_t[63] = 21'b000000000011110010010;
        
        h_t_prev[0] = 21'b111111111101100110011;
        h_t_prev[1] = 21'b111111111110101010100;
        h_t_prev[2] = 21'b111111111110010110111;
        h_t_prev[3] = 21'b111111111110100001110;
        h_t_prev[4] = 21'b111111111110010101000;
        h_t_prev[5] = 21'b111111111101011100100;
        h_t_prev[6] = 21'b111111111100111011111;
        h_t_prev[7] = 21'b000000000000101001010;
        h_t_prev[8] = 21'b111111111111110010001;
        h_t_prev[9] = 21'b111111111111110010110;
        h_t_prev[10] = 21'b000000000000100010111;
        h_t_prev[11] = 21'b000000000000101101000;
        h_t_prev[12] = 21'b111111111111110111100;
        h_t_prev[13] = 21'b111111111110011011111;
        h_t_prev[14] = 21'b000000000000111111110;
        h_t_prev[15] = 21'b000000000000111111101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 36 timeout!");
                $fdisplay(fd_cycles, "Test Vector  36: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  36: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 36");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 37
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111111100001101;
        x_t[1] = 21'b000000000000101110101;
        x_t[2] = 21'b111111111111110111111;
        x_t[3] = 21'b111111111111100000100;
        x_t[4] = 21'b111111111111000010011;
        x_t[5] = 21'b111111111110001000111;
        x_t[6] = 21'b111111111101111010001;
        x_t[7] = 21'b000000000010111100111;
        x_t[8] = 21'b000000000001011001010;
        x_t[9] = 21'b000000000001000011000;
        x_t[10] = 21'b000000000001001110111;
        x_t[11] = 21'b000000000000001110100;
        x_t[12] = 21'b111111111111101011111;
        x_t[13] = 21'b111111111100110101101;
        x_t[14] = 21'b000000000010111001001;
        x_t[15] = 21'b000000000010011011010;
        x_t[16] = 21'b000000000001111101011;
        x_t[17] = 21'b000000000001010111110;
        x_t[18] = 21'b000000000001100111000;
        x_t[19] = 21'b000000000001001100101;
        x_t[20] = 21'b000000000000001000000;
        x_t[21] = 21'b111111111110010100001;
        x_t[22] = 21'b111111111101010100110;
        x_t[23] = 21'b111111111101101110000;
        x_t[24] = 21'b111111111110011101011;
        x_t[25] = 21'b111111111110101100011;
        x_t[26] = 21'b111111111101100111011;
        x_t[27] = 21'b111111111110000011111;
        x_t[28] = 21'b111111111101001100111;
        x_t[29] = 21'b111111111111110100010;
        x_t[30] = 21'b111111111100001011111;
        x_t[31] = 21'b000000000000011110011;
        x_t[32] = 21'b111111111111110000011;
        x_t[33] = 21'b111111111110100000011;
        x_t[34] = 21'b111111111101101010111;
        x_t[35] = 21'b111111111101010110011;
        x_t[36] = 21'b111111111110000010011;
        x_t[37] = 21'b111111111010011110010;
        x_t[38] = 21'b000000000000011101101;
        x_t[39] = 21'b111111111100011010011;
        x_t[40] = 21'b000000000001101111101;
        x_t[41] = 21'b111111111101001101001;
        x_t[42] = 21'b000000000000111001101;
        x_t[43] = 21'b111111111100010110001;
        x_t[44] = 21'b111111111110111011010;
        x_t[45] = 21'b111111111110101010011;
        x_t[46] = 21'b000000000011110101011;
        x_t[47] = 21'b000000000100001110011;
        x_t[48] = 21'b000000000100001101101;
        x_t[49] = 21'b000000000101010010100;
        x_t[50] = 21'b000000000100000011110;
        x_t[51] = 21'b000000000011010010000;
        x_t[52] = 21'b000000000010100000111;
        x_t[53] = 21'b000000000000111011101;
        x_t[54] = 21'b000000000000100011000;
        x_t[55] = 21'b000000000101011111001;
        x_t[56] = 21'b000000000110001100100;
        x_t[57] = 21'b000000000110101100011;
        x_t[58] = 21'b000000000100000000101;
        x_t[59] = 21'b000000000011011000011;
        x_t[60] = 21'b000000000110110100001;
        x_t[61] = 21'b000000000110001000100;
        x_t[62] = 21'b000000000100110110001;
        x_t[63] = 21'b000000000101100000011;
        
        h_t_prev[0] = 21'b111111111111100001101;
        h_t_prev[1] = 21'b000000000000101110101;
        h_t_prev[2] = 21'b111111111111110111111;
        h_t_prev[3] = 21'b111111111111100000100;
        h_t_prev[4] = 21'b111111111111000010011;
        h_t_prev[5] = 21'b111111111110001000111;
        h_t_prev[6] = 21'b111111111101111010001;
        h_t_prev[7] = 21'b000000000010111100111;
        h_t_prev[8] = 21'b000000000001011001010;
        h_t_prev[9] = 21'b000000000001000011000;
        h_t_prev[10] = 21'b000000000001001110111;
        h_t_prev[11] = 21'b000000000000001110100;
        h_t_prev[12] = 21'b111111111111101011111;
        h_t_prev[13] = 21'b111111111100110101101;
        h_t_prev[14] = 21'b000000000010111001001;
        h_t_prev[15] = 21'b000000000010011011010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 37 timeout!");
                $fdisplay(fd_cycles, "Test Vector  37: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  37: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 37");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 38
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000000010011000;
        x_t[1] = 21'b000000000000001100011;
        x_t[2] = 21'b111111111111000111011;
        x_t[3] = 21'b111111111110010011010;
        x_t[4] = 21'b111111111101101100100;
        x_t[5] = 21'b111111111101000000110;
        x_t[6] = 21'b111111111101001000010;
        x_t[7] = 21'b000000000011000111000;
        x_t[8] = 21'b000000000001001111000;
        x_t[9] = 21'b000000000000010101111;
        x_t[10] = 21'b111111111111111011110;
        x_t[11] = 21'b111111111110010100001;
        x_t[12] = 21'b111111111110011001111;
        x_t[13] = 21'b111111111100011010011;
        x_t[14] = 21'b000000000011011110000;
        x_t[15] = 21'b000000000010100101011;
        x_t[16] = 21'b000000000001101110100;
        x_t[17] = 21'b000000000000111111001;
        x_t[18] = 21'b000000000001000010001;
        x_t[19] = 21'b000000000000100000101;
        x_t[20] = 21'b111111111111111011100;
        x_t[21] = 21'b111111111110101010010;
        x_t[22] = 21'b111111111101100100101;
        x_t[23] = 21'b111111111110001011000;
        x_t[24] = 21'b111111111111000010000;
        x_t[25] = 21'b111111111111001110100;
        x_t[26] = 21'b111111111101100111011;
        x_t[27] = 21'b111111111110001111101;
        x_t[28] = 21'b111111111101101100011;
        x_t[29] = 21'b000000000000110110111;
        x_t[30] = 21'b111111111101100101101;
        x_t[31] = 21'b000000000000011110011;
        x_t[32] = 21'b000000000000000010100;
        x_t[33] = 21'b111111111110110111100;
        x_t[34] = 21'b111111111101110100100;
        x_t[35] = 21'b111111111101101111000;
        x_t[36] = 21'b111111111110000111011;
        x_t[37] = 21'b111111111010101110100;
        x_t[38] = 21'b000000000010111110111;
        x_t[39] = 21'b111111111101100011111;
        x_t[40] = 21'b000000000011100111010;
        x_t[41] = 21'b000000000000110010101;
        x_t[42] = 21'b000000000010111100001;
        x_t[43] = 21'b111111111010011101011;
        x_t[44] = 21'b000000000000001001100;
        x_t[45] = 21'b111111111110100010110;
        x_t[46] = 21'b000000000101101100101;
        x_t[47] = 21'b000000000101101100111;
        x_t[48] = 21'b000000000101011110101;
        x_t[49] = 21'b000000000110011000000;
        x_t[50] = 21'b000000000100101001110;
        x_t[51] = 21'b000000000011110011110;
        x_t[52] = 21'b000000000011001001111;
        x_t[53] = 21'b000000000001010111100;
        x_t[54] = 21'b000000000000011101000;
        x_t[55] = 21'b000000000111001011001;
        x_t[56] = 21'b000000000111011110001;
        x_t[57] = 21'b000000000111110000101;
        x_t[58] = 21'b000000000100011010111;
        x_t[59] = 21'b000000000011110000000;
        x_t[60] = 21'b000000001000010100000;
        x_t[61] = 21'b000000000111001010110;
        x_t[62] = 21'b000000000100101110110;
        x_t[63] = 21'b000000000101101101100;
        
        h_t_prev[0] = 21'b000000000000010011000;
        h_t_prev[1] = 21'b000000000000001100011;
        h_t_prev[2] = 21'b111111111111000111011;
        h_t_prev[3] = 21'b111111111110010011010;
        h_t_prev[4] = 21'b111111111101101100100;
        h_t_prev[5] = 21'b111111111101000000110;
        h_t_prev[6] = 21'b111111111101001000010;
        h_t_prev[7] = 21'b000000000011000111000;
        h_t_prev[8] = 21'b000000000001001111000;
        h_t_prev[9] = 21'b000000000000010101111;
        h_t_prev[10] = 21'b111111111111111011110;
        h_t_prev[11] = 21'b111111111110010100001;
        h_t_prev[12] = 21'b111111111110011001111;
        h_t_prev[13] = 21'b111111111100011010011;
        h_t_prev[14] = 21'b000000000011011110000;
        h_t_prev[15] = 21'b000000000010100101011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 38 timeout!");
                $fdisplay(fd_cycles, "Test Vector  38: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  38: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 38");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 39
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000010011000010;
        x_t[1] = 21'b000000000010010000100;
        x_t[2] = 21'b000000000000101101011;
        x_t[3] = 21'b111111111111101010010;
        x_t[4] = 21'b111111111110111101011;
        x_t[5] = 21'b111111111101111000010;
        x_t[6] = 21'b111111111101110011111;
        x_t[7] = 21'b000000000101100100111;
        x_t[8] = 21'b000000000011100100100;
        x_t[9] = 21'b000000000010011000001;
        x_t[10] = 21'b000000000001011000101;
        x_t[11] = 21'b111111111111101010110;
        x_t[12] = 21'b111111111111011010010;
        x_t[13] = 21'b111111111101101100001;
        x_t[14] = 21'b000000000101111100010;
        x_t[15] = 21'b000000000100111110000;
        x_t[16] = 21'b000000000011101010011;
        x_t[17] = 21'b000000000010011100111;
        x_t[18] = 21'b000000000010010001010;
        x_t[19] = 21'b000000000001101101100;
        x_t[20] = 21'b000000000001000110101;
        x_t[21] = 21'b111111111111011110101;
        x_t[22] = 21'b111111111110001010101;
        x_t[23] = 21'b111111111110011100100;
        x_t[24] = 21'b111111111111101100101;
        x_t[25] = 21'b111111111111110110111;
        x_t[26] = 21'b111111111110011010000;
        x_t[27] = 21'b111111111110100111010;
        x_t[28] = 21'b111111111101101001010;
        x_t[29] = 21'b000000000001100100101;
        x_t[30] = 21'b111111111111000111010;
        x_t[31] = 21'b000000000001001010110;
        x_t[32] = 21'b000000000001000010001;
        x_t[33] = 21'b111111111111110011101;
        x_t[34] = 21'b111111111110110010011;
        x_t[35] = 21'b111111111110010110100;
        x_t[36] = 21'b111111111101101001100;
        x_t[37] = 21'b111111111010001001110;
        x_t[38] = 21'b000000000011100010010;
        x_t[39] = 21'b111111111100101001001;
        x_t[40] = 21'b000000000011011100011;
        x_t[41] = 21'b111111111110011001101;
        x_t[42] = 21'b000000000001101111000;
        x_t[43] = 21'b111111111011010100010;
        x_t[44] = 21'b000000000001111001001;
        x_t[45] = 21'b111111111111000001101;
        x_t[46] = 21'b000000000110101111111;
        x_t[47] = 21'b000000000110110111100;
        x_t[48] = 21'b000000000110101010111;
        x_t[49] = 21'b000000000111100010001;
        x_t[50] = 21'b000000000101100111101;
        x_t[51] = 21'b000000000100100100001;
        x_t[52] = 21'b000000000100000010001;
        x_t[53] = 21'b000000000010010100110;
        x_t[54] = 21'b000000000001101010111;
        x_t[55] = 21'b000000000111100101000;
        x_t[56] = 21'b000000000111111100010;
        x_t[57] = 21'b000000001000001010001;
        x_t[58] = 21'b000000000101000010001;
        x_t[59] = 21'b000000000100101011010;
        x_t[60] = 21'b000000001001000010000;
        x_t[61] = 21'b000000000111110000000;
        x_t[62] = 21'b000000000101001000101;
        x_t[63] = 21'b000000000110011001100;
        
        h_t_prev[0] = 21'b000000000010011000010;
        h_t_prev[1] = 21'b000000000010010000100;
        h_t_prev[2] = 21'b000000000000101101011;
        h_t_prev[3] = 21'b111111111111101010010;
        h_t_prev[4] = 21'b111111111110111101011;
        h_t_prev[5] = 21'b111111111101111000010;
        h_t_prev[6] = 21'b111111111101110011111;
        h_t_prev[7] = 21'b000000000101100100111;
        h_t_prev[8] = 21'b000000000011100100100;
        h_t_prev[9] = 21'b000000000010011000001;
        h_t_prev[10] = 21'b000000000001011000101;
        h_t_prev[11] = 21'b111111111111101010110;
        h_t_prev[12] = 21'b111111111111011010010;
        h_t_prev[13] = 21'b111111111101101100001;
        h_t_prev[14] = 21'b000000000101111100010;
        h_t_prev[15] = 21'b000000000100111110000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 39 timeout!");
                $fdisplay(fd_cycles, "Test Vector  39: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  39: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 39");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 40
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000001111010101;
        x_t[1] = 21'b000000000010010101011;
        x_t[2] = 21'b000000000000101101011;
        x_t[3] = 21'b000000000000000111010;
        x_t[4] = 21'b111111111111010110101;
        x_t[5] = 21'b111111111110000011011;
        x_t[6] = 21'b111111111110000000011;
        x_t[7] = 21'b000000000101001011011;
        x_t[8] = 21'b000000000011111110011;
        x_t[9] = 21'b000000000010101100010;
        x_t[10] = 21'b000000000010011101001;
        x_t[11] = 21'b000000000000110010001;
        x_t[12] = 21'b000000000000011010101;
        x_t[13] = 21'b111111111110011011111;
        x_t[14] = 21'b000000000101010111010;
        x_t[15] = 21'b000000000101001101010;
        x_t[16] = 21'b000000000100010111000;
        x_t[17] = 21'b000000000011001001010;
        x_t[18] = 21'b000000000010110110001;
        x_t[19] = 21'b000000000010001110100;
        x_t[20] = 21'b000000000001011111101;
        x_t[21] = 21'b111111111110111000000;
        x_t[22] = 21'b111111111101011011000;
        x_t[23] = 21'b111111111101110000111;
        x_t[24] = 21'b111111111110111000111;
        x_t[25] = 21'b111111111111000101010;
        x_t[26] = 21'b111111111101001110000;
        x_t[27] = 21'b111111111101100100011;
        x_t[28] = 21'b111111111100110011110;
        x_t[29] = 21'b000000000000011001110;
        x_t[30] = 21'b111111111110010100100;
        x_t[31] = 21'b000000000000010001000;
        x_t[32] = 21'b111111111111100111010;
        x_t[33] = 21'b111111111110010111001;
        x_t[34] = 21'b111111111101100110001;
        x_t[35] = 21'b111111111100111000110;
        x_t[36] = 21'b111111111100110010111;
        x_t[37] = 21'b111111111001101101010;
        x_t[38] = 21'b000000000001111000011;
        x_t[39] = 21'b111111111011111101000;
        x_t[40] = 21'b000000000001011111011;
        x_t[41] = 21'b111111111110100111100;
        x_t[42] = 21'b000000000010011110100;
        x_t[43] = 21'b111111111000101111110;
        x_t[44] = 21'b000000000001110011101;
        x_t[45] = 21'b111111111110001011100;
        x_t[46] = 21'b000000000100111110000;
        x_t[47] = 21'b000000000101110001111;
        x_t[48] = 21'b000000000101110110100;
        x_t[49] = 21'b000000000111000001110;
        x_t[50] = 21'b000000000101001011001;
        x_t[51] = 21'b000000000011111000101;
        x_t[52] = 21'b000000000011001111000;
        x_t[53] = 21'b000000000001100010101;
        x_t[54] = 21'b000000000001011110111;
        x_t[55] = 21'b000000000110110101100;
        x_t[56] = 21'b000000000111010101100;
        x_t[57] = 21'b000000000111010111000;
        x_t[58] = 21'b000000000100010010001;
        x_t[59] = 21'b000000000011110111111;
        x_t[60] = 21'b000000001001000010000;
        x_t[61] = 21'b000000000111111000010;
        x_t[62] = 21'b000000000101110101000;
        x_t[63] = 21'b000000000111010010110;
        
        h_t_prev[0] = 21'b000000000001111010101;
        h_t_prev[1] = 21'b000000000010010101011;
        h_t_prev[2] = 21'b000000000000101101011;
        h_t_prev[3] = 21'b000000000000000111010;
        h_t_prev[4] = 21'b111111111111010110101;
        h_t_prev[5] = 21'b111111111110000011011;
        h_t_prev[6] = 21'b111111111110000000011;
        h_t_prev[7] = 21'b000000000101001011011;
        h_t_prev[8] = 21'b000000000011111110011;
        h_t_prev[9] = 21'b000000000010101100010;
        h_t_prev[10] = 21'b000000000010011101001;
        h_t_prev[11] = 21'b000000000000110010001;
        h_t_prev[12] = 21'b000000000000011010101;
        h_t_prev[13] = 21'b111111111110011011111;
        h_t_prev[14] = 21'b000000000101010111010;
        h_t_prev[15] = 21'b000000000101001101010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 40 timeout!");
                $fdisplay(fd_cycles, "Test Vector  40: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  40: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 40");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 41
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000000011000000;
        x_t[1] = 21'b000000000001000111001;
        x_t[2] = 21'b000000000000010000010;
        x_t[3] = 21'b111111111111101010010;
        x_t[4] = 21'b111111111111000111100;
        x_t[5] = 21'b111111111101100111101;
        x_t[6] = 21'b111111111101011011000;
        x_t[7] = 21'b000000000011011011011;
        x_t[8] = 21'b000000000011001010110;
        x_t[9] = 21'b000000000010100010010;
        x_t[10] = 21'b000000000010100110111;
        x_t[11] = 21'b000000000001000110100;
        x_t[12] = 21'b111111111111110001110;
        x_t[13] = 21'b111111111100100001010;
        x_t[14] = 21'b000000000100100111111;
        x_t[15] = 21'b000000000100101110101;
        x_t[16] = 21'b000000000011111110010;
        x_t[17] = 21'b000000000010101011101;
        x_t[18] = 21'b000000000010010110100;
        x_t[19] = 21'b000000000001001100101;
        x_t[20] = 21'b111111111111100010100;
        x_t[21] = 21'b111111111111000000010;
        x_t[22] = 21'b111111111101100111110;
        x_t[23] = 21'b111111111101110110110;
        x_t[24] = 21'b111111111111001000000;
        x_t[25] = 21'b111111111111010100110;
        x_t[26] = 21'b111111111101101011101;
        x_t[27] = 21'b111111111101111111111;
        x_t[28] = 21'b111111111101011001100;
        x_t[29] = 21'b000000000000101110100;
        x_t[30] = 21'b111111111110110111101;
        x_t[31] = 21'b000000000000110100100;
        x_t[32] = 21'b000000000000101011100;
        x_t[33] = 21'b111111111111100001001;
        x_t[34] = 21'b111111111110011111011;
        x_t[35] = 21'b111111111110000111101;
        x_t[36] = 21'b111111111101101001100;
        x_t[37] = 21'b111111111011011011011;
        x_t[38] = 21'b000000000010000010011;
        x_t[39] = 21'b111111111100110111111;
        x_t[40] = 21'b000000000010100000101;
        x_t[41] = 21'b111111111101000110001;
        x_t[42] = 21'b000000000011011001110;
        x_t[43] = 21'b111111111101000010000;
        x_t[44] = 21'b000000000001101000011;
        x_t[45] = 21'b111111111101101100100;
        x_t[46] = 21'b000000000100110011101;
        x_t[47] = 21'b000000000101100111111;
        x_t[48] = 21'b000000000101101100111;
        x_t[49] = 21'b000000000110100001010;
        x_t[50] = 21'b000000000101000001100;
        x_t[51] = 21'b000000000011001101001;
        x_t[52] = 21'b000000000010010110101;
        x_t[53] = 21'b000000000000010100101;
        x_t[54] = 21'b000000000000011101000;
        x_t[55] = 21'b000000000111001011001;
        x_t[56] = 21'b000000000111011110001;
        x_t[57] = 21'b000000000110111101011;
        x_t[58] = 21'b000000000011010101001;
        x_t[59] = 21'b000000000011000100101;
        x_t[60] = 21'b000000001000011011110;
        x_t[61] = 21'b000000000111000110101;
        x_t[62] = 21'b000000000101101101101;
        x_t[63] = 21'b000000000110011001100;
        
        h_t_prev[0] = 21'b000000000000011000000;
        h_t_prev[1] = 21'b000000000001000111001;
        h_t_prev[2] = 21'b000000000000010000010;
        h_t_prev[3] = 21'b111111111111101010010;
        h_t_prev[4] = 21'b111111111111000111100;
        h_t_prev[5] = 21'b111111111101100111101;
        h_t_prev[6] = 21'b111111111101011011000;
        h_t_prev[7] = 21'b000000000011011011011;
        h_t_prev[8] = 21'b000000000011001010110;
        h_t_prev[9] = 21'b000000000010100010010;
        h_t_prev[10] = 21'b000000000010100110111;
        h_t_prev[11] = 21'b000000000001000110100;
        h_t_prev[12] = 21'b111111111111110001110;
        h_t_prev[13] = 21'b111111111100100001010;
        h_t_prev[14] = 21'b000000000100100111111;
        h_t_prev[15] = 21'b000000000100101110101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 41 timeout!");
                $fdisplay(fd_cycles, "Test Vector  41: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  41: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 41");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 42
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000010001001011;
        x_t[1] = 21'b000000000011101000101;
        x_t[2] = 21'b000000000010110101010;
        x_t[3] = 21'b000000000010011000010;
        x_t[4] = 21'b000000000001011010000;
        x_t[5] = 21'b111111111111010110101;
        x_t[6] = 21'b111111111101111010001;
        x_t[7] = 21'b000000000110010010101;
        x_t[8] = 21'b000000000101100000011;
        x_t[9] = 21'b000000000100111000100;
        x_t[10] = 21'b000000000100010010100;
        x_t[11] = 21'b000000000010110110101;
        x_t[12] = 21'b000000000000110010001;
        x_t[13] = 21'b111111111100011010011;
        x_t[14] = 21'b000000000111100000011;
        x_t[15] = 21'b000000000110100011101;
        x_t[16] = 21'b000000000101100110011;
        x_t[17] = 21'b000000000100000100100;
        x_t[18] = 21'b000000000011101010110;
        x_t[19] = 21'b000000000010010100000;
        x_t[20] = 21'b000000000000001000000;
        x_t[21] = 21'b111111111111001011011;
        x_t[22] = 21'b111111111110000001001;
        x_t[23] = 21'b111111111110011100100;
        x_t[24] = 21'b111111111111101111101;
        x_t[25] = 21'b000000000000000000010;
        x_t[26] = 21'b111111111111010001000;
        x_t[27] = 21'b111111111111010010100;
        x_t[28] = 21'b111111111110010010001;
        x_t[29] = 21'b000000000001110001001;
        x_t[30] = 21'b111111111111111101111;
        x_t[31] = 21'b000000000010101100010;
        x_t[32] = 21'b000000000010011000100;
        x_t[33] = 21'b000000000001011001011;
        x_t[34] = 21'b000000000000011011001;
        x_t[35] = 21'b111111111111101010011;
        x_t[36] = 21'b111111111110101111001;
        x_t[37] = 21'b111111111100000000000;
        x_t[38] = 21'b000000000010100101110;
        x_t[39] = 21'b111111111101010101010;
        x_t[40] = 21'b000000000010011011001;
        x_t[41] = 21'b111111111100111000010;
        x_t[42] = 21'b000000000011110111011;
        x_t[43] = 21'b111111111110001110110;
        x_t[44] = 21'b000000000011100011010;
        x_t[45] = 21'b000000000000000111010;
        x_t[46] = 21'b000000000110111010010;
        x_t[47] = 21'b000000000111011111010;
        x_t[48] = 21'b000000000110110100011;
        x_t[49] = 21'b000000001000000010101;
        x_t[50] = 21'b000000000110010111001;
        x_t[51] = 21'b000000000100110111011;
        x_t[52] = 21'b000000000100001100011;
        x_t[53] = 21'b000000000010000100000;
        x_t[54] = 21'b000000000010001000111;
        x_t[55] = 21'b000000001000011000110;
        x_t[56] = 21'b000000001000101111110;
        x_t[57] = 21'b000000001000001010001;
        x_t[58] = 21'b000000000100010110100;
        x_t[59] = 21'b000000000100000011110;
        x_t[60] = 21'b000000001000011011110;
        x_t[61] = 21'b000000000111000010100;
        x_t[62] = 21'b000000000101111100011;
        x_t[63] = 21'b000000000110011101111;
        
        h_t_prev[0] = 21'b000000000010001001011;
        h_t_prev[1] = 21'b000000000011101000101;
        h_t_prev[2] = 21'b000000000010110101010;
        h_t_prev[3] = 21'b000000000010011000010;
        h_t_prev[4] = 21'b000000000001011010000;
        h_t_prev[5] = 21'b111111111111010110101;
        h_t_prev[6] = 21'b111111111101111010001;
        h_t_prev[7] = 21'b000000000110010010101;
        h_t_prev[8] = 21'b000000000101100000011;
        h_t_prev[9] = 21'b000000000100111000100;
        h_t_prev[10] = 21'b000000000100010010100;
        h_t_prev[11] = 21'b000000000010110110101;
        h_t_prev[12] = 21'b000000000000110010001;
        h_t_prev[13] = 21'b111111111100011010011;
        h_t_prev[14] = 21'b000000000111100000011;
        h_t_prev[15] = 21'b000000000110100011101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 42 timeout!");
                $fdisplay(fd_cycles, "Test Vector  42: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  42: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 42");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 43
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000010110000111;
        x_t[1] = 21'b000000000011011001111;
        x_t[2] = 21'b000000000010101011101;
        x_t[3] = 21'b000000000010100110110;
        x_t[4] = 21'b000000000001101110001;
        x_t[5] = 21'b000000000000001000100;
        x_t[6] = 21'b111111111111100011111;
        x_t[7] = 21'b000000000100110111000;
        x_t[8] = 21'b000000000100011000001;
        x_t[9] = 21'b000000000100000001011;
        x_t[10] = 21'b000000000011110101010;
        x_t[11] = 21'b000000000011001011000;
        x_t[12] = 21'b000000000001100110110;
        x_t[13] = 21'b111111111110111101111;
        x_t[14] = 21'b000000000101100001111;
        x_t[15] = 21'b000000000101001000001;
        x_t[16] = 21'b000000000100110100110;
        x_t[17] = 21'b000000000011100110111;
        x_t[18] = 21'b000000000100000101001;
        x_t[19] = 21'b000000000011100000111;
        x_t[20] = 21'b000000000010010001101;
        x_t[21] = 21'b111111111110101111110;
        x_t[22] = 21'b111111111101011110010;
        x_t[23] = 21'b111111111110001110000;
        x_t[24] = 21'b111111111111001011001;
        x_t[25] = 21'b111111111111010111111;
        x_t[26] = 21'b111111111110011010000;
        x_t[27] = 21'b111111111110111010111;
        x_t[28] = 21'b111111111110001000110;
        x_t[29] = 21'b000000000001101100111;
        x_t[30] = 21'b111111111111101010011;
        x_t[31] = 21'b000000000001111011100;
        x_t[32] = 21'b000000000000111001001;
        x_t[33] = 21'b000000000000001111011;
        x_t[34] = 21'b111111111111100010000;
        x_t[35] = 21'b111111111110101111001;
        x_t[36] = 21'b111111111110011011010;
        x_t[37] = 21'b111111111100000100001;
        x_t[38] = 21'b000000000011011101010;
        x_t[39] = 21'b111111111110111100001;
        x_t[40] = 21'b000000000101001001000;
        x_t[41] = 21'b000000000011011001100;
        x_t[42] = 21'b000000000101101000000;
        x_t[43] = 21'b111111111110100100110;
        x_t[44] = 21'b000000000011101110100;
        x_t[45] = 21'b000000000001100100001;
        x_t[46] = 21'b000000000101100010010;
        x_t[47] = 21'b000000000101100111111;
        x_t[48] = 21'b000000000100110011110;
        x_t[49] = 21'b000000000110100101111;
        x_t[50] = 21'b000000000100111100110;
        x_t[51] = 21'b000000000100010000110;
        x_t[52] = 21'b000000000100000111010;
        x_t[53] = 21'b000000000010101011000;
        x_t[54] = 21'b000000000010101100111;
        x_t[55] = 21'b000000000110011111111;
        x_t[56] = 21'b000000000111000100011;
        x_t[57] = 21'b000000000110111001001;
        x_t[58] = 21'b000000000100000101000;
        x_t[59] = 21'b000000000100000011110;
        x_t[60] = 21'b000000001000010000010;
        x_t[61] = 21'b000000000111000110101;
        x_t[62] = 21'b000000000110001011001;
        x_t[63] = 21'b000000000110101011001;
        
        h_t_prev[0] = 21'b000000000010110000111;
        h_t_prev[1] = 21'b000000000011011001111;
        h_t_prev[2] = 21'b000000000010101011101;
        h_t_prev[3] = 21'b000000000010100110110;
        h_t_prev[4] = 21'b000000000001101110001;
        h_t_prev[5] = 21'b000000000000001000100;
        h_t_prev[6] = 21'b111111111111100011111;
        h_t_prev[7] = 21'b000000000100110111000;
        h_t_prev[8] = 21'b000000000100011000001;
        h_t_prev[9] = 21'b000000000100000001011;
        h_t_prev[10] = 21'b000000000011110101010;
        h_t_prev[11] = 21'b000000000011001011000;
        h_t_prev[12] = 21'b000000000001100110110;
        h_t_prev[13] = 21'b111111111110111101111;
        h_t_prev[14] = 21'b000000000101100001111;
        h_t_prev[15] = 21'b000000000101001000001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 43 timeout!");
                $fdisplay(fd_cycles, "Test Vector  43: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  43: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 43");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 44
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000010100010000;
        x_t[1] = 21'b000000000010100100000;
        x_t[2] = 21'b000000000001110001011;
        x_t[3] = 21'b000000000001111011010;
        x_t[4] = 21'b000000000001001010111;
        x_t[5] = 21'b111111111111111101011;
        x_t[6] = 21'b000000000001000001010;
        x_t[7] = 21'b000000000011101111110;
        x_t[8] = 21'b000000000011001111111;
        x_t[9] = 21'b000000000010110110010;
        x_t[10] = 21'b000000000011001001001;
        x_t[11] = 21'b000000000011010000001;
        x_t[12] = 21'b000000000010001111110;
        x_t[13] = 21'b000000000001101000010;
        x_t[14] = 21'b000000000011111000011;
        x_t[15] = 21'b000000000011111011111;
        x_t[16] = 21'b000000000011101111011;
        x_t[17] = 21'b000000000011001001010;
        x_t[18] = 21'b000000000100000101001;
        x_t[19] = 21'b000000000100000001111;
        x_t[20] = 21'b000000000100001110111;
        x_t[21] = 21'b111111111111001110001;
        x_t[22] = 21'b111111111101111110000;
        x_t[23] = 21'b111111111110011100100;
        x_t[24] = 21'b111111111111110101110;
        x_t[25] = 21'b000000000000000000010;
        x_t[26] = 21'b111111111111001000100;
        x_t[27] = 21'b111111111111010010100;
        x_t[28] = 21'b111111111110010010001;
        x_t[29] = 21'b000000000010011110111;
        x_t[30] = 21'b000000000000011001001;
        x_t[31] = 21'b000000000010100011100;
        x_t[32] = 21'b000000000001110100001;
        x_t[33] = 21'b000000000001001011100;
        x_t[34] = 21'b000000000000010110011;
        x_t[35] = 21'b111111111111111001001;
        x_t[36] = 21'b111111111111100000110;
        x_t[37] = 21'b111111111101001001011;
        x_t[38] = 21'b000000000011101100011;
        x_t[39] = 21'b000000000001001111001;
        x_t[40] = 21'b000000000100100011000;
        x_t[41] = 21'b000000000101010110110;
        x_t[42] = 21'b000000000101101000000;
        x_t[43] = 21'b000000000000110011011;
        x_t[44] = 21'b000000000010001111100;
        x_t[45] = 21'b000000000011011000010;
        x_t[46] = 21'b000000000100111000110;
        x_t[47] = 21'b000000000101001111000;
        x_t[48] = 21'b000000000100100101100;
        x_t[49] = 21'b000000000110011000000;
        x_t[50] = 21'b000000000101000110011;
        x_t[51] = 21'b000000000100101101110;
        x_t[52] = 21'b000000000101000100101;
        x_t[53] = 21'b000000000100001001101;
        x_t[54] = 21'b000000000100011000110;
        x_t[55] = 21'b000000000101110100110;
        x_t[56] = 21'b000000000110010101001;
        x_t[57] = 21'b000000000110011111101;
        x_t[58] = 21'b000000000100101000000;
        x_t[59] = 21'b000000000100110011001;
        x_t[60] = 21'b000000000111010110110;
        x_t[61] = 21'b000000000110100101100;
        x_t[62] = 21'b000000000110010110010;
        x_t[63] = 21'b000000000101111111001;
        
        h_t_prev[0] = 21'b000000000010100010000;
        h_t_prev[1] = 21'b000000000010100100000;
        h_t_prev[2] = 21'b000000000001110001011;
        h_t_prev[3] = 21'b000000000001111011010;
        h_t_prev[4] = 21'b000000000001001010111;
        h_t_prev[5] = 21'b111111111111111101011;
        h_t_prev[6] = 21'b000000000001000001010;
        h_t_prev[7] = 21'b000000000011101111110;
        h_t_prev[8] = 21'b000000000011001111111;
        h_t_prev[9] = 21'b000000000010110110010;
        h_t_prev[10] = 21'b000000000011001001001;
        h_t_prev[11] = 21'b000000000011010000001;
        h_t_prev[12] = 21'b000000000010001111110;
        h_t_prev[13] = 21'b000000000001101000010;
        h_t_prev[14] = 21'b000000000011111000011;
        h_t_prev[15] = 21'b000000000011111011111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 44 timeout!");
                $fdisplay(fd_cycles, "Test Vector  44: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  44: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 44");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 45
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000011100010001;
        x_t[1] = 21'b000000000011111100001;
        x_t[2] = 21'b000000000011100001000;
        x_t[3] = 21'b000000000011001101011;
        x_t[4] = 21'b000000000010011011101;
        x_t[5] = 21'b000000000001100001010;
        x_t[6] = 21'b000000000010010010001;
        x_t[7] = 21'b000000000101000110010;
        x_t[8] = 21'b000000000100101100110;
        x_t[9] = 21'b000000000100000110011;
        x_t[10] = 21'b000000000100001000110;
        x_t[11] = 21'b000000000011111000111;
        x_t[12] = 21'b000000000011100001101;
        x_t[13] = 21'b000000000010000011100;
        x_t[14] = 21'b000000000100111100111;
        x_t[15] = 21'b000000000100011111011;
        x_t[16] = 21'b000000000100001000001;
        x_t[17] = 21'b000000000011100110111;
        x_t[18] = 21'b000000000100001111110;
        x_t[19] = 21'b000000000100001100110;
        x_t[20] = 21'b000000000100100001101;
        x_t[21] = 21'b111111111111011001001;
        x_t[22] = 21'b111111111101110111101;
        x_t[23] = 21'b111111111110001011000;
        x_t[24] = 21'b111111111111101111101;
        x_t[25] = 21'b000000000000000110100;
        x_t[26] = 21'b111111111111100001111;
        x_t[27] = 21'b111111111111101010000;
        x_t[28] = 21'b111111111110001011111;
        x_t[29] = 21'b000000000001111001011;
        x_t[30] = 21'b000000000000101100101;
        x_t[31] = 21'b000000000011010100010;
        x_t[32] = 21'b000000000010010011111;
        x_t[33] = 21'b000000000001011001011;
        x_t[34] = 21'b000000000000101110010;
        x_t[35] = 21'b000000000000001100111;
        x_t[36] = 21'b000000000000010010100;
        x_t[37] = 21'b111111111110010110111;
        x_t[38] = 21'b000000000100001111101;
        x_t[39] = 21'b000000000000111001000;
        x_t[40] = 21'b000000000101010011111;
        x_t[41] = 21'b000000000010101000111;
        x_t[42] = 21'b000000000011011111101;
        x_t[43] = 21'b000000000010101100000;
        x_t[44] = 21'b000000000010001001111;
        x_t[45] = 21'b000000000011100000000;
        x_t[46] = 21'b000000000100011001110;
        x_t[47] = 21'b000000000100011000010;
        x_t[48] = 21'b000000000011101100010;
        x_t[49] = 21'b000000000101000100101;
        x_t[50] = 21'b000000000011111111000;
        x_t[51] = 21'b000000000011100000100;
        x_t[52] = 21'b000000000011101101101;
        x_t[53] = 21'b000000000010111011110;
        x_t[54] = 21'b000000000011001010110;
        x_t[55] = 21'b000000000100001000111;
        x_t[56] = 21'b000000000100101001101;
        x_t[57] = 21'b000000000100010111001;
        x_t[58] = 21'b000000000010111111010;
        x_t[59] = 21'b000000000010100101000;
        x_t[60] = 21'b000000000101010000100;
        x_t[61] = 21'b000000000011110111101;
        x_t[62] = 21'b000000000100100011101;
        x_t[63] = 21'b000000000010110100110;
        
        h_t_prev[0] = 21'b000000000011100010001;
        h_t_prev[1] = 21'b000000000011111100001;
        h_t_prev[2] = 21'b000000000011100001000;
        h_t_prev[3] = 21'b000000000011001101011;
        h_t_prev[4] = 21'b000000000010011011101;
        h_t_prev[5] = 21'b000000000001100001010;
        h_t_prev[6] = 21'b000000000010010010001;
        h_t_prev[7] = 21'b000000000101000110010;
        h_t_prev[8] = 21'b000000000100101100110;
        h_t_prev[9] = 21'b000000000100000110011;
        h_t_prev[10] = 21'b000000000100001000110;
        h_t_prev[11] = 21'b000000000011111000111;
        h_t_prev[12] = 21'b000000000011100001101;
        h_t_prev[13] = 21'b000000000010000011100;
        h_t_prev[14] = 21'b000000000100111100111;
        h_t_prev[15] = 21'b000000000100011111011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 45 timeout!");
                $fdisplay(fd_cycles, "Test Vector  45: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  45: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 45");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 46
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000011010011011;
        x_t[1] = 21'b000000000100000110000;
        x_t[2] = 21'b000000000011010010100;
        x_t[3] = 21'b000000000010111010001;
        x_t[4] = 21'b000000000001111101011;
        x_t[5] = 21'b000000000001010000101;
        x_t[6] = 21'b000000000001101100110;
        x_t[7] = 21'b000000000101101001111;
        x_t[8] = 21'b000000000100110111001;
        x_t[9] = 21'b000000000100010101100;
        x_t[10] = 21'b000000000100010111100;
        x_t[11] = 21'b000000000011011010010;
        x_t[12] = 21'b000000000011010000001;
        x_t[13] = 21'b000000000001100001100;
        x_t[14] = 21'b000000000101111100010;
        x_t[15] = 21'b000000000100111110000;
        x_t[16] = 21'b000000000100010111000;
        x_t[17] = 21'b000000000011110000110;
        x_t[18] = 21'b000000000100001111110;
        x_t[19] = 21'b000000000100000111010;
        x_t[20] = 21'b000000000100001000100;
        x_t[21] = 21'b111111111111011001001;
        x_t[22] = 21'b111111111110000100010;
        x_t[23] = 21'b111111111101111111100;
        x_t[24] = 21'b111111111111110010101;
        x_t[25] = 21'b000000000000000110100;
        x_t[26] = 21'b111111111111100110001;
        x_t[27] = 21'b111111111111111001110;
        x_t[28] = 21'b111111111110010101011;
        x_t[29] = 21'b000000000001101100111;
        x_t[30] = 21'b000000000001011011100;
        x_t[31] = 21'b000000000011011000101;
        x_t[32] = 21'b000000000010110011110;
        x_t[33] = 21'b000000000001100111010;
        x_t[34] = 21'b000000000000101110010;
        x_t[35] = 21'b000000000000011011110;
        x_t[36] = 21'b000000000000000011101;
        x_t[37] = 21'b111111111110100111010;
        x_t[38] = 21'b000000000101000111001;
        x_t[39] = 21'b000000000000101010011;
        x_t[40] = 21'b000000000100101000100;
        x_t[41] = 21'b000000000001100011010;
        x_t[42] = 21'b000000000011110111011;
        x_t[43] = 21'b000000000100011001110;
        x_t[44] = 21'b000000000010110001000;
        x_t[45] = 21'b000000000101010100000;
        x_t[46] = 21'b000000000101001101100;
        x_t[47] = 21'b000000000101010100000;
        x_t[48] = 21'b000000000100100000110;
        x_t[49] = 21'b000000000101111100010;
        x_t[50] = 21'b000000000101001011001;
        x_t[51] = 21'b000000000100111100010;
        x_t[52] = 21'b000000000101001001110;
        x_t[53] = 21'b000000000100010100110;
        x_t[54] = 21'b000000000100111100101;
        x_t[55] = 21'b000000000100011010001;
        x_t[56] = 21'b000000000101000011011;
        x_t[57] = 21'b000000000101001110101;
        x_t[58] = 21'b000000000100011010111;
        x_t[59] = 21'b000000000100000011110;
        x_t[60] = 21'b000000000100000000000;
        x_t[61] = 21'b000000000010010100011;
        x_t[62] = 21'b000000000011100001000;
        x_t[63] = 21'b000000000001101001111;
        
        h_t_prev[0] = 21'b000000000011010011011;
        h_t_prev[1] = 21'b000000000100000110000;
        h_t_prev[2] = 21'b000000000011010010100;
        h_t_prev[3] = 21'b000000000010111010001;
        h_t_prev[4] = 21'b000000000001111101011;
        h_t_prev[5] = 21'b000000000001010000101;
        h_t_prev[6] = 21'b000000000001101100110;
        h_t_prev[7] = 21'b000000000101101001111;
        h_t_prev[8] = 21'b000000000100110111001;
        h_t_prev[9] = 21'b000000000100010101100;
        h_t_prev[10] = 21'b000000000100010111100;
        h_t_prev[11] = 21'b000000000011011010010;
        h_t_prev[12] = 21'b000000000011010000001;
        h_t_prev[13] = 21'b000000000001100001100;
        h_t_prev[14] = 21'b000000000101111100010;
        h_t_prev[15] = 21'b000000000100111110000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 46 timeout!");
                $fdisplay(fd_cycles, "Test Vector  46: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  46: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 46");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 47
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000100101100001;
        x_t[1] = 21'b000000000101011110000;
        x_t[2] = 21'b000000000100011011010;
        x_t[3] = 21'b000000000100011111101;
        x_t[4] = 21'b000000000011010011010;
        x_t[5] = 21'b000000000001110001111;
        x_t[6] = 21'b000000000001100110101;
        x_t[7] = 21'b000000000110100001111;
        x_t[8] = 21'b000000000101101010101;
        x_t[9] = 21'b000000000110001000110;
        x_t[10] = 21'b000000000110000011001;
        x_t[11] = 21'b000000000101010100101;
        x_t[12] = 21'b000000000100010000100;
        x_t[13] = 21'b000000000010001010011;
        x_t[14] = 21'b000000000101010111010;
        x_t[15] = 21'b000000000101100110101;
        x_t[16] = 21'b000000000101101011010;
        x_t[17] = 21'b000000000101010011100;
        x_t[18] = 21'b000000000101111110011;
        x_t[19] = 21'b000000000101100100101;
        x_t[20] = 21'b000000000100110100011;
        x_t[21] = 21'b111111111111010110011;
        x_t[22] = 21'b111111111110010111011;
        x_t[23] = 21'b111111111110011001100;
        x_t[24] = 21'b111111111111110010101;
        x_t[25] = 21'b000000000000000110100;
        x_t[26] = 21'b000000000000001100001;
        x_t[27] = 21'b000000000000000001101;
        x_t[28] = 21'b111111111110101000010;
        x_t[29] = 21'b000000000010111011111;
        x_t[30] = 21'b000000000000011001001;
        x_t[31] = 21'b000000000011001111110;
        x_t[32] = 21'b000000000010111100111;
        x_t[33] = 21'b000000000010000011000;
        x_t[34] = 21'b000000000001000001010;
        x_t[35] = 21'b000000000000001100111;
        x_t[36] = 21'b111111111111100101110;
        x_t[37] = 21'b111111111101110010010;
        x_t[38] = 21'b000000000011011000001;
        x_t[39] = 21'b000000000000011011101;
        x_t[40] = 21'b000000000001001001101;
        x_t[41] = 21'b000000000010100001111;
        x_t[42] = 21'b000000000101110011111;
        x_t[43] = 21'b000000000100000011111;
        x_t[44] = 21'b000000000010001111100;
        x_t[45] = 21'b000000000100101101011;
        x_t[46] = 21'b000000000100000101000;
        x_t[47] = 21'b000000000100010011011;
        x_t[48] = 21'b000000000011111010101;
        x_t[49] = 21'b000000000101001001010;
        x_t[50] = 21'b000000000100111100110;
        x_t[51] = 21'b000000000101001010110;
        x_t[52] = 21'b000000000101000100101;
        x_t[53] = 21'b000000000100000100001;
        x_t[54] = 21'b000000000100001100110;
        x_t[55] = 21'b000000000011011001011;
        x_t[56] = 21'b000000000100011100110;
        x_t[57] = 21'b000000000100111101100;
        x_t[58] = 21'b000000000100101000000;
        x_t[59] = 21'b000000000100001011101;
        x_t[60] = 21'b000000000011011101100;
        x_t[61] = 21'b000000000010010100011;
        x_t[62] = 21'b000000000011110011100;
        x_t[63] = 21'b000000000010011010010;
        
        h_t_prev[0] = 21'b000000000100101100001;
        h_t_prev[1] = 21'b000000000101011110000;
        h_t_prev[2] = 21'b000000000100011011010;
        h_t_prev[3] = 21'b000000000100011111101;
        h_t_prev[4] = 21'b000000000011010011010;
        h_t_prev[5] = 21'b000000000001110001111;
        h_t_prev[6] = 21'b000000000001100110101;
        h_t_prev[7] = 21'b000000000110100001111;
        h_t_prev[8] = 21'b000000000101101010101;
        h_t_prev[9] = 21'b000000000110001000110;
        h_t_prev[10] = 21'b000000000110000011001;
        h_t_prev[11] = 21'b000000000101010100101;
        h_t_prev[12] = 21'b000000000100010000100;
        h_t_prev[13] = 21'b000000000010001010011;
        h_t_prev[14] = 21'b000000000101010111010;
        h_t_prev[15] = 21'b000000000101100110101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 47 timeout!");
                $fdisplay(fd_cycles, "Test Vector  47: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  47: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 47");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 48
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000010101011111;
        x_t[1] = 21'b000000000011011110110;
        x_t[2] = 21'b000000000011001000110;
        x_t[3] = 21'b000000000011111101110;
        x_t[4] = 21'b000000000011000100001;
        x_t[5] = 21'b000000000001100001010;
        x_t[6] = 21'b000000000001111001010;
        x_t[7] = 21'b000000000010110111110;
        x_t[8] = 21'b000000000011111110011;
        x_t[9] = 21'b000000000100011111100;
        x_t[10] = 21'b000000000100101111111;
        x_t[11] = 21'b000000000100010010011;
        x_t[12] = 21'b000000000100000100110;
        x_t[13] = 21'b000000000010000011100;
        x_t[14] = 21'b000000000011101000100;
        x_t[15] = 21'b000000000100010000001;
        x_t[16] = 21'b000000000100100000111;
        x_t[17] = 21'b000000000100001001011;
        x_t[18] = 21'b000000000101011001100;
        x_t[19] = 21'b000000000101000011110;
        x_t[20] = 21'b000000000100010101001;
        x_t[21] = 21'b111111111111001110001;
        x_t[22] = 21'b111111111110010001000;
        x_t[23] = 21'b111111111110010110101;
        x_t[24] = 21'b111111111111100011100;
        x_t[25] = 21'b111111111111110011111;
        x_t[26] = 21'b111111111111111011010;
        x_t[27] = 21'b111111111111111101101;
        x_t[28] = 21'b111111111110100001111;
        x_t[29] = 21'b000000000010011010101;
        x_t[30] = 21'b111111111111110110000;
        x_t[31] = 21'b000000000011001011011;
        x_t[32] = 21'b000000000010000001110;
        x_t[33] = 21'b000000000001011001011;
        x_t[34] = 21'b000000000000110011000;
        x_t[35] = 21'b111111111111110100010;
        x_t[36] = 21'b111111111111111001101;
        x_t[37] = 21'b111111111110011111000;
        x_t[38] = 21'b000000000010111001111;
        x_t[39] = 21'b000000000001000000011;
        x_t[40] = 21'b000000000011100001110;
        x_t[41] = 21'b000000000011111100010;
        x_t[42] = 21'b000000000110000101110;
        x_t[43] = 21'b111111111110100100110;
        x_t[44] = 21'b000000000011010010100;
        x_t[45] = 21'b000000000100110101001;
        x_t[46] = 21'b000000000011010110011;
        x_t[47] = 21'b000000000100010011011;
        x_t[48] = 21'b000000000011110101110;
        x_t[49] = 21'b000000000101001101111;
        x_t[50] = 21'b000000000101001011001;
        x_t[51] = 21'b000000000101111011000;
        x_t[52] = 21'b000000000101101000011;
        x_t[53] = 21'b000000000100110110001;
        x_t[54] = 21'b000000000100111100101;
        x_t[55] = 21'b000000000011101010101;
        x_t[56] = 21'b000000000100111010111;
        x_t[57] = 21'b000000000101111101100;
        x_t[58] = 21'b000000000101111111001;
        x_t[59] = 21'b000000000101100110100;
        x_t[60] = 21'b000000000011110000101;
        x_t[61] = 21'b000000000011100111001;
        x_t[62] = 21'b000000000101010111011;
        x_t[63] = 21'b000000000100010101100;
        
        h_t_prev[0] = 21'b000000000010101011111;
        h_t_prev[1] = 21'b000000000011011110110;
        h_t_prev[2] = 21'b000000000011001000110;
        h_t_prev[3] = 21'b000000000011111101110;
        h_t_prev[4] = 21'b000000000011000100001;
        h_t_prev[5] = 21'b000000000001100001010;
        h_t_prev[6] = 21'b000000000001111001010;
        h_t_prev[7] = 21'b000000000010110111110;
        h_t_prev[8] = 21'b000000000011111110011;
        h_t_prev[9] = 21'b000000000100011111100;
        h_t_prev[10] = 21'b000000000100101111111;
        h_t_prev[11] = 21'b000000000100010010011;
        h_t_prev[12] = 21'b000000000100000100110;
        h_t_prev[13] = 21'b000000000010000011100;
        h_t_prev[14] = 21'b000000000011101000100;
        h_t_prev[15] = 21'b000000000100010000001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 48 timeout!");
                $fdisplay(fd_cycles, "Test Vector  48: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  48: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 48");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 49
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111100111010000;
        x_t[1] = 21'b111111111010111111100;
        x_t[2] = 21'b111111111000110100011;
        x_t[3] = 21'b111111110110111110010;
        x_t[4] = 21'b111111110111100010100;
        x_t[5] = 21'b111111110111000010000;
        x_t[6] = 21'b111111111000110000010;
        x_t[7] = 21'b111111111101110111001;
        x_t[8] = 21'b111111111000110001100;
        x_t[9] = 21'b111111111000001100110;
        x_t[10] = 21'b111111110111100110011;
        x_t[11] = 21'b111111110110101010111;
        x_t[12] = 21'b111111111000000000001;
        x_t[13] = 21'b111111110110111000000;
        x_t[14] = 21'b111111111010001111011;
        x_t[15] = 21'b111111111001100001101;
        x_t[16] = 21'b111111111000100000101;
        x_t[17] = 21'b111111110111111101110;
        x_t[18] = 21'b111111111001010111111;
        x_t[19] = 21'b111111111001110100010;
        x_t[20] = 21'b111111111001011000010;
        x_t[21] = 21'b111111111101010100100;
        x_t[22] = 21'b111111111011001111011;
        x_t[23] = 21'b111111111011001011101;
        x_t[24] = 21'b111111111111001000000;
        x_t[25] = 21'b111111111110111011111;
        x_t[26] = 21'b111111111000001101000;
        x_t[27] = 21'b111111110111110110111;
        x_t[28] = 21'b111111111010011100101;
        x_t[29] = 21'b111111111101101111001;
        x_t[30] = 21'b111111111100100111010;
        x_t[31] = 21'b111111110111100110101;
        x_t[32] = 21'b111111111000001010010;
        x_t[33] = 21'b111111110111001000100;
        x_t[34] = 21'b111111110110110000000;
        x_t[35] = 21'b111111111000000001111;
        x_t[36] = 21'b111111110111010010000;
        x_t[37] = 21'b111111111101000001010;
        x_t[38] = 21'b111111111011101111000;
        x_t[39] = 21'b111111110110101011000;
        x_t[40] = 21'b111111111001101011011;
        x_t[41] = 21'b111111110110110010110;
        x_t[42] = 21'b111111111010101100011;
        x_t[43] = 21'b111111111100010110001;
        x_t[44] = 21'b111111111011010000101;
        x_t[45] = 21'b111111111100000111111;
        x_t[46] = 21'b111111111011000101111;
        x_t[47] = 21'b111111111010101010101;
        x_t[48] = 21'b111111111010001111001;
        x_t[49] = 21'b111111111001111011001;
        x_t[50] = 21'b111111111001000100101;
        x_t[51] = 21'b111111111011010010000;
        x_t[52] = 21'b111111111100000010100;
        x_t[53] = 21'b111111111101010001111;
        x_t[54] = 21'b111111111011111101011;
        x_t[55] = 21'b111111111110011110011;
        x_t[56] = 21'b111111111100010000101;
        x_t[57] = 21'b111111111100101000101;
        x_t[58] = 21'b111111111110010010010;
        x_t[59] = 21'b111111111110011100101;
        x_t[60] = 21'b000000000000110100111;
        x_t[61] = 21'b111111111110110000110;
        x_t[62] = 21'b000000000000011101000;
        x_t[63] = 21'b000000000001001011001;
        
        h_t_prev[0] = 21'b111111111100111010000;
        h_t_prev[1] = 21'b111111111010111111100;
        h_t_prev[2] = 21'b111111111000110100011;
        h_t_prev[3] = 21'b111111110110111110010;
        h_t_prev[4] = 21'b111111110111100010100;
        h_t_prev[5] = 21'b111111110111000010000;
        h_t_prev[6] = 21'b111111111000110000010;
        h_t_prev[7] = 21'b111111111101110111001;
        h_t_prev[8] = 21'b111111111000110001100;
        h_t_prev[9] = 21'b111111111000001100110;
        h_t_prev[10] = 21'b111111110111100110011;
        h_t_prev[11] = 21'b111111110110101010111;
        h_t_prev[12] = 21'b111111111000000000001;
        h_t_prev[13] = 21'b111111110110111000000;
        h_t_prev[14] = 21'b111111111010001111011;
        h_t_prev[15] = 21'b111111111001100001101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 49 timeout!");
                $fdisplay(fd_cycles, "Test Vector  49: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  49: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 49");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 50
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111010111001110;
        x_t[1] = 21'b111111111001001111000;
        x_t[2] = 21'b111111110110100111100;
        x_t[3] = 21'b111111110100100011101;
        x_t[4] = 21'b111111110100011101100;
        x_t[5] = 21'b111111110011011110101;
        x_t[6] = 21'b111111110110010100101;
        x_t[7] = 21'b111111111011111101000;
        x_t[8] = 21'b111111110111001010011;
        x_t[9] = 21'b111111110110011110100;
        x_t[10] = 21'b111111110101110001000;
        x_t[11] = 21'b111111110101000101000;
        x_t[12] = 21'b111111110101000100111;
        x_t[13] = 21'b111111110101011000101;
        x_t[14] = 21'b111111111001001010111;
        x_t[15] = 21'b111111111000000110001;
        x_t[16] = 21'b111111110111001100011;
        x_t[17] = 21'b111111110110110011101;
        x_t[18] = 21'b111111110111101110100;
        x_t[19] = 21'b111111110111110110000;
        x_t[20] = 21'b111111110111101101111;
        x_t[21] = 21'b111111111100110000101;
        x_t[22] = 21'b111111111010110110000;
        x_t[23] = 21'b111111111010111010010;
        x_t[24] = 21'b111111111110111011111;
        x_t[25] = 21'b111111111110101111100;
        x_t[26] = 21'b111111110111000101001;
        x_t[27] = 21'b111111110110111000000;
        x_t[28] = 21'b111111111010001100111;
        x_t[29] = 21'b111111111101110011011;
        x_t[30] = 21'b111111111100011111011;
        x_t[31] = 21'b111111110110010110110;
        x_t[32] = 21'b111111110111000001101;
        x_t[33] = 21'b111111110101110000101;
        x_t[34] = 21'b111111110101010101100;
        x_t[35] = 21'b111111110110101001000;
        x_t[36] = 21'b111111110110000010100;
        x_t[37] = 21'b111111111100100100110;
        x_t[38] = 21'b111111111011111110001;
        x_t[39] = 21'b111111110110000110010;
        x_t[40] = 21'b111111111010001100000;
        x_t[41] = 21'b111111110100111100101;
        x_t[42] = 21'b111111111101110000001;
        x_t[43] = 21'b111111111000011001110;
        x_t[44] = 21'b111111111100011110111;
        x_t[45] = 21'b111111111011101001000;
        x_t[46] = 21'b111111111100001110100;
        x_t[47] = 21'b111111111011001000100;
        x_t[48] = 21'b111111111010100111000;
        x_t[49] = 21'b111111111010101001011;
        x_t[50] = 21'b111111111001111000111;
        x_t[51] = 21'b111111111011111000110;
        x_t[52] = 21'b111111111100001100110;
        x_t[53] = 21'b111111111101010001111;
        x_t[54] = 21'b111111111100011011010;
        x_t[55] = 21'b111111111110111000010;
        x_t[56] = 21'b111111111100101110101;
        x_t[57] = 21'b111111111101111101111;
        x_t[58] = 21'b111111111110011011000;
        x_t[59] = 21'b111111111110010000110;
        x_t[60] = 21'b111111111111100000100;
        x_t[61] = 21'b111111111101111011000;
        x_t[62] = 21'b111111111111000100010;
        x_t[63] = 21'b111111111110011011000;
        
        h_t_prev[0] = 21'b111111111010111001110;
        h_t_prev[1] = 21'b111111111001001111000;
        h_t_prev[2] = 21'b111111110110100111100;
        h_t_prev[3] = 21'b111111110100100011101;
        h_t_prev[4] = 21'b111111110100011101100;
        h_t_prev[5] = 21'b111111110011011110101;
        h_t_prev[6] = 21'b111111110110010100101;
        h_t_prev[7] = 21'b111111111011111101000;
        h_t_prev[8] = 21'b111111110111001010011;
        h_t_prev[9] = 21'b111111110110011110100;
        h_t_prev[10] = 21'b111111110101110001000;
        h_t_prev[11] = 21'b111111110101000101000;
        h_t_prev[12] = 21'b111111110101000100111;
        h_t_prev[13] = 21'b111111110101011000101;
        h_t_prev[14] = 21'b111111111001001010111;
        h_t_prev[15] = 21'b111111111000000110001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 50 timeout!");
                $fdisplay(fd_cycles, "Test Vector  50: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  50: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 50");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 51
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111011001000100;
        x_t[1] = 21'b111111111001000101001;
        x_t[2] = 21'b111111110111001001100;
        x_t[3] = 21'b111111110101001111001;
        x_t[4] = 21'b111111110101001010111;
        x_t[5] = 21'b111111110100110001111;
        x_t[6] = 21'b111111110111010010111;
        x_t[7] = 21'b111111111100100101110;
        x_t[8] = 21'b111111111000011100111;
        x_t[9] = 21'b111111110111111000101;
        x_t[10] = 21'b111111110111011100101;
        x_t[11] = 21'b111111110110110101001;
        x_t[12] = 21'b111111110101111111011;
        x_t[13] = 21'b111111110110001111001;
        x_t[14] = 21'b111111111010111110111;
        x_t[15] = 21'b111111111001111011001;
        x_t[16] = 21'b111111111001001101010;
        x_t[17] = 21'b111111111000101111000;
        x_t[18] = 21'b111111111001100010100;
        x_t[19] = 21'b111111111001011000111;
        x_t[20] = 21'b111111111000100110010;
        x_t[21] = 21'b111111111101001111000;
        x_t[22] = 21'b111111111011010101110;
        x_t[23] = 21'b111111111011011010001;
        x_t[24] = 21'b111111111111100011100;
        x_t[25] = 21'b111111111111011011000;
        x_t[26] = 21'b111111111000001101000;
        x_t[27] = 21'b111111110111110110111;
        x_t[28] = 21'b111111111010101001001;
        x_t[29] = 21'b111111111110101101101;
        x_t[30] = 21'b111111111101100101101;
        x_t[31] = 21'b111111111000001010001;
        x_t[32] = 21'b111111111000100001000;
        x_t[33] = 21'b111111110111001000100;
        x_t[34] = 21'b111111110110111110010;
        x_t[35] = 21'b111111111000010101101;
        x_t[36] = 21'b111111110111100101111;
        x_t[37] = 21'b111111111110010110111;
        x_t[38] = 21'b111111111110010101011;
        x_t[39] = 21'b111111111000110110101;
        x_t[40] = 21'b111111111110110110111;
        x_t[41] = 21'b111111111000000110010;
        x_t[42] = 21'b111111111110101011011;
        x_t[43] = 21'b111111111001100110101;
        x_t[44] = 21'b111111111110111011010;
        x_t[45] = 21'b111111111110100010110;
        x_t[46] = 21'b111111111110010000000;
        x_t[47] = 21'b111111111101010011110;
        x_t[48] = 21'b111111111100110101111;
        x_t[49] = 21'b111111111101010000010;
        x_t[50] = 21'b111111111100110110111;
        x_t[51] = 21'b111111111110001110011;
        x_t[52] = 21'b111111111110010001110;
        x_t[53] = 21'b111111111110111011101;
        x_t[54] = 21'b111111111110010011001;
        x_t[55] = 21'b111111111111001101110;
        x_t[56] = 21'b111111111101101111001;
        x_t[57] = 21'b000000000000000010000;
        x_t[58] = 21'b111111111111100101001;
        x_t[59] = 21'b111111111110100100100;
        x_t[60] = 21'b111111111111000001110;
        x_t[61] = 21'b111111111110000111011;
        x_t[62] = 21'b111111111111001011101;
        x_t[63] = 21'b111111111101110111111;
        
        h_t_prev[0] = 21'b111111111011001000100;
        h_t_prev[1] = 21'b111111111001000101001;
        h_t_prev[2] = 21'b111111110111001001100;
        h_t_prev[3] = 21'b111111110101001111001;
        h_t_prev[4] = 21'b111111110101001010111;
        h_t_prev[5] = 21'b111111110100110001111;
        h_t_prev[6] = 21'b111111110111010010111;
        h_t_prev[7] = 21'b111111111100100101110;
        h_t_prev[8] = 21'b111111111000011100111;
        h_t_prev[9] = 21'b111111110111111000101;
        h_t_prev[10] = 21'b111111110111011100101;
        h_t_prev[11] = 21'b111111110110110101001;
        h_t_prev[12] = 21'b111111110101111111011;
        h_t_prev[13] = 21'b111111110110001111001;
        h_t_prev[14] = 21'b111111111010111110111;
        h_t_prev[15] = 21'b111111111001111011001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 51 timeout!");
                $fdisplay(fd_cycles, "Test Vector  51: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  51: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 51");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 52
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111101101011010;
        x_t[1] = 21'b111111111100001000111;
        x_t[2] = 21'b111111111001111101001;
        x_t[3] = 21'b111111110111111101001;
        x_t[4] = 21'b111111111000000000110;
        x_t[5] = 21'b111111110111110100000;
        x_t[6] = 21'b111111111010110010111;
        x_t[7] = 21'b000000000000110011100;
        x_t[8] = 21'b111111111011110101100;
        x_t[9] = 21'b111111111011101110010;
        x_t[10] = 21'b111111111011010001010;
        x_t[11] = 21'b111111111001100010011;
        x_t[12] = 21'b111111111001011000000;
        x_t[13] = 21'b111111111001000111001;
        x_t[14] = 21'b111111111110110001011;
        x_t[15] = 21'b111111111101011010111;
        x_t[16] = 21'b111111111100100111011;
        x_t[17] = 21'b111111111100010111000;
        x_t[18] = 21'b111111111100100101100;
        x_t[19] = 21'b111111111100001110001;
        x_t[20] = 21'b111111111010110110001;
        x_t[21] = 21'b111111111110000011100;
        x_t[22] = 21'b111111111100001110111;
        x_t[23] = 21'b111111111100001000100;
        x_t[24] = 21'b000000000000011010010;
        x_t[25] = 21'b000000000000010010111;
        x_t[26] = 21'b111111111001010000100;
        x_t[27] = 21'b111111111000111101101;
        x_t[28] = 21'b111111111011011011100;
        x_t[29] = 21'b111111111111111000100;
        x_t[30] = 21'b111111111110101000000;
        x_t[31] = 21'b111111111001010101100;
        x_t[32] = 21'b111111111010010111001;
        x_t[33] = 21'b111111111001000000110;
        x_t[34] = 21'b111111111000101011110;
        x_t[35] = 21'b111111111010000111001;
        x_t[36] = 21'b111111111001110001000;
        x_t[37] = 21'b111111111111101100100;
        x_t[38] = 21'b000000000000001110100;
        x_t[39] = 21'b111111111010101100001;
        x_t[40] = 21'b111111111111000001110;
        x_t[41] = 21'b111111111100000000101;
        x_t[42] = 21'b111111111110110111010;
        x_t[43] = 21'b111111111111111100100;
        x_t[44] = 21'b111111111111101101100;
        x_t[45] = 21'b111111111111000001101;
        x_t[46] = 21'b111111111101101011110;
        x_t[47] = 21'b111111111101110001101;
        x_t[48] = 21'b111111111101100101101;
        x_t[49] = 21'b111111111110000011001;
        x_t[50] = 21'b111111111110011010110;
        x_t[51] = 21'b111111111111000011100;
        x_t[52] = 21'b111111111110110101101;
        x_t[53] = 21'b111111111111000001001;
        x_t[54] = 21'b111111111101111011010;
        x_t[55] = 21'b111111111110100010101;
        x_t[56] = 21'b111111111101010101011;
        x_t[57] = 21'b000000000000001010101;
        x_t[58] = 21'b111111111111001011000;
        x_t[59] = 21'b111111111101010001101;
        x_t[60] = 21'b111111111110101010110;
        x_t[61] = 21'b111111111110001011100;
        x_t[62] = 21'b111111111111011010011;
        x_t[63] = 21'b111111111101101111000;
        
        h_t_prev[0] = 21'b111111111101101011010;
        h_t_prev[1] = 21'b111111111100001000111;
        h_t_prev[2] = 21'b111111111001111101001;
        h_t_prev[3] = 21'b111111110111111101001;
        h_t_prev[4] = 21'b111111111000000000110;
        h_t_prev[5] = 21'b111111110111110100000;
        h_t_prev[6] = 21'b111111111010110010111;
        h_t_prev[7] = 21'b000000000000110011100;
        h_t_prev[8] = 21'b111111111011110101100;
        h_t_prev[9] = 21'b111111111011101110010;
        h_t_prev[10] = 21'b111111111011010001010;
        h_t_prev[11] = 21'b111111111001100010011;
        h_t_prev[12] = 21'b111111111001011000000;
        h_t_prev[13] = 21'b111111111001000111001;
        h_t_prev[14] = 21'b111111111110110001011;
        h_t_prev[15] = 21'b111111111101011010111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 52 timeout!");
                $fdisplay(fd_cycles, "Test Vector  52: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  52: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 52");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 53
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111111101011100;
        x_t[1] = 21'b111111111110000011010;
        x_t[2] = 21'b111111111100001010000;
        x_t[3] = 21'b111111111010110000000;
        x_t[4] = 21'b111111111010101100100;
        x_t[5] = 21'b111111111010001111010;
        x_t[6] = 21'b111111111101001000010;
        x_t[7] = 21'b000000000001100110011;
        x_t[8] = 21'b111111111100110011011;
        x_t[9] = 21'b111111111101011100100;
        x_t[10] = 21'b111111111101011111001;
        x_t[11] = 21'b111111111011010111101;
        x_t[12] = 21'b111111111011100100100;
        x_t[13] = 21'b111111111011001000101;
        x_t[14] = 21'b111111111101110010001;
        x_t[15] = 21'b111111111101100101000;
        x_t[16] = 21'b111111111101100111110;
        x_t[17] = 21'b111111111101011100001;
        x_t[18] = 21'b111111111101101010000;
        x_t[19] = 21'b111111111101001010100;
        x_t[20] = 21'b111111111011110100110;
        x_t[21] = 21'b111111111110011111001;
        x_t[22] = 21'b111111111100111110100;
        x_t[23] = 21'b111111111101000101011;
        x_t[24] = 21'b000000000000101111101;
        x_t[25] = 21'b000000000000101011110;
        x_t[26] = 21'b111111111010011100101;
        x_t[27] = 21'b111111111010011000000;
        x_t[28] = 21'b111111111100101010010;
        x_t[29] = 21'b000000000000001101010;
        x_t[30] = 21'b111111111111101110010;
        x_t[31] = 21'b111111111011000100011;
        x_t[32] = 21'b111111111011011111110;
        x_t[33] = 21'b111111111010011101010;
        x_t[34] = 21'b111111111010001011000;
        x_t[35] = 21'b111111111011011111111;
        x_t[36] = 21'b111111111011011110011;
        x_t[37] = 21'b000000000000110101111;
        x_t[38] = 21'b000000000000000100011;
        x_t[39] = 21'b111111111100000100011;
        x_t[40] = 21'b111111111110011011110;
        x_t[41] = 21'b111111111011101011110;
        x_t[42] = 21'b000000000001110101000;
        x_t[43] = 21'b111111111111011011101;
        x_t[44] = 21'b000000000000100101011;
        x_t[45] = 21'b111111111101110100010;
        x_t[46] = 21'b111111111101100110100;
        x_t[47] = 21'b111111111101001110110;
        x_t[48] = 21'b111111111101001001000;
        x_t[49] = 21'b111111111101110000101;
        x_t[50] = 21'b111111111110011010110;
        x_t[51] = 21'b111111111110110000010;
        x_t[52] = 21'b111111111110010110111;
        x_t[53] = 21'b111111111110010100101;
        x_t[54] = 21'b111111111100000011011;
        x_t[55] = 21'b111111111101011101101;
        x_t[56] = 21'b111111111100010100111;
        x_t[57] = 21'b111111111111010011001;
        x_t[58] = 21'b111111111101100110101;
        x_t[59] = 21'b111111111011101110111;
        x_t[60] = 21'b111111111101101001101;
        x_t[61] = 21'b111111111101000101001;
        x_t[62] = 21'b111111111110000101011;
        x_t[63] = 21'b111111111100110101111;
        
        h_t_prev[0] = 21'b111111111111101011100;
        h_t_prev[1] = 21'b111111111110000011010;
        h_t_prev[2] = 21'b111111111100001010000;
        h_t_prev[3] = 21'b111111111010110000000;
        h_t_prev[4] = 21'b111111111010101100100;
        h_t_prev[5] = 21'b111111111010001111010;
        h_t_prev[6] = 21'b111111111101001000010;
        h_t_prev[7] = 21'b000000000001100110011;
        h_t_prev[8] = 21'b111111111100110011011;
        h_t_prev[9] = 21'b111111111101011100100;
        h_t_prev[10] = 21'b111111111101011111001;
        h_t_prev[11] = 21'b111111111011010111101;
        h_t_prev[12] = 21'b111111111011100100100;
        h_t_prev[13] = 21'b111111111011001000101;
        h_t_prev[14] = 21'b111111111101110010001;
        h_t_prev[15] = 21'b111111111101100101000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 53 timeout!");
                $fdisplay(fd_cycles, "Test Vector  53: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  53: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 53");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 54
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111111010111110;
        x_t[1] = 21'b111111111101111001100;
        x_t[2] = 21'b111111111100010011110;
        x_t[3] = 21'b111111111011001101000;
        x_t[4] = 21'b111111111011000101110;
        x_t[5] = 21'b111111111010011111111;
        x_t[6] = 21'b111111111100101111011;
        x_t[7] = 21'b000000000000111101101;
        x_t[8] = 21'b111111111100011110110;
        x_t[9] = 21'b111111111100111110011;
        x_t[10] = 21'b111111111100110011001;
        x_t[11] = 21'b111111111010101110111;
        x_t[12] = 21'b111111111011011000110;
        x_t[13] = 21'b111111111011100011111;
        x_t[14] = 21'b111111111101100111101;
        x_t[15] = 21'b111111111101000110100;
        x_t[16] = 21'b111111111101000101001;
        x_t[17] = 21'b111111111100100101110;
        x_t[18] = 21'b111111111100101010110;
        x_t[19] = 21'b111111111100001000101;
        x_t[20] = 21'b111111111010111100011;
        x_t[21] = 21'b111111111110100100101;
        x_t[22] = 21'b111111111101001000000;
        x_t[23] = 21'b111111111101011100101;
        x_t[24] = 21'b000000000000110010101;
        x_t[25] = 21'b000000000000101011110;
        x_t[26] = 21'b111111111010100000110;
        x_t[27] = 21'b111111111010110111100;
        x_t[28] = 21'b111111111101000011100;
        x_t[29] = 21'b000000000000011001110;
        x_t[30] = 21'b111111111111110110000;
        x_t[31] = 21'b111111111011010001110;
        x_t[32] = 21'b111111111011011011010;
        x_t[33] = 21'b111111111010001111011;
        x_t[34] = 21'b111111111010001011000;
        x_t[35] = 21'b111111111011101001110;
        x_t[36] = 21'b111111111011011110011;
        x_t[37] = 21'b000000000001100110110;
        x_t[38] = 21'b111111111111110101010;
        x_t[39] = 21'b111111111100010011001;
        x_t[40] = 21'b000000000001011001111;
        x_t[41] = 21'b111111111011000010000;
        x_t[42] = 21'b000000000001001011100;
        x_t[43] = 21'b111111111001011011101;
        x_t[44] = 21'b000000000010100000010;
        x_t[45] = 21'b111111111011001010000;
        x_t[46] = 21'b111111111110001010110;
        x_t[47] = 21'b111111111101011000110;
        x_t[48] = 21'b111111111100111010110;
        x_t[49] = 21'b111111111100111101101;
        x_t[50] = 21'b111111111100110110111;
        x_t[51] = 21'b111111111100100100001;
        x_t[52] = 21'b111111111100000111101;
        x_t[53] = 21'b111111111100000011111;
        x_t[54] = 21'b111111111010000101100;
        x_t[55] = 21'b111111111100101110001;
        x_t[56] = 21'b111111111011100101101;
        x_t[57] = 21'b111111111101101100111;
        x_t[58] = 21'b111111111010111100100;
        x_t[59] = 21'b111111111001110100100;
        x_t[60] = 21'b111111111100010001100;
        x_t[61] = 21'b111111111011001101001;
        x_t[62] = 21'b111111111011010111100;
        x_t[63] = 21'b111111111011110011111;
        
        h_t_prev[0] = 21'b111111111111010111110;
        h_t_prev[1] = 21'b111111111101111001100;
        h_t_prev[2] = 21'b111111111100010011110;
        h_t_prev[3] = 21'b111111111011001101000;
        h_t_prev[4] = 21'b111111111011000101110;
        h_t_prev[5] = 21'b111111111010011111111;
        h_t_prev[6] = 21'b111111111100101111011;
        h_t_prev[7] = 21'b000000000000111101101;
        h_t_prev[8] = 21'b111111111100011110110;
        h_t_prev[9] = 21'b111111111100111110011;
        h_t_prev[10] = 21'b111111111100110011001;
        h_t_prev[11] = 21'b111111111010101110111;
        h_t_prev[12] = 21'b111111111011011000110;
        h_t_prev[13] = 21'b111111111011100011111;
        h_t_prev[14] = 21'b111111111101100111101;
        h_t_prev[15] = 21'b111111111101000110100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 54 timeout!");
                $fdisplay(fd_cycles, "Test Vector  54: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  54: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 54");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 55
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111111001110000;
        x_t[1] = 21'b111111111101100001000;
        x_t[2] = 21'b111111111011011110010;
        x_t[3] = 21'b111111111010000100100;
        x_t[4] = 21'b111111111010000100001;
        x_t[5] = 21'b111111111001101000100;
        x_t[6] = 21'b111111111011101011000;
        x_t[7] = 21'b000000000000111000100;
        x_t[8] = 21'b111111111100101110001;
        x_t[9] = 21'b111111111100001100010;
        x_t[10] = 21'b111111111011011111111;
        x_t[11] = 21'b111111111001010011001;
        x_t[12] = 21'b111111111010011110010;
        x_t[13] = 21'b111111111001111101101;
        x_t[14] = 21'b111111111111000001010;
        x_t[15] = 21'b111111111101000001011;
        x_t[16] = 21'b111111111100010011100;
        x_t[17] = 21'b111111111011001101000;
        x_t[18] = 21'b111111111011011011110;
        x_t[19] = 21'b111111111010111011110;
        x_t[20] = 21'b111111111001110111101;
        x_t[21] = 21'b111111111110011111001;
        x_t[22] = 21'b111111111100111000001;
        x_t[23] = 21'b111111111100110100000;
        x_t[24] = 21'b000000000000101111101;
        x_t[25] = 21'b000000000000101011110;
        x_t[26] = 21'b111111111001111111000;
        x_t[27] = 21'b111111111010001000010;
        x_t[28] = 21'b111111111100011010100;
        x_t[29] = 21'b000000000000100010000;
        x_t[30] = 21'b111111111111010010111;
        x_t[31] = 21'b111111111010010011101;
        x_t[32] = 21'b111111111010110110111;
        x_t[33] = 21'b111111111001011100100;
        x_t[34] = 21'b111111111001010001111;
        x_t[35] = 21'b111111111010111000011;
        x_t[36] = 21'b111111111010000100111;
        x_t[37] = 21'b000000000000001001000;
        x_t[38] = 21'b000000000001001011000;
        x_t[39] = 21'b111111111001110001011;
        x_t[40] = 21'b000000000010110000111;
        x_t[41] = 21'b111111110100101110101;
        x_t[42] = 21'b000000000010000110110;
        x_t[43] = 21'b111111111110111010110;
        x_t[44] = 21'b000000000010010101001;
        x_t[45] = 21'b111111111100011111001;
        x_t[46] = 21'b111111111101110110000;
        x_t[47] = 21'b111111111101001001110;
        x_t[48] = 21'b111111111100011001011;
        x_t[49] = 21'b111111111011111100110;
        x_t[50] = 21'b111111111011100110001;
        x_t[51] = 21'b111111111010111110110;
        x_t[52] = 21'b111111111011000000000;
        x_t[53] = 21'b111111111011011100111;
        x_t[54] = 21'b111111111010111011011;
        x_t[55] = 21'b111111111100001111111;
        x_t[56] = 21'b111111111011010000001;
        x_t[57] = 21'b111111111100011011111;
        x_t[58] = 21'b111111111010000011111;
        x_t[59] = 21'b111111111001110100100;
        x_t[60] = 21'b111111111011000100110;
        x_t[61] = 21'b111111111001110110010;
        x_t[62] = 21'b111111111001000111010;
        x_t[63] = 21'b111111111011010000101;
        
        h_t_prev[0] = 21'b111111111111001110000;
        h_t_prev[1] = 21'b111111111101100001000;
        h_t_prev[2] = 21'b111111111011011110010;
        h_t_prev[3] = 21'b111111111010000100100;
        h_t_prev[4] = 21'b111111111010000100001;
        h_t_prev[5] = 21'b111111111001101000100;
        h_t_prev[6] = 21'b111111111011101011000;
        h_t_prev[7] = 21'b000000000000111000100;
        h_t_prev[8] = 21'b111111111100101110001;
        h_t_prev[9] = 21'b111111111100001100010;
        h_t_prev[10] = 21'b111111111011011111111;
        h_t_prev[11] = 21'b111111111001010011001;
        h_t_prev[12] = 21'b111111111010011110010;
        h_t_prev[13] = 21'b111111111001111101101;
        h_t_prev[14] = 21'b111111111111000001010;
        h_t_prev[15] = 21'b111111111101000001011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 55 timeout!");
                $fdisplay(fd_cycles, "Test Vector  55: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  55: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 55");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 56
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111110111010010;
        x_t[1] = 21'b111111111100110101000;
        x_t[2] = 21'b111111111010101101110;
        x_t[3] = 21'b111111111001101100011;
        x_t[4] = 21'b111111111001100101111;
        x_t[5] = 21'b111111111001001100110;
        x_t[6] = 21'b111111111010011010000;
        x_t[7] = 21'b000000000000000101101;
        x_t[8] = 21'b111111111011111111110;
        x_t[9] = 21'b111111111011011010001;
        x_t[10] = 21'b111111111011000010101;
        x_t[11] = 21'b111111111001001000111;
        x_t[12] = 21'b111111111010000001000;
        x_t[13] = 21'b111111111000000011000;
        x_t[14] = 21'b111111111110010001110;
        x_t[15] = 21'b111111111100011000110;
        x_t[16] = 21'b111111111011011101000;
        x_t[17] = 21'b111111111010100000100;
        x_t[18] = 21'b111111111010111100001;
        x_t[19] = 21'b111111111010100000010;
        x_t[20] = 21'b111111111001101011001;
        x_t[21] = 21'b111111111101111110000;
        x_t[22] = 21'b111111111100011011101;
        x_t[23] = 21'b111111111100010001010;
        x_t[24] = 21'b000000000000100000011;
        x_t[25] = 21'b000000000000011100010;
        x_t[26] = 21'b111111111001101110001;
        x_t[27] = 21'b111111111001101000111;
        x_t[28] = 21'b111111111100001010110;
        x_t[29] = 21'b000000000000100010000;
        x_t[30] = 21'b111111111111010110110;
        x_t[31] = 21'b111111111010001010110;
        x_t[32] = 21'b111111111010001001100;
        x_t[33] = 21'b111111111001000101011;
        x_t[34] = 21'b111111111000111010001;
        x_t[35] = 21'b111111111010011010110;
        x_t[36] = 21'b111111111001110001000;
        x_t[37] = 21'b111111111111010000000;
        x_t[38] = 21'b000000000000001001011;
        x_t[39] = 21'b111111111001011011011;
        x_t[40] = 21'b000000000001000100010;
        x_t[41] = 21'b111111111000100010001;
        x_t[42] = 21'b000000000001100011001;
        x_t[43] = 21'b111111111110100100110;
        x_t[44] = 21'b000000000000101011000;
        x_t[45] = 21'b111111111110010011010;
        x_t[46] = 21'b111111111110100100101;
        x_t[47] = 21'b111111111101001110110;
        x_t[48] = 21'b111111111100001111110;
        x_t[49] = 21'b111111111011110011100;
        x_t[50] = 21'b111111111011100001011;
        x_t[51] = 21'b111111111011011011110;
        x_t[52] = 21'b111111111011111000011;
        x_t[53] = 21'b111111111100110110000;
        x_t[54] = 21'b111111111101000101010;
        x_t[55] = 21'b111111111100011000100;
        x_t[56] = 21'b111111111011100001010;
        x_t[57] = 21'b111111111100101100111;
        x_t[58] = 21'b111111111100000110110;
        x_t[59] = 21'b111111111100101110000;
        x_t[60] = 21'b111111111010110101100;
        x_t[61] = 21'b111111111010001010111;
        x_t[62] = 21'b111111111001011001110;
        x_t[63] = 21'b111111111100011011011;
        
        h_t_prev[0] = 21'b111111111110111010010;
        h_t_prev[1] = 21'b111111111100110101000;
        h_t_prev[2] = 21'b111111111010101101110;
        h_t_prev[3] = 21'b111111111001101100011;
        h_t_prev[4] = 21'b111111111001100101111;
        h_t_prev[5] = 21'b111111111001001100110;
        h_t_prev[6] = 21'b111111111010011010000;
        h_t_prev[7] = 21'b000000000000000101101;
        h_t_prev[8] = 21'b111111111011111111110;
        h_t_prev[9] = 21'b111111111011011010001;
        h_t_prev[10] = 21'b111111111011000010101;
        h_t_prev[11] = 21'b111111111001001000111;
        h_t_prev[12] = 21'b111111111010000001000;
        h_t_prev[13] = 21'b111111111000000011000;
        h_t_prev[14] = 21'b111111111110010001110;
        h_t_prev[15] = 21'b111111111100011000110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 56 timeout!");
                $fdisplay(fd_cycles, "Test Vector  56: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  56: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 56");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 57
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111110110000011;
        x_t[1] = 21'b111111111011111010010;
        x_t[2] = 21'b111111111001111101001;
        x_t[3] = 21'b111111111000110111001;
        x_t[4] = 21'b111111111001000010100;
        x_t[5] = 21'b111111111001010010010;
        x_t[6] = 21'b111111111011000101101;
        x_t[7] = 21'b000000000000000000100;
        x_t[8] = 21'b111111111011010001011;
        x_t[9] = 21'b111111111011000001001;
        x_t[10] = 21'b111111111010100101010;
        x_t[11] = 21'b111111111001001000111;
        x_t[12] = 21'b111111111010010010100;
        x_t[13] = 21'b111111111001100010011;
        x_t[14] = 21'b111111111110000111010;
        x_t[15] = 21'b111111111100100010111;
        x_t[16] = 21'b111111111011100001111;
        x_t[17] = 21'b111111111010100101100;
        x_t[18] = 21'b111111111011011011110;
        x_t[19] = 21'b111111111011000110101;
        x_t[20] = 21'b111111111010010110111;
        x_t[21] = 21'b111111111101100010011;
        x_t[22] = 21'b111111111100001000100;
        x_t[23] = 21'b111111111011111111111;
        x_t[24] = 21'b000000000000000100111;
        x_t[25] = 21'b000000000000000011011;
        x_t[26] = 21'b111111111001011101010;
        x_t[27] = 21'b111111111001011101000;
        x_t[28] = 21'b111111111011110111111;
        x_t[29] = 21'b000000000000010101100;
        x_t[30] = 21'b111111111110110011101;
        x_t[31] = 21'b111111111001110100100;
        x_t[32] = 21'b111111111001100101001;
        x_t[33] = 21'b111111111001000000110;
        x_t[34] = 21'b111111111000110101011;
        x_t[35] = 21'b111111111010010000111;
        x_t[36] = 21'b111111111010011000110;
        x_t[37] = 21'b111111111111001011111;
        x_t[38] = 21'b111111111111010111000;
        x_t[39] = 21'b111111111011001001101;
        x_t[40] = 21'b111111111111100111110;
        x_t[41] = 21'b111111111011111001101;
        x_t[42] = 21'b111111111110101011011;
        x_t[43] = 21'b111111111011101010010;
        x_t[44] = 21'b000000000000001111000;
        x_t[45] = 21'b111111111101000101111;
        x_t[46] = 21'b111111111110010101001;
        x_t[47] = 21'b111111111110000000100;
        x_t[48] = 21'b111111111100110101111;
        x_t[49] = 21'b111111111101000110111;
        x_t[50] = 21'b111111111100011010011;
        x_t[51] = 21'b111111111101011110001;
        x_t[52] = 21'b111111111101111101011;
        x_t[53] = 21'b111111111111010111011;
        x_t[54] = 21'b111111111111100001001;
        x_t[55] = 21'b111111111110000000001;
        x_t[56] = 21'b111111111101001100110;
        x_t[57] = 21'b111111111110100100010;
        x_t[58] = 21'b111111111111111011000;
        x_t[59] = 21'b000000000001100001111;
        x_t[60] = 21'b111111111100011101000;
        x_t[61] = 21'b111111111100110000100;
        x_t[62] = 21'b111111111101000110100;
        x_t[63] = 21'b111111111111000111000;
        
        h_t_prev[0] = 21'b111111111110110000011;
        h_t_prev[1] = 21'b111111111011111010010;
        h_t_prev[2] = 21'b111111111001111101001;
        h_t_prev[3] = 21'b111111111000110111001;
        h_t_prev[4] = 21'b111111111001000010100;
        h_t_prev[5] = 21'b111111111001010010010;
        h_t_prev[6] = 21'b111111111011000101101;
        h_t_prev[7] = 21'b000000000000000000100;
        h_t_prev[8] = 21'b111111111011010001011;
        h_t_prev[9] = 21'b111111111011000001001;
        h_t_prev[10] = 21'b111111111010100101010;
        h_t_prev[11] = 21'b111111111001001000111;
        h_t_prev[12] = 21'b111111111010010010100;
        h_t_prev[13] = 21'b111111111001100010011;
        h_t_prev[14] = 21'b111111111110000111010;
        h_t_prev[15] = 21'b111111111100100010111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 57 timeout!");
                $fdisplay(fd_cycles, "Test Vector  57: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  57: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 57");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 58
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111101110101001;
        x_t[1] = 21'b111111111011011000000;
        x_t[2] = 21'b111111111001100100111;
        x_t[3] = 21'b111111111000011010001;
        x_t[4] = 21'b111111111001000010100;
        x_t[5] = 21'b111111111001000111001;
        x_t[6] = 21'b111111111010111111011;
        x_t[7] = 21'b111111111111010111111;
        x_t[8] = 21'b111111111011001100010;
        x_t[9] = 21'b111111111011000001001;
        x_t[10] = 21'b111111111010111000110;
        x_t[11] = 21'b111111111001011000010;
        x_t[12] = 21'b111111111010101001111;
        x_t[13] = 21'b111111111001111101101;
        x_t[14] = 21'b111111111101111100101;
        x_t[15] = 21'b111111111100111100011;
        x_t[16] = 21'b111111111100001110100;
        x_t[17] = 21'b111111111010111001010;
        x_t[18] = 21'b111111111100010101110;
        x_t[19] = 21'b111111111100001000101;
        x_t[20] = 21'b111111111011001111001;
        x_t[21] = 21'b111111111101001100010;
        x_t[22] = 21'b111111111011011100001;
        x_t[23] = 21'b111111111011010100011;
        x_t[24] = 21'b111111111111011010010;
        x_t[25] = 21'b111111111111010111111;
        x_t[26] = 21'b111111111000101010100;
        x_t[27] = 21'b111111111000100110000;
        x_t[28] = 21'b111111111011001000101;
        x_t[29] = 21'b111111111110111010000;
        x_t[30] = 21'b111111111101110001011;
        x_t[31] = 21'b111111111000111010111;
        x_t[32] = 21'b111111111000111100010;
        x_t[33] = 21'b111111111000001101111;
        x_t[34] = 21'b111111111000001111010;
        x_t[35] = 21'b111111111001010101110;
        x_t[36] = 21'b111111111001001110010;
        x_t[37] = 21'b111111111101110010010;
        x_t[38] = 21'b111111111111001100111;
        x_t[39] = 21'b111111111001011011011;
        x_t[40] = 21'b111111111110011011110;
        x_t[41] = 21'b111111110110111001110;
        x_t[42] = 21'b111111111110111101001;
        x_t[43] = 21'b111111111101001101000;
        x_t[44] = 21'b000000000000001001100;
        x_t[45] = 21'b111111111111010001001;
        x_t[46] = 21'b111111111110010000000;
        x_t[47] = 21'b111111111110101000010;
        x_t[48] = 21'b111111111110000010001;
        x_t[49] = 21'b111111111110010001001;
        x_t[50] = 21'b111111111101001110101;
        x_t[51] = 21'b111111111111100101011;
        x_t[52] = 21'b000000000000010001101;
        x_t[53] = 21'b000000000010001111001;
        x_t[54] = 21'b000000000011001010110;
        x_t[55] = 21'b111111111111101100000;
        x_t[56] = 21'b111111111110111000001;
        x_t[57] = 21'b000000000000010111011;
        x_t[58] = 21'b000000000011111000000;
        x_t[59] = 21'b000000000110100001101;
        x_t[60] = 21'b111111111111000101101;
        x_t[61] = 21'b000000000000110101001;
        x_t[62] = 21'b000000000010111100000;
        x_t[63] = 21'b000000000010011110110;
        
        h_t_prev[0] = 21'b111111111101110101001;
        h_t_prev[1] = 21'b111111111011011000000;
        h_t_prev[2] = 21'b111111111001100100111;
        h_t_prev[3] = 21'b111111111000011010001;
        h_t_prev[4] = 21'b111111111001000010100;
        h_t_prev[5] = 21'b111111111001000111001;
        h_t_prev[6] = 21'b111111111010111111011;
        h_t_prev[7] = 21'b111111111111010111111;
        h_t_prev[8] = 21'b111111111011001100010;
        h_t_prev[9] = 21'b111111111011000001001;
        h_t_prev[10] = 21'b111111111010111000110;
        h_t_prev[11] = 21'b111111111001011000010;
        h_t_prev[12] = 21'b111111111010101001111;
        h_t_prev[13] = 21'b111111111001111101101;
        h_t_prev[14] = 21'b111111111101111100101;
        h_t_prev[15] = 21'b111111111100111100011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 58 timeout!");
                $fdisplay(fd_cycles, "Test Vector  58: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  58: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 58");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 59
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111101110000010;
        x_t[1] = 21'b111111111011111111001;
        x_t[2] = 21'b111111111001101001110;
        x_t[3] = 21'b111111111000010101010;
        x_t[4] = 21'b111111111000110011010;
        x_t[5] = 21'b111111111000101011100;
        x_t[6] = 21'b111111111001101000010;
        x_t[7] = 21'b111111111111010010110;
        x_t[8] = 21'b111111111011110101100;
        x_t[9] = 21'b111111111011010101001;
        x_t[10] = 21'b111111111011001100011;
        x_t[11] = 21'b111111111001110001101;
        x_t[12] = 21'b111111111010011000011;
        x_t[13] = 21'b111111111000100101001;
        x_t[14] = 21'b111111111110011100011;
        x_t[15] = 21'b111111111101011111111;
        x_t[16] = 21'b111111111100111011001;
        x_t[17] = 21'b111111111011010001111;
        x_t[18] = 21'b111111111100110101011;
        x_t[19] = 21'b111111111100110100100;
        x_t[20] = 21'b111111111100000001010;
        x_t[21] = 21'b111111111101111000100;
        x_t[22] = 21'b111111111100001000100;
        x_t[23] = 21'b111111111100000101101;
        x_t[24] = 21'b000000000000001011000;
        x_t[25] = 21'b000000000000000011011;
        x_t[26] = 21'b111111111001100101101;
        x_t[27] = 21'b111111111001011001001;
        x_t[28] = 21'b111111111011101000001;
        x_t[29] = 21'b111111111111111100101;
        x_t[30] = 21'b111111111110101011111;
        x_t[31] = 21'b111111111001111101011;
        x_t[32] = 21'b111111111010001001100;
        x_t[33] = 21'b111111111000110111100;
        x_t[34] = 21'b111111111000110000101;
        x_t[35] = 21'b111111111010001100000;
        x_t[36] = 21'b111111111001010011010;
        x_t[37] = 21'b111111111101011001110;
        x_t[38] = 21'b000000000000011101101;
        x_t[39] = 21'b111111111000101111010;
        x_t[40] = 21'b000000000000101001000;
        x_t[41] = 21'b111111110111000000110;
        x_t[42] = 21'b000000000010100100011;
        x_t[43] = 21'b111111111100001011001;
        x_t[44] = 21'b000000000010100101111;
        x_t[45] = 21'b000000000010000011001;
        x_t[46] = 21'b000000000000011011111;
        x_t[47] = 21'b000000000000001011110;
        x_t[48] = 21'b111111111111001001101;
        x_t[49] = 21'b111111111110100011101;
        x_t[50] = 21'b111111111101011000001;
        x_t[51] = 21'b000000000000001100000;
        x_t[52] = 21'b000000000001001111001;
        x_t[53] = 21'b000000000011101101110;
        x_t[54] = 21'b000000000101000010101;
        x_t[55] = 21'b000000000001111010100;
        x_t[56] = 21'b000000000000001110001;
        x_t[57] = 21'b000000000000011011101;
        x_t[58] = 21'b000000000101000110100;
        x_t[59] = 21'b000000001000011100000;
        x_t[60] = 21'b000000000001110010001;
        x_t[61] = 21'b000000000100000000000;
        x_t[62] = 21'b000000000111100111101;
        x_t[63] = 21'b000000000101000101111;
        
        h_t_prev[0] = 21'b111111111101110000010;
        h_t_prev[1] = 21'b111111111011111111001;
        h_t_prev[2] = 21'b111111111001101001110;
        h_t_prev[3] = 21'b111111111000010101010;
        h_t_prev[4] = 21'b111111111000110011010;
        h_t_prev[5] = 21'b111111111000101011100;
        h_t_prev[6] = 21'b111111111001101000010;
        h_t_prev[7] = 21'b111111111111010010110;
        h_t_prev[8] = 21'b111111111011110101100;
        h_t_prev[9] = 21'b111111111011010101001;
        h_t_prev[10] = 21'b111111111011001100011;
        h_t_prev[11] = 21'b111111111001110001101;
        h_t_prev[12] = 21'b111111111010011000011;
        h_t_prev[13] = 21'b111111111000100101001;
        h_t_prev[14] = 21'b111111111110011100011;
        h_t_prev[15] = 21'b111111111101011111111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 59 timeout!");
                $fdisplay(fd_cycles, "Test Vector  59: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  59: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 59");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 60
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111111101011100;
        x_t[1] = 21'b111111111101111110011;
        x_t[2] = 21'b111111111011001111110;
        x_t[3] = 21'b111111111001110110000;
        x_t[4] = 21'b111111111001011011110;
        x_t[5] = 21'b111111111001000111001;
        x_t[6] = 21'b111111111010010011111;
        x_t[7] = 21'b000000000001000010110;
        x_t[8] = 21'b111111111101001101001;
        x_t[9] = 21'b111111111100010001010;
        x_t[10] = 21'b111111111011111000011;
        x_t[11] = 21'b111111111010001011001;
        x_t[12] = 21'b111111111011000111001;
        x_t[13] = 21'b111111111001110110111;
        x_t[14] = 21'b000000000000000000100;
        x_t[15] = 21'b111111111110000011100;
        x_t[16] = 21'b111111111101000101001;
        x_t[17] = 21'b111111111011100101101;
        x_t[18] = 21'b111111111101000101001;
        x_t[19] = 21'b111111111101100000100;
        x_t[20] = 21'b111111111101010010101;
        x_t[21] = 21'b111111111110001011110;
        x_t[22] = 21'b111111111100000010010;
        x_t[23] = 21'b111111111011110100010;
        x_t[24] = 21'b000000000000011101010;
        x_t[25] = 21'b000000000000010010111;
        x_t[26] = 21'b111111111001111111000;
        x_t[27] = 21'b111111111001000001100;
        x_t[28] = 21'b111111111010111100000;
        x_t[29] = 21'b000000000000100110010;
        x_t[30] = 21'b111111111111010110110;
        x_t[31] = 21'b111111111001110000001;
        x_t[32] = 21'b111111111010110110111;
        x_t[33] = 21'b111111111001100001001;
        x_t[34] = 21'b111111111000110000101;
        x_t[35] = 21'b111111111010010000111;
        x_t[36] = 21'b111111111000100001100;
        x_t[37] = 21'b111111111101000001010;
        x_t[38] = 21'b000000000000110001110;
        x_t[39] = 21'b111111111000110110101;
        x_t[40] = 21'b000000000010010101110;
        x_t[41] = 21'b111111111001000100111;
        x_t[42] = 21'b000000000010001100101;
        x_t[43] = 21'b111111111011110101010;
        x_t[44] = 21'b000000000010110001000;
        x_t[45] = 21'b111111111111100000101;
        x_t[46] = 21'b000000000001001111101;
        x_t[47] = 21'b000000000000011010101;
        x_t[48] = 21'b111111111111000000001;
        x_t[49] = 21'b111111111110010001001;
        x_t[50] = 21'b111111111101000000011;
        x_t[51] = 21'b000000000000000111001;
        x_t[52] = 21'b000000000001011001010;
        x_t[53] = 21'b000000000011101101110;
        x_t[54] = 21'b000000000100101010101;
        x_t[55] = 21'b000000000010101001111;
        x_t[56] = 21'b000000000000100011100;
        x_t[57] = 21'b000000000000001110111;
        x_t[58] = 21'b000000000101010111111;
        x_t[59] = 21'b000000001000110111101;
        x_t[60] = 21'b000000000011011001101;
        x_t[61] = 21'b000000000100111001111;
        x_t[62] = 21'b000000001001001111010;
        x_t[63] = 21'b000000000101011011111;
        
        h_t_prev[0] = 21'b111111111111101011100;
        h_t_prev[1] = 21'b111111111101111110011;
        h_t_prev[2] = 21'b111111111011001111110;
        h_t_prev[3] = 21'b111111111001110110000;
        h_t_prev[4] = 21'b111111111001011011110;
        h_t_prev[5] = 21'b111111111001000111001;
        h_t_prev[6] = 21'b111111111010010011111;
        h_t_prev[7] = 21'b000000000001000010110;
        h_t_prev[8] = 21'b111111111101001101001;
        h_t_prev[9] = 21'b111111111100010001010;
        h_t_prev[10] = 21'b111111111011111000011;
        h_t_prev[11] = 21'b111111111010001011001;
        h_t_prev[12] = 21'b111111111011000111001;
        h_t_prev[13] = 21'b111111111001110110111;
        h_t_prev[14] = 21'b000000000000000000100;
        h_t_prev[15] = 21'b111111111110000011100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 60 timeout!");
                $fdisplay(fd_cycles, "Test Vector  60: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  60: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 60");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 61
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111111100110101;
        x_t[1] = 21'b111111111101010111010;
        x_t[2] = 21'b111111111010110111100;
        x_t[3] = 21'b111111111001001111011;
        x_t[4] = 21'b111111111000101001010;
        x_t[5] = 21'b111111111000001111110;
        x_t[6] = 21'b111111111001000010111;
        x_t[7] = 21'b000000000000110011100;
        x_t[8] = 21'b111111111100101110001;
        x_t[9] = 21'b111111111011111101010;
        x_t[10] = 21'b111111111011111000011;
        x_t[11] = 21'b111111111001100111100;
        x_t[12] = 21'b111111111010111011100;
        x_t[13] = 21'b111111111001111101101;
        x_t[14] = 21'b000000000000000101110;
        x_t[15] = 21'b111111111101101010001;
        x_t[16] = 21'b111111111101000000001;
        x_t[17] = 21'b111111111011111001011;
        x_t[18] = 21'b111111111101100100110;
        x_t[19] = 21'b111111111110000001011;
        x_t[20] = 21'b111111111101111110011;
        x_t[21] = 21'b111111111101000100000;
        x_t[22] = 21'b111111111010101100100;
        x_t[23] = 21'b111111111010100000001;
        x_t[24] = 21'b111111111111100110100;
        x_t[25] = 21'b111111111111011011000;
        x_t[26] = 21'b111111111000101010100;
        x_t[27] = 21'b111111110111010111011;
        x_t[28] = 21'b111111111001110000100;
        x_t[29] = 21'b000000000001001111110;
        x_t[30] = 21'b111111111110010000101;
        x_t[31] = 21'b111111111000111010111;
        x_t[32] = 21'b111111111001111011111;
        x_t[33] = 21'b111111111000011011110;
        x_t[34] = 21'b111111110111011010111;
        x_t[35] = 21'b111111111000110011001;
        x_t[36] = 21'b111111110111100000111;
        x_t[37] = 21'b111111111100110101000;
        x_t[38] = 21'b000000000001011111001;
        x_t[39] = 21'b111111110111111011110;
        x_t[40] = 21'b000000000010100110000;
        x_t[41] = 21'b111111111000110000000;
        x_t[42] = 21'b000000000001101111000;
        x_t[43] = 21'b000000000010000000001;
        x_t[44] = 21'b000000000011111111010;
        x_t[45] = 21'b000000000001110011101;
        x_t[46] = 21'b000000000011010110011;
        x_t[47] = 21'b000000000010010010000;
        x_t[48] = 21'b000000000000011111011;
        x_t[49] = 21'b111111111111110111000;
        x_t[50] = 21'b111111111110110010100;
        x_t[51] = 21'b000000000001110110010;
        x_t[52] = 21'b000000000010111111101;
        x_t[53] = 21'b000000000101011101001;
        x_t[54] = 21'b000000000110010110100;
        x_t[55] = 21'b000000000101000101010;
        x_t[56] = 21'b000000000010101101000;
        x_t[57] = 21'b000000000001110101001;
        x_t[58] = 21'b000000000110100110011;
        x_t[59] = 21'b000000001001010111010;
        x_t[60] = 21'b000000000100110001111;
        x_t[61] = 21'b000000000101000010001;
        x_t[62] = 21'b000000001001000100001;
        x_t[63] = 21'b000000000101101001001;
        
        h_t_prev[0] = 21'b111111111111100110101;
        h_t_prev[1] = 21'b111111111101010111010;
        h_t_prev[2] = 21'b111111111010110111100;
        h_t_prev[3] = 21'b111111111001001111011;
        h_t_prev[4] = 21'b111111111000101001010;
        h_t_prev[5] = 21'b111111111000001111110;
        h_t_prev[6] = 21'b111111111001000010111;
        h_t_prev[7] = 21'b000000000000110011100;
        h_t_prev[8] = 21'b111111111100101110001;
        h_t_prev[9] = 21'b111111111011111101010;
        h_t_prev[10] = 21'b111111111011111000011;
        h_t_prev[11] = 21'b111111111001100111100;
        h_t_prev[12] = 21'b111111111010111011100;
        h_t_prev[13] = 21'b111111111001111101101;
        h_t_prev[14] = 21'b000000000000000101110;
        h_t_prev[15] = 21'b111111111101101010001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 61 timeout!");
                $fdisplay(fd_cycles, "Test Vector  61: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  61: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 61");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 62
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000000100110110;
        x_t[1] = 21'b111111111110010010000;
        x_t[2] = 21'b111111111011011110010;
        x_t[3] = 21'b111111111000101101100;
        x_t[4] = 21'b111111111000011111001;
        x_t[5] = 21'b111111111000001111110;
        x_t[6] = 21'b111111111001110100110;
        x_t[7] = 21'b000000000010101000100;
        x_t[8] = 21'b111111111110011010100;
        x_t[9] = 21'b111111111101100110100;
        x_t[10] = 21'b111111111101010000100;
        x_t[11] = 21'b111111111010011111100;
        x_t[12] = 21'b111111111011011000110;
        x_t[13] = 21'b111111111011101010101;
        x_t[14] = 21'b000000000010011001100;
        x_t[15] = 21'b000000000000001100111;
        x_t[16] = 21'b111111111111001111111;
        x_t[17] = 21'b111111111101101111111;
        x_t[18] = 21'b111111111111001110001;
        x_t[19] = 21'b111111111111011110110;
        x_t[20] = 21'b111111111111101111000;
        x_t[21] = 21'b111111111101010111010;
        x_t[22] = 21'b111111111010111111101;
        x_t[23] = 21'b111111111011000000000;
        x_t[24] = 21'b111111111111111000110;
        x_t[25] = 21'b111111111111101010100;
        x_t[26] = 21'b111111111000101110110;
        x_t[27] = 21'b111111110111100011010;
        x_t[28] = 21'b111111111010011001011;
        x_t[29] = 21'b000000000001000111100;
        x_t[30] = 21'b111111111110101111110;
        x_t[31] = 21'b111111111000110110100;
        x_t[32] = 21'b111111111010010010101;
        x_t[33] = 21'b111111111000010010100;
        x_t[34] = 21'b111111110111010001010;
        x_t[35] = 21'b111111111000110011001;
        x_t[36] = 21'b111111110111111110110;
        x_t[37] = 21'b111111111101111110011;
        x_t[38] = 21'b000000000010000111100;
        x_t[39] = 21'b111111111001000101010;
        x_t[40] = 21'b000000000001111010100;
        x_t[41] = 21'b111111111001001011110;
        x_t[42] = 21'b000000000100100000111;
        x_t[43] = 21'b111111111110101111110;
        x_t[44] = 21'b000000000110110010000;
        x_t[45] = 21'b000000000011011000010;
        x_t[46] = 21'b000000000110101010110;
        x_t[47] = 21'b000000000100001110011;
        x_t[48] = 21'b000000000001111001111;
        x_t[49] = 21'b000000000001001111000;
        x_t[50] = 21'b111111111111110101000;
        x_t[51] = 21'b000000000010000100110;
        x_t[52] = 21'b000000000010110000010;
        x_t[53] = 21'b000000000101000001010;
        x_t[54] = 21'b000000000101110010101;
        x_t[55] = 21'b000000000111000010100;
        x_t[56] = 21'b000000000100001011101;
        x_t[57] = 21'b000000000010100100000;
        x_t[58] = 21'b000000000101110110100;
        x_t[59] = 21'b000000001000000100011;
        x_t[60] = 21'b000000000110010001101;
        x_t[61] = 21'b000000000101010110111;
        x_t[62] = 21'b000000001000011011011;
        x_t[63] = 21'b000000000110111100110;
        
        h_t_prev[0] = 21'b000000000000100110110;
        h_t_prev[1] = 21'b111111111110010010000;
        h_t_prev[2] = 21'b111111111011011110010;
        h_t_prev[3] = 21'b111111111000101101100;
        h_t_prev[4] = 21'b111111111000011111001;
        h_t_prev[5] = 21'b111111111000001111110;
        h_t_prev[6] = 21'b111111111001110100110;
        h_t_prev[7] = 21'b000000000010101000100;
        h_t_prev[8] = 21'b111111111110011010100;
        h_t_prev[9] = 21'b111111111101100110100;
        h_t_prev[10] = 21'b111111111101010000100;
        h_t_prev[11] = 21'b111111111010011111100;
        h_t_prev[12] = 21'b111111111011011000110;
        h_t_prev[13] = 21'b111111111011101010101;
        h_t_prev[14] = 21'b000000000010011001100;
        h_t_prev[15] = 21'b000000000000001100111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 62 timeout!");
                $fdisplay(fd_cycles, "Test Vector  62: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  62: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 62");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 63
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000000000100010;
        x_t[1] = 21'b111111111110110100010;
        x_t[2] = 21'b111111111100000101001;
        x_t[3] = 21'b111111111001010100001;
        x_t[4] = 21'b111111111000000101111;
        x_t[5] = 21'b111111110111001101001;
        x_t[6] = 21'b111111111001001111011;
        x_t[7] = 21'b000000000010100011011;
        x_t[8] = 21'b111111111110101010000;
        x_t[9] = 21'b111111111110010011101;
        x_t[10] = 21'b111111111101010101011;
        x_t[11] = 21'b111111111001100010011;
        x_t[12] = 21'b111111111001011000000;
        x_t[13] = 21'b111111111001111101101;
        x_t[14] = 21'b000000000011011110000;
        x_t[15] = 21'b000000000000101011011;
        x_t[16] = 21'b111111111111100011101;
        x_t[17] = 21'b111111111101111001110;
        x_t[18] = 21'b111111111110101001010;
        x_t[19] = 21'b111111111110000110111;
        x_t[20] = 21'b111111111101101011101;
        x_t[21] = 21'b111111111101111000100;
        x_t[22] = 21'b111111111011100010100;
        x_t[23] = 21'b111111111011011010001;
        x_t[24] = 21'b000000000000011101010;
        x_t[25] = 21'b000000000000001111110;
        x_t[26] = 21'b111111111001010000100;
        x_t[27] = 21'b111111110111101111000;
        x_t[28] = 21'b111111111001110110110;
        x_t[29] = 21'b000000000001110101010;
        x_t[30] = 21'b111111111111010010111;
        x_t[31] = 21'b111111111001010001000;
        x_t[32] = 21'b111111111011001001001;
        x_t[33] = 21'b111111111001001110101;
        x_t[34] = 21'b111111111000000000111;
        x_t[35] = 21'b111111111001010101110;
        x_t[36] = 21'b111111111000001000101;
        x_t[37] = 21'b111111111110000010100;
        x_t[38] = 21'b000000000010010001100;
        x_t[39] = 21'b111111111001010100000;
        x_t[40] = 21'b000000000011010110111;
        x_t[41] = 21'b111111111011011101111;
        x_t[42] = 21'b000000000101011100010;
        x_t[43] = 21'b111111111101011000000;
        x_t[44] = 21'b000000000110110010000;
        x_t[45] = 21'b000000000000100110010;
        x_t[46] = 21'b000000000110000001010;
        x_t[47] = 21'b000000000100001001011;
        x_t[48] = 21'b000000000001101011101;
        x_t[49] = 21'b000000000001001010011;
        x_t[50] = 21'b111111111111011000100;
        x_t[51] = 21'b000000000000110111100;
        x_t[52] = 21'b000000000001010100001;
        x_t[53] = 21'b000000000010110110001;
        x_t[54] = 21'b000000000011100010110;
        x_t[55] = 21'b000000000110110101100;
        x_t[56] = 21'b000000000011111110101;
        x_t[57] = 21'b000000000010000110010;
        x_t[58] = 21'b000000000011110011101;
        x_t[59] = 21'b000000000100010111100;
        x_t[60] = 21'b000000000110101100100;
        x_t[61] = 21'b000000000100010100101;
        x_t[62] = 21'b000000000110011101101;
        x_t[63] = 21'b000000000110011101111;
        
        h_t_prev[0] = 21'b000000000000000100010;
        h_t_prev[1] = 21'b111111111110110100010;
        h_t_prev[2] = 21'b111111111100000101001;
        h_t_prev[3] = 21'b111111111001010100001;
        h_t_prev[4] = 21'b111111111000000101111;
        h_t_prev[5] = 21'b111111110111001101001;
        h_t_prev[6] = 21'b111111111001001111011;
        h_t_prev[7] = 21'b000000000010100011011;
        h_t_prev[8] = 21'b111111111110101010000;
        h_t_prev[9] = 21'b111111111110010011101;
        h_t_prev[10] = 21'b111111111101010101011;
        h_t_prev[11] = 21'b111111111001100010011;
        h_t_prev[12] = 21'b111111111001011000000;
        h_t_prev[13] = 21'b111111111001111101101;
        h_t_prev[14] = 21'b000000000011011110000;
        h_t_prev[15] = 21'b000000000000101011011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 63 timeout!");
                $fdisplay(fd_cycles, "Test Vector  63: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  63: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 63");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 64
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000000111010100;
        x_t[1] = 21'b111111111111010110100;
        x_t[2] = 21'b111111111100011101011;
        x_t[3] = 21'b111111111001110110000;
        x_t[4] = 21'b111111111000111000011;
        x_t[5] = 21'b111111110111101000111;
        x_t[6] = 21'b111111111001011011110;
        x_t[7] = 21'b000000000010110111110;
        x_t[8] = 21'b111111111110101111001;
        x_t[9] = 21'b111111111110000100101;
        x_t[10] = 21'b111111111100101001011;
        x_t[11] = 21'b111111111001100010011;
        x_t[12] = 21'b111111111000110100111;
        x_t[13] = 21'b111111111001111101101;
        x_t[14] = 21'b000000000010111001001;
        x_t[15] = 21'b000000000000010111000;
        x_t[16] = 21'b111111111111001010111;
        x_t[17] = 21'b111111111101101010111;
        x_t[18] = 21'b111111111110000100011;
        x_t[19] = 21'b111111111101001010100;
        x_t[20] = 21'b111111111100100110110;
        x_t[21] = 21'b111111111110100100101;
        x_t[22] = 21'b111111111100011011101;
        x_t[23] = 21'b111111111100010111000;
        x_t[24] = 21'b000000000001000001111;
        x_t[25] = 21'b000000000000110101001;
        x_t[26] = 21'b111111111010000111100;
        x_t[27] = 21'b111111111000111001101;
        x_t[28] = 21'b111111111011100101000;
        x_t[29] = 21'b000000000010100011000;
        x_t[30] = 21'b111111111111011010110;
        x_t[31] = 21'b111111111010100000111;
        x_t[32] = 21'b111111111011001101101;
        x_t[33] = 21'b111111111001101010011;
        x_t[34] = 21'b111111111000110101011;
        x_t[35] = 21'b111111111010000010001;
        x_t[36] = 21'b111111111000111010011;
        x_t[37] = 21'b111111111110011111000;
        x_t[38] = 21'b000000000011000100000;
        x_t[39] = 21'b111111111010100100111;
        x_t[40] = 21'b000000000101001110100;
        x_t[41] = 21'b111111111101011011000;
        x_t[42] = 21'b000000000101101110000;
        x_t[43] = 21'b111111111100100001001;
        x_t[44] = 21'b000000000110101100011;
        x_t[45] = 21'b111111111111110000001;
        x_t[46] = 21'b000000000101001101100;
        x_t[47] = 21'b000000000011010111101;
        x_t[48] = 21'b000000000001010011110;
        x_t[49] = 21'b000000000001000001001;
        x_t[50] = 21'b111111111111101011100;
        x_t[51] = 21'b000000000000101001000;
        x_t[52] = 21'b000000000000110000011;
        x_t[53] = 21'b000000000001100010101;
        x_t[54] = 21'b000000000001100100111;
        x_t[55] = 21'b000000000110000001110;
        x_t[56] = 21'b000000000011011000000;
        x_t[57] = 21'b000000000010000010000;
        x_t[58] = 21'b000000000010101101110;
        x_t[59] = 21'b000000000010000101100;
        x_t[60] = 21'b000000000101110110111;
        x_t[61] = 21'b000000000010110001011;
        x_t[62] = 21'b000000000100010001001;
        x_t[63] = 21'b000000000101011011111;
        
        h_t_prev[0] = 21'b000000000000111010100;
        h_t_prev[1] = 21'b111111111111010110100;
        h_t_prev[2] = 21'b111111111100011101011;
        h_t_prev[3] = 21'b111111111001110110000;
        h_t_prev[4] = 21'b111111111000111000011;
        h_t_prev[5] = 21'b111111110111101000111;
        h_t_prev[6] = 21'b111111111001011011110;
        h_t_prev[7] = 21'b000000000010110111110;
        h_t_prev[8] = 21'b111111111110101111001;
        h_t_prev[9] = 21'b111111111110000100101;
        h_t_prev[10] = 21'b111111111100101001011;
        h_t_prev[11] = 21'b111111111001100010011;
        h_t_prev[12] = 21'b111111111000110100111;
        h_t_prev[13] = 21'b111111111001111101101;
        h_t_prev[14] = 21'b000000000010111001001;
        h_t_prev[15] = 21'b000000000000010111000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 64 timeout!");
                $fdisplay(fd_cycles, "Test Vector  64: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  64: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 64");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 65
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111001001101010;
        x_t[1] = 21'b111111111011110000100;
        x_t[2] = 21'b111111111100001010000;
        x_t[3] = 21'b111111111110100110100;
        x_t[4] = 21'b111111111111000111100;
        x_t[5] = 21'b111111111111000000011;
        x_t[6] = 21'b111111111101000010001;
        x_t[7] = 21'b111111111011011001011;
        x_t[8] = 21'b111111111101100001110;
        x_t[9] = 21'b111111111110011000101;
        x_t[10] = 21'b111111111111011001100;
        x_t[11] = 21'b111111111111111111001;
        x_t[12] = 21'b000000000000011010101;
        x_t[13] = 21'b111111111111001011100;
        x_t[14] = 21'b111111111101100010011;
        x_t[15] = 21'b111111111110100010000;
        x_t[16] = 21'b111111111110111100000;
        x_t[17] = 21'b000000000000011100100;
        x_t[18] = 21'b000000000000100111110;
        x_t[19] = 21'b000000000001000111001;
        x_t[20] = 21'b000000000001011111101;
        x_t[21] = 21'b111111111001011110101;
        x_t[22] = 21'b111111111001001010001;
        x_t[23] = 21'b111111111010010001101;
        x_t[24] = 21'b111111111001000010010;
        x_t[25] = 21'b111111111001000110111;
        x_t[26] = 21'b111111111010110001110;
        x_t[27] = 21'b111111111011000111001;
        x_t[28] = 21'b111111111010101111100;
        x_t[29] = 21'b111111111000100110101;
        x_t[30] = 21'b111111111010010110110;
        x_t[31] = 21'b111111111011011010101;
        x_t[32] = 21'b111111111011101000111;
        x_t[33] = 21'b111111111100011010001;
        x_t[34] = 21'b111111111101010011001;
        x_t[35] = 21'b111111111101000111100;
        x_t[36] = 21'b111111111100111100110;
        x_t[37] = 21'b111111111101001101100;
        x_t[38] = 21'b111111111001010010110;
        x_t[39] = 21'b111111111101010101010;
        x_t[40] = 21'b111111111001110000110;
        x_t[41] = 21'b000000000000000010000;
        x_t[42] = 21'b111111110111101110110;
        x_t[43] = 21'b000000000000110011011;
        x_t[44] = 21'b111111111100001000100;
        x_t[45] = 21'b111111111111100000101;
        x_t[46] = 21'b111111111111101000000;
        x_t[47] = 21'b111111111111011111000;
        x_t[48] = 21'b000000000000010101111;
        x_t[49] = 21'b000000000000100101011;
        x_t[50] = 21'b000000000000101110000;
        x_t[51] = 21'b000000000010001110011;
        x_t[52] = 21'b000000000001011001010;
        x_t[53] = 21'b000000000010000100000;
        x_t[54] = 21'b000000000001011000111;
        x_t[55] = 21'b000000000001100100111;
        x_t[56] = 21'b000000000001101000010;
        x_t[57] = 21'b000000000011011111110;
        x_t[58] = 21'b000000000011011101110;
        x_t[59] = 21'b000000000010110000111;
        x_t[60] = 21'b000000000011100101001;
        x_t[61] = 21'b000000000100110101110;
        x_t[62] = 21'b000000000001011011111;
        x_t[63] = 21'b000000000011010011100;
        
        h_t_prev[0] = 21'b111111111001001101010;
        h_t_prev[1] = 21'b111111111011110000100;
        h_t_prev[2] = 21'b111111111100001010000;
        h_t_prev[3] = 21'b111111111110100110100;
        h_t_prev[4] = 21'b111111111111000111100;
        h_t_prev[5] = 21'b111111111111000000011;
        h_t_prev[6] = 21'b111111111101000010001;
        h_t_prev[7] = 21'b111111111011011001011;
        h_t_prev[8] = 21'b111111111101100001110;
        h_t_prev[9] = 21'b111111111110011000101;
        h_t_prev[10] = 21'b111111111111011001100;
        h_t_prev[11] = 21'b111111111111111111001;
        h_t_prev[12] = 21'b000000000000011010101;
        h_t_prev[13] = 21'b111111111111001011100;
        h_t_prev[14] = 21'b111111111101100010011;
        h_t_prev[15] = 21'b111111111110100010000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 65 timeout!");
                $fdisplay(fd_cycles, "Test Vector  65: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  65: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 65");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 66
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111001101111110;
        x_t[1] = 21'b111111111100100001011;
        x_t[2] = 21'b111111111100111010100;
        x_t[3] = 21'b111111111110101011011;
        x_t[4] = 21'b111111111111010110101;
        x_t[5] = 21'b111111111111110010010;
        x_t[6] = 21'b111111111110111110100;
        x_t[7] = 21'b111111111100010001011;
        x_t[8] = 21'b111111111110001011000;
        x_t[9] = 21'b111111111110100010101;
        x_t[10] = 21'b111111111110101101011;
        x_t[11] = 21'b111111111111111010000;
        x_t[12] = 21'b000000000000100110011;
        x_t[13] = 21'b000000000000101011000;
        x_t[14] = 21'b111111111101010111110;
        x_t[15] = 21'b111111111110010111111;
        x_t[16] = 21'b111111111110101101001;
        x_t[17] = 21'b111111111111011100011;
        x_t[18] = 21'b111111111110111110011;
        x_t[19] = 21'b111111111111110100110;
        x_t[20] = 21'b000000000000100111011;
        x_t[21] = 21'b111111111001001011011;
        x_t[22] = 21'b111111111001011101010;
        x_t[23] = 21'b111111111010110100011;
        x_t[24] = 21'b111111111000111001001;
        x_t[25] = 21'b111111111001000011111;
        x_t[26] = 21'b111111111010111010001;
        x_t[27] = 21'b111111111011111010010;
        x_t[28] = 21'b111111111011101011010;
        x_t[29] = 21'b111111111000110111010;
        x_t[30] = 21'b111111111011000101101;
        x_t[31] = 21'b111111111011111001101;
        x_t[32] = 21'b111111111011101000111;
        x_t[33] = 21'b111111111100011110110;
        x_t[34] = 21'b111111111101100001011;
        x_t[35] = 21'b111111111101011011010;
        x_t[36] = 21'b111111111110001100010;
        x_t[37] = 21'b111111111110000010100;
        x_t[38] = 21'b111111111001011100110;
        x_t[39] = 21'b111111111111100000111;
        x_t[40] = 21'b111111111010000001001;
        x_t[41] = 21'b000000000101001000110;
        x_t[42] = 21'b111111110111111010100;
        x_t[43] = 21'b111111111011110101010;
        x_t[44] = 21'b111111111010111111111;
        x_t[45] = 21'b111111111101010101010;
        x_t[46] = 21'b111111111110011010011;
        x_t[47] = 21'b111111111111001011001;
        x_t[48] = 21'b000000000000011010101;
        x_t[49] = 21'b000000000000000100111;
        x_t[50] = 21'b111111111111110000010;
        x_t[51] = 21'b000000000000111100010;
        x_t[52] = 21'b000000000000010001101;
        x_t[53] = 21'b000000000001010111100;
        x_t[54] = 21'b000000000000101111000;
        x_t[55] = 21'b000000000001011100010;
        x_t[56] = 21'b000000000001010111001;
        x_t[57] = 21'b000000000011000110001;
        x_t[58] = 21'b000000000011000011101;
        x_t[59] = 21'b000000000010100101000;
        x_t[60] = 21'b000000000011000110100;
        x_t[61] = 21'b000000000100010100101;
        x_t[62] = 21'b000000000000101011110;
        x_t[63] = 21'b000000000010111001001;
        
        h_t_prev[0] = 21'b111111111001101111110;
        h_t_prev[1] = 21'b111111111100100001011;
        h_t_prev[2] = 21'b111111111100111010100;
        h_t_prev[3] = 21'b111111111110101011011;
        h_t_prev[4] = 21'b111111111111010110101;
        h_t_prev[5] = 21'b111111111111110010010;
        h_t_prev[6] = 21'b111111111110111110100;
        h_t_prev[7] = 21'b111111111100010001011;
        h_t_prev[8] = 21'b111111111110001011000;
        h_t_prev[9] = 21'b111111111110100010101;
        h_t_prev[10] = 21'b111111111110101101011;
        h_t_prev[11] = 21'b111111111111111010000;
        h_t_prev[12] = 21'b000000000000100110011;
        h_t_prev[13] = 21'b000000000000101011000;
        h_t_prev[14] = 21'b111111111101010111110;
        h_t_prev[15] = 21'b111111111110010111111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 66 timeout!");
                $fdisplay(fd_cycles, "Test Vector  66: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  66: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 66");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 67
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111010100110000;
        x_t[1] = 21'b111111111101010111010;
        x_t[2] = 21'b111111111101010111110;
        x_t[3] = 21'b111111111110100001110;
        x_t[4] = 21'b111111111111000111100;
        x_t[5] = 21'b111111111111110010010;
        x_t[6] = 21'b000000000000000011000;
        x_t[7] = 21'b111111111101011000101;
        x_t[8] = 21'b111111111110110100010;
        x_t[9] = 21'b111111111110001110101;
        x_t[10] = 21'b111111111101110111101;
        x_t[11] = 21'b111111111111000010000;
        x_t[12] = 21'b000000000000001111000;
        x_t[13] = 21'b000000000001010011111;
        x_t[14] = 21'b111111111101111100101;
        x_t[15] = 21'b111111111110111011100;
        x_t[16] = 21'b111111111110100011010;
        x_t[17] = 21'b111111111110111110110;
        x_t[18] = 21'b111111111101111111001;
        x_t[19] = 21'b111111111110111101110;
        x_t[20] = 21'b000000000000101101101;
        x_t[21] = 21'b111111111010000101011;
        x_t[22] = 21'b111111111010000110100;
        x_t[23] = 21'b111111111011001110100;
        x_t[24] = 21'b111111111001110110001;
        x_t[25] = 21'b111111111001111000101;
        x_t[26] = 21'b111111111011010111110;
        x_t[27] = 21'b111111111100000110000;
        x_t[28] = 21'b111111111011101011010;
        x_t[29] = 21'b111111111010001010011;
        x_t[30] = 21'b111111111011001101011;
        x_t[31] = 21'b111111111100011000101;
        x_t[32] = 21'b111111111100011010111;
        x_t[33] = 21'b111111111100111010100;
        x_t[34] = 21'b111111111101101111101;
        x_t[35] = 21'b111111111101110011111;
        x_t[36] = 21'b111111111110001100010;
        x_t[37] = 21'b111111111101110010010;
        x_t[38] = 21'b111111111011011010111;
        x_t[39] = 21'b111111111111000011100;
        x_t[40] = 21'b111111111100000011100;
        x_t[41] = 21'b000000000010011011000;
        x_t[42] = 21'b111111110111011100111;
        x_t[43] = 21'b000000000000110011011;
        x_t[44] = 21'b111111111100011110111;
        x_t[45] = 21'b111111111111000001101;
        x_t[46] = 21'b111111111111110111101;
        x_t[47] = 21'b000000000000000110110;
        x_t[48] = 21'b000000000001001010010;
        x_t[49] = 21'b000000000000011100001;
        x_t[50] = 21'b111111111111111001110;
        x_t[51] = 21'b000000000000101001000;
        x_t[52] = 21'b000000000000000010011;
        x_t[53] = 21'b000000000001110011011;
        x_t[54] = 21'b000000000001111100111;
        x_t[55] = 21'b000000000001101101100;
        x_t[56] = 21'b000000000001100100000;
        x_t[57] = 21'b000000000011001010011;
        x_t[58] = 21'b000000000011010101001;
        x_t[59] = 21'b000000000011000100101;
        x_t[60] = 21'b000000000010110111001;
        x_t[61] = 21'b000000000100001000010;
        x_t[62] = 21'b000000000000101011110;
        x_t[63] = 21'b000000000010111101100;
        
        h_t_prev[0] = 21'b111111111010100110000;
        h_t_prev[1] = 21'b111111111101010111010;
        h_t_prev[2] = 21'b111111111101010111110;
        h_t_prev[3] = 21'b111111111110100001110;
        h_t_prev[4] = 21'b111111111111000111100;
        h_t_prev[5] = 21'b111111111111110010010;
        h_t_prev[6] = 21'b000000000000000011000;
        h_t_prev[7] = 21'b111111111101011000101;
        h_t_prev[8] = 21'b111111111110110100010;
        h_t_prev[9] = 21'b111111111110001110101;
        h_t_prev[10] = 21'b111111111101110111101;
        h_t_prev[11] = 21'b111111111111000010000;
        h_t_prev[12] = 21'b000000000000001111000;
        h_t_prev[13] = 21'b000000000001010011111;
        h_t_prev[14] = 21'b111111111101111100101;
        h_t_prev[15] = 21'b111111111110111011100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 67 timeout!");
                $fdisplay(fd_cycles, "Test Vector  67: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  67: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 67");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 68
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111100001101101;
        x_t[1] = 21'b111111111110010010000;
        x_t[2] = 21'b111111111101111001101;
        x_t[3] = 21'b111111111110100110100;
        x_t[4] = 21'b111111111110111101011;
        x_t[5] = 21'b111111111111010001000;
        x_t[6] = 21'b111111111110111110100;
        x_t[7] = 21'b111111111110101010000;
        x_t[8] = 21'b111111111111011000011;
        x_t[9] = 21'b111111111110100111101;
        x_t[10] = 21'b111111111110011110110;
        x_t[11] = 21'b111111111110011110011;
        x_t[12] = 21'b111111111110111101000;
        x_t[13] = 21'b111111111110010101000;
        x_t[14] = 21'b111111111111000110100;
        x_t[15] = 21'b111111111111001111110;
        x_t[16] = 21'b111111111111000001000;
        x_t[17] = 21'b111111111111000011110;
        x_t[18] = 21'b111111111101011010010;
        x_t[19] = 21'b111111111101111011111;
        x_t[20] = 21'b111111111111000011010;
        x_t[21] = 21'b111111111010000101011;
        x_t[22] = 21'b111111111001111100111;
        x_t[23] = 21'b111111111011000101111;
        x_t[24] = 21'b111111111001111111010;
        x_t[25] = 21'b111111111010001000010;
        x_t[26] = 21'b111111111011100000001;
        x_t[27] = 21'b111111111100000110000;
        x_t[28] = 21'b111111111011101011010;
        x_t[29] = 21'b111111111010011111010;
        x_t[30] = 21'b111111111011111000011;
        x_t[31] = 21'b111111111100001111110;
        x_t[32] = 21'b111111111100011111011;
        x_t[33] = 21'b111111111100111010100;
        x_t[34] = 21'b111111111101110100100;
        x_t[35] = 21'b111111111110000010110;
        x_t[36] = 21'b111111111101011111101;
        x_t[37] = 21'b111111111101100110000;
        x_t[38] = 21'b111111111010111100101;
        x_t[39] = 21'b111111111100101001001;
        x_t[40] = 21'b111111111010110111100;
        x_t[41] = 21'b111111111010000011100;
        x_t[42] = 21'b111111111000011110001;
        x_t[43] = 21'b111111111100110111000;
        x_t[44] = 21'b111111111100001000100;
        x_t[45] = 21'b111111111101011101000;
        x_t[46] = 21'b111111111110101111000;
        x_t[47] = 21'b111111111110110010010;
        x_t[48] = 21'b111111111111101011000;
        x_t[49] = 21'b111111111111011011010;
        x_t[50] = 21'b111111111111100010000;
        x_t[51] = 21'b111111111111110011111;
        x_t[52] = 21'b111111111111000101000;
        x_t[53] = 21'b000000000000001111001;
        x_t[54] = 21'b000000000000010111000;
        x_t[55] = 21'b111111111111000101001;
        x_t[56] = 21'b111111111111010110010;
        x_t[57] = 21'b000000000001101100101;
        x_t[58] = 21'b000000000001110000110;
        x_t[59] = 21'b000000000001100101111;
        x_t[60] = 21'b000000000001100010111;
        x_t[61] = 21'b000000000010110101100;
        x_t[62] = 21'b111111111111101100111;
        x_t[63] = 21'b000000000001011100101;
        
        h_t_prev[0] = 21'b111111111100001101101;
        h_t_prev[1] = 21'b111111111110010010000;
        h_t_prev[2] = 21'b111111111101111001101;
        h_t_prev[3] = 21'b111111111110100110100;
        h_t_prev[4] = 21'b111111111110111101011;
        h_t_prev[5] = 21'b111111111111010001000;
        h_t_prev[6] = 21'b111111111110111110100;
        h_t_prev[7] = 21'b111111111110101010000;
        h_t_prev[8] = 21'b111111111111011000011;
        h_t_prev[9] = 21'b111111111110100111101;
        h_t_prev[10] = 21'b111111111110011110110;
        h_t_prev[11] = 21'b111111111110011110011;
        h_t_prev[12] = 21'b111111111110111101000;
        h_t_prev[13] = 21'b111111111110010101000;
        h_t_prev[14] = 21'b111111111111000110100;
        h_t_prev[15] = 21'b111111111111001111110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 68 timeout!");
                $fdisplay(fd_cycles, "Test Vector  68: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  68: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 68");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 69
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111011111001111;
        x_t[1] = 21'b111111111101111001100;
        x_t[2] = 21'b111111111101110000000;
        x_t[3] = 21'b111111111110100110100;
        x_t[4] = 21'b111111111110111000010;
        x_t[5] = 21'b111111111110111010111;
        x_t[6] = 21'b111111111101101101101;
        x_t[7] = 21'b111111111101100010110;
        x_t[8] = 21'b111111111110111001011;
        x_t[9] = 21'b111111111110110110101;
        x_t[10] = 21'b111111111111001010110;
        x_t[11] = 21'b111111111111100000101;
        x_t[12] = 21'b111111111110110001010;
        x_t[13] = 21'b111111111101111001110;
        x_t[14] = 21'b111111111101001101010;
        x_t[15] = 21'b111111111110010111111;
        x_t[16] = 21'b111111111111001010111;
        x_t[17] = 21'b111111111111100001011;
        x_t[18] = 21'b111111111110101001010;
        x_t[19] = 21'b111111111110110010111;
        x_t[20] = 21'b111111111111100010100;
        x_t[21] = 21'b111111111001011011111;
        x_t[22] = 21'b111111111001000111000;
        x_t[23] = 21'b111111111010000110000;
        x_t[24] = 21'b111111111001000101011;
        x_t[25] = 21'b111111111001010110100;
        x_t[26] = 21'b111111111011000110111;
        x_t[27] = 21'b111111111011011010111;
        x_t[28] = 21'b111111111010111000111;
        x_t[29] = 21'b111111111001101101010;
        x_t[30] = 21'b111111111100101111000;
        x_t[31] = 21'b111111111100100001100;
        x_t[32] = 21'b111111111100011010111;
        x_t[33] = 21'b111111111100111111001;
        x_t[34] = 21'b111111111101111001010;
        x_t[35] = 21'b111111111101110011111;
        x_t[36] = 21'b111111111100111100110;
        x_t[37] = 21'b111111111110000010100;
        x_t[38] = 21'b111111111011010000110;
        x_t[39] = 21'b111111111101110010101;
        x_t[40] = 21'b111111111100101001101;
        x_t[41] = 21'b000000000010000110001;
        x_t[42] = 21'b111111111000011000010;
        x_t[43] = 21'b111111111101000010000;
        x_t[44] = 21'b111111111100010011101;
        x_t[45] = 21'b111111111110011011000;
        x_t[46] = 21'b111111111101101011110;
        x_t[47] = 21'b111111111110001010100;
        x_t[48] = 21'b111111111111111110000;
        x_t[49] = 21'b000000000000001001100;
        x_t[50] = 21'b000000000000110010110;
        x_t[51] = 21'b000000000001100111110;
        x_t[52] = 21'b000000000001001111001;
        x_t[53] = 21'b000000000001110011011;
        x_t[54] = 21'b000000000001110000111;
        x_t[55] = 21'b111111111110100010101;
        x_t[56] = 21'b111111111111010001111;
        x_t[57] = 21'b000000000010001010100;
        x_t[58] = 21'b000000000010110110100;
        x_t[59] = 21'b000000000010100101000;
        x_t[60] = 21'b000000000000000011000;
        x_t[61] = 21'b000000000001100010110;
        x_t[62] = 21'b111111111111000100010;
        x_t[63] = 21'b111111111111101110101;
        
        h_t_prev[0] = 21'b111111111011111001111;
        h_t_prev[1] = 21'b111111111101111001100;
        h_t_prev[2] = 21'b111111111101110000000;
        h_t_prev[3] = 21'b111111111110100110100;
        h_t_prev[4] = 21'b111111111110111000010;
        h_t_prev[5] = 21'b111111111110111010111;
        h_t_prev[6] = 21'b111111111101101101101;
        h_t_prev[7] = 21'b111111111101100010110;
        h_t_prev[8] = 21'b111111111110111001011;
        h_t_prev[9] = 21'b111111111110110110101;
        h_t_prev[10] = 21'b111111111111001010110;
        h_t_prev[11] = 21'b111111111111100000101;
        h_t_prev[12] = 21'b111111111110110001010;
        h_t_prev[13] = 21'b111111111101111001110;
        h_t_prev[14] = 21'b111111111101001101010;
        h_t_prev[15] = 21'b111111111110010111111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 69 timeout!");
                $fdisplay(fd_cycles, "Test Vector  69: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  69: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 69");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 70
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111011111110110;
        x_t[1] = 21'b111111111110000011010;
        x_t[2] = 21'b111111111110100000100;
        x_t[3] = 21'b111111111111110011111;
        x_t[4] = 21'b000000000000010011010;
        x_t[5] = 21'b000000000000011110101;
        x_t[6] = 21'b111111111111101010001;
        x_t[7] = 21'b111111111110010000101;
        x_t[8] = 21'b111111111111100010110;
        x_t[9] = 21'b111111111111101101110;
        x_t[10] = 21'b000000000000000000101;
        x_t[11] = 21'b000000000000100010111;
        x_t[12] = 21'b000000000000111101110;
        x_t[13] = 21'b000000000000100100001;
        x_t[14] = 21'b111111111100111101011;
        x_t[15] = 21'b111111111110101100010;
        x_t[16] = 21'b111111111111101000101;
        x_t[17] = 21'b000000000000100001100;
        x_t[18] = 21'b000000000000100111110;
        x_t[19] = 21'b000000000000110001001;
        x_t[20] = 21'b000000000000101101101;
        x_t[21] = 21'b111111111001101111010;
        x_t[22] = 21'b111111111001110110101;
        x_t[23] = 21'b111111111010110001100;
        x_t[24] = 21'b111111111001010111101;
        x_t[25] = 21'b111111111001100010111;
        x_t[26] = 21'b111111111011100000001;
        x_t[27] = 21'b111111111011111010010;
        x_t[28] = 21'b111111111011001111000;
        x_t[29] = 21'b111111111010100111100;
        x_t[30] = 21'b111111111011111000011;
        x_t[31] = 21'b111111111100011000101;
        x_t[32] = 21'b111111111100011111011;
        x_t[33] = 21'b111111111101000011110;
        x_t[34] = 21'b111111111110001100010;
        x_t[35] = 21'b111111111101110011111;
        x_t[36] = 21'b111111111101010101101;
        x_t[37] = 21'b111111111110010110111;
        x_t[38] = 21'b111111111011000001101;
        x_t[39] = 21'b111111111101101011010;
        x_t[40] = 21'b111111111010000001001;
        x_t[41] = 21'b111111111100110001010;
        x_t[42] = 21'b111111110111101000110;
        x_t[43] = 21'b000000000000011101011;
        x_t[44] = 21'b111111111011011011111;
        x_t[45] = 21'b111111111100110110011;
        x_t[46] = 21'b111111111100110010110;
        x_t[47] = 21'b111111111100111111111;
        x_t[48] = 21'b111111111110110110101;
        x_t[49] = 21'b111111111110111111011;
        x_t[50] = 21'b000000000000000011010;
        x_t[51] = 21'b000000000001100010111;
        x_t[52] = 21'b000000000000111111110;
        x_t[53] = 21'b000000000001000110110;
        x_t[54] = 21'b000000000000101111000;
        x_t[55] = 21'b111111111101101110111;
        x_t[56] = 21'b111111111110011010000;
        x_t[57] = 21'b000000000001010111011;
        x_t[58] = 21'b000000000010000010010;
        x_t[59] = 21'b000000000001100101111;
        x_t[60] = 21'b111111111110111010001;
        x_t[61] = 21'b000000000000100100101;
        x_t[62] = 21'b111111111110101010011;
        x_t[63] = 21'b111111111110010010010;
        
        h_t_prev[0] = 21'b111111111011111110110;
        h_t_prev[1] = 21'b111111111110000011010;
        h_t_prev[2] = 21'b111111111110100000100;
        h_t_prev[3] = 21'b111111111111110011111;
        h_t_prev[4] = 21'b000000000000010011010;
        h_t_prev[5] = 21'b000000000000011110101;
        h_t_prev[6] = 21'b111111111111101010001;
        h_t_prev[7] = 21'b111111111110010000101;
        h_t_prev[8] = 21'b111111111111100010110;
        h_t_prev[9] = 21'b111111111111101101110;
        h_t_prev[10] = 21'b000000000000000000101;
        h_t_prev[11] = 21'b000000000000100010111;
        h_t_prev[12] = 21'b000000000000111101110;
        h_t_prev[13] = 21'b000000000000100100001;
        h_t_prev[14] = 21'b111111111100111101011;
        h_t_prev[15] = 21'b111111111110101100010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 70 timeout!");
                $fdisplay(fd_cycles, "Test Vector  70: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  70: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 70");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 71
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111010001000011;
        x_t[1] = 21'b111111111100011100100;
        x_t[2] = 21'b111111111100110101110;
        x_t[3] = 21'b111111111110110101000;
        x_t[4] = 21'b111111111111011011101;
        x_t[5] = 21'b111111111111011100001;
        x_t[6] = 21'b111111111110001100110;
        x_t[7] = 21'b111111111011110111111;
        x_t[8] = 21'b111111111101110001010;
        x_t[9] = 21'b111111111101110101100;
        x_t[10] = 21'b111111111110011110110;
        x_t[11] = 21'b111111111111110101000;
        x_t[12] = 21'b000000000000100110011;
        x_t[13] = 21'b111111111111000100110;
        x_t[14] = 21'b111111111011111000111;
        x_t[15] = 21'b111111111100111100011;
        x_t[16] = 21'b111111111110000101100;
        x_t[17] = 21'b111111111111100001011;
        x_t[18] = 21'b000000000000001101011;
        x_t[19] = 21'b000000000000110001001;
        x_t[20] = 21'b000000000000001110010;
        x_t[21] = 21'b111111111001001110001;
        x_t[22] = 21'b111111111001011101010;
        x_t[23] = 21'b111111111010101110101;
        x_t[24] = 21'b111111111000111111010;
        x_t[25] = 21'b111111111001000110111;
        x_t[26] = 21'b111111111010111010001;
        x_t[27] = 21'b111111111011111010010;
        x_t[28] = 21'b111111111011011000011;
        x_t[29] = 21'b111111111001110001100;
        x_t[30] = 21'b111111111011110000100;
        x_t[31] = 21'b111111111100000010100;
        x_t[32] = 21'b111111111011101101011;
        x_t[33] = 21'b111111111100011010001;
        x_t[34] = 21'b111111111101110100100;
        x_t[35] = 21'b111111111101101111000;
        x_t[36] = 21'b111111111101110011100;
        x_t[37] = 21'b111111111110010010110;
        x_t[38] = 21'b111111111001011100110;
        x_t[39] = 21'b111111111110010111011;
        x_t[40] = 21'b111111111000101010001;
        x_t[41] = 21'b111111111100111000010;
        x_t[42] = 21'b111111111000010010010;
        x_t[43] = 21'b111111111111011011101;
        x_t[44] = 21'b111111111011100001011;
        x_t[45] = 21'b111111111110001011100;
        x_t[46] = 21'b111111111101101011110;
        x_t[47] = 21'b111111111101100111101;
        x_t[48] = 21'b111111111111000000001;
        x_t[49] = 21'b111111111111010010000;
        x_t[50] = 21'b000000000000110010110;
        x_t[51] = 21'b000000000010101011011;
        x_t[52] = 21'b000000000010000111011;
        x_t[53] = 21'b000000000010010100110;
        x_t[54] = 21'b000000000001110110111;
        x_t[55] = 21'b111111111111000101001;
        x_t[56] = 21'b111111111111100011001;
        x_t[57] = 21'b000000000010101100101;
        x_t[58] = 21'b000000000011000011101;
        x_t[59] = 21'b000000000010100001001;
        x_t[60] = 21'b111111111111000001110;
        x_t[61] = 21'b000000000000100100101;
        x_t[62] = 21'b111111111110110101011;
        x_t[63] = 21'b111111111110000101000;
        
        h_t_prev[0] = 21'b111111111010001000011;
        h_t_prev[1] = 21'b111111111100011100100;
        h_t_prev[2] = 21'b111111111100110101110;
        h_t_prev[3] = 21'b111111111110110101000;
        h_t_prev[4] = 21'b111111111111011011101;
        h_t_prev[5] = 21'b111111111111011100001;
        h_t_prev[6] = 21'b111111111110001100110;
        h_t_prev[7] = 21'b111111111011110111111;
        h_t_prev[8] = 21'b111111111101110001010;
        h_t_prev[9] = 21'b111111111101110101100;
        h_t_prev[10] = 21'b111111111110011110110;
        h_t_prev[11] = 21'b111111111111110101000;
        h_t_prev[12] = 21'b000000000000100110011;
        h_t_prev[13] = 21'b111111111111000100110;
        h_t_prev[14] = 21'b111111111011111000111;
        h_t_prev[15] = 21'b111111111100111100011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 71 timeout!");
                $fdisplay(fd_cycles, "Test Vector  71: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  71: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 71");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 72
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111010101010111;
        x_t[1] = 21'b111111111101001101100;
        x_t[2] = 21'b111111111101001110000;
        x_t[3] = 21'b111111111111010110111;
        x_t[4] = 21'b000000000000011101011;
        x_t[5] = 21'b000000000001000101100;
        x_t[6] = 21'b111111111111010001010;
        x_t[7] = 21'b111111111101011000101;
        x_t[8] = 21'b111111111110010000001;
        x_t[9] = 21'b111111111110011101101;
        x_t[10] = 21'b111111111111011110011;
        x_t[11] = 21'b000000000001010101110;
        x_t[12] = 21'b000000000010011011011;
        x_t[13] = 21'b000000000001000110010;
        x_t[14] = 21'b111111111100111101011;
        x_t[15] = 21'b111111111101010101110;
        x_t[16] = 21'b111111111110101000010;
        x_t[17] = 21'b000000000000011100100;
        x_t[18] = 21'b000000000010000110101;
        x_t[19] = 21'b000000000010100100100;
        x_t[20] = 21'b000000000010011000000;
        x_t[21] = 21'b111111111010001010111;
        x_t[22] = 21'b111111111010011100101;
        x_t[23] = 21'b111111111011010001011;
        x_t[24] = 21'b111111111001110011000;
        x_t[25] = 21'b111111111001110101100;
        x_t[26] = 21'b111111111100000010000;
        x_t[27] = 21'b111111111100110101010;
        x_t[28] = 21'b111111111011111011000;
        x_t[29] = 21'b111111111010011111010;
        x_t[30] = 21'b111111111101001110010;
        x_t[31] = 21'b111111111101011011010;
        x_t[32] = 21'b111111111100011111011;
        x_t[33] = 21'b111111111101010001101;
        x_t[34] = 21'b111111111110110111001;
        x_t[35] = 21'b111111111110110100001;
        x_t[36] = 21'b111111111110111001000;
        x_t[37] = 21'b111111111110001110110;
        x_t[38] = 21'b111111111011100101000;
        x_t[39] = 21'b111111111111011001100;
        x_t[40] = 21'b111111111100111111011;
        x_t[41] = 21'b111111111110100111100;
        x_t[42] = 21'b111111111000111011110;
        x_t[43] = 21'b000000000000101000011;
        x_t[44] = 21'b111111111100101010000;
        x_t[45] = 21'b000000000000000111010;
        x_t[46] = 21'b111111111110101111000;
        x_t[47] = 21'b111111111110011001011;
        x_t[48] = 21'b111111111111010011001;
        x_t[49] = 21'b000000000000001110001;
        x_t[50] = 21'b000000000001110000100;
        x_t[51] = 21'b000000000011101111000;
        x_t[52] = 21'b000000000010111111101;
        x_t[53] = 21'b000000000011010010000;
        x_t[54] = 21'b000000000010101100111;
        x_t[55] = 21'b000000000000001010010;
        x_t[56] = 21'b000000000000010110101;
        x_t[57] = 21'b000000000011010111010;
        x_t[58] = 21'b000000000011101111010;
        x_t[59] = 21'b000000000011001000100;
        x_t[60] = 21'b000000000000010010011;
        x_t[61] = 21'b000000000010001000000;
        x_t[62] = 21'b000000000000010001111;
        x_t[63] = 21'b111111111111101110101;
        
        h_t_prev[0] = 21'b111111111010101010111;
        h_t_prev[1] = 21'b111111111101001101100;
        h_t_prev[2] = 21'b111111111101001110000;
        h_t_prev[3] = 21'b111111111111010110111;
        h_t_prev[4] = 21'b000000000000011101011;
        h_t_prev[5] = 21'b000000000001000101100;
        h_t_prev[6] = 21'b111111111111010001010;
        h_t_prev[7] = 21'b111111111101011000101;
        h_t_prev[8] = 21'b111111111110010000001;
        h_t_prev[9] = 21'b111111111110011101101;
        h_t_prev[10] = 21'b111111111111011110011;
        h_t_prev[11] = 21'b000000000001010101110;
        h_t_prev[12] = 21'b000000000010011011011;
        h_t_prev[13] = 21'b000000000001000110010;
        h_t_prev[14] = 21'b111111111100111101011;
        h_t_prev[15] = 21'b111111111101010101110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 72 timeout!");
                $fdisplay(fd_cycles, "Test Vector  72: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  72: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 72");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 73
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111100011100011;
        x_t[1] = 21'b111111111110001101001;
        x_t[2] = 21'b111111111110000011011;
        x_t[3] = 21'b000000000000000010011;
        x_t[4] = 21'b000000000000110001100;
        x_t[5] = 21'b000000000000111010011;
        x_t[6] = 21'b111111111111011101101;
        x_t[7] = 21'b111111111101101101000;
        x_t[8] = 21'b111111111110010000001;
        x_t[9] = 21'b111111111110110110101;
        x_t[10] = 21'b111111111111110110110;
        x_t[11] = 21'b000000000001000110100;
        x_t[12] = 21'b000000000001101100101;
        x_t[13] = 21'b000000000000001000111;
        x_t[14] = 21'b111111111100001000101;
        x_t[15] = 21'b111111111101010000101;
        x_t[16] = 21'b111111111110111100000;
        x_t[17] = 21'b000000000000100110011;
        x_t[18] = 21'b000000000001100111000;
        x_t[19] = 21'b000000000001101101100;
        x_t[20] = 21'b000000000001010011001;
        x_t[21] = 21'b111111111010111111011;
        x_t[22] = 21'b111111111011001001001;
        x_t[23] = 21'b111111111011101011100;
        x_t[24] = 21'b111111111010100110110;
        x_t[25] = 21'b111111111010101101100;
        x_t[26] = 21'b111111111100110000011;
        x_t[27] = 21'b111111111100111001001;
        x_t[28] = 21'b111111111011101011010;
        x_t[29] = 21'b111111111011010101010;
        x_t[30] = 21'b111111111110010100100;
        x_t[31] = 21'b111111111101010110110;
        x_t[32] = 21'b111111111101010101111;
        x_t[33] = 21'b111111111101101101011;
        x_t[34] = 21'b111111111110111011111;
        x_t[35] = 21'b111111111111000010111;
        x_t[36] = 21'b111111111110000111011;
        x_t[37] = 21'b111111111110001110110;
        x_t[38] = 21'b111111111100101011100;
        x_t[39] = 21'b111111111110010111011;
        x_t[40] = 21'b111111111011110011010;
        x_t[41] = 21'b000000000001010101011;
        x_t[42] = 21'b111111111000101111111;
        x_t[43] = 21'b111111111101101101111;
        x_t[44] = 21'b111111111100111010110;
        x_t[45] = 21'b111111111101000101111;
        x_t[46] = 21'b111111111111000011110;
        x_t[47] = 21'b111111111110001010100;
        x_t[48] = 21'b111111111111001110011;
        x_t[49] = 21'b111111111111101001001;
        x_t[50] = 21'b000000000000110111100;
        x_t[51] = 21'b000000000001100010111;
        x_t[52] = 21'b000000000000101011010;
        x_t[53] = 21'b000000000000100101011;
        x_t[54] = 21'b111111111111100001001;
        x_t[55] = 21'b111111111111100111110;
        x_t[56] = 21'b111111111111110000000;
        x_t[57] = 21'b000000000001101100101;
        x_t[58] = 21'b000000000001001001100;
        x_t[59] = 21'b000000000000001111000;
        x_t[60] = 21'b000000000000110100111;
        x_t[61] = 21'b000000000001111111101;
        x_t[62] = 21'b111111111111111011110;
        x_t[63] = 21'b111111111111011000101;
        
        h_t_prev[0] = 21'b111111111100011100011;
        h_t_prev[1] = 21'b111111111110001101001;
        h_t_prev[2] = 21'b111111111110000011011;
        h_t_prev[3] = 21'b000000000000000010011;
        h_t_prev[4] = 21'b000000000000110001100;
        h_t_prev[5] = 21'b000000000000111010011;
        h_t_prev[6] = 21'b111111111111011101101;
        h_t_prev[7] = 21'b111111111101101101000;
        h_t_prev[8] = 21'b111111111110010000001;
        h_t_prev[9] = 21'b111111111110110110101;
        h_t_prev[10] = 21'b111111111111110110110;
        h_t_prev[11] = 21'b000000000001000110100;
        h_t_prev[12] = 21'b000000000001101100101;
        h_t_prev[13] = 21'b000000000000001000111;
        h_t_prev[14] = 21'b111111111100001000101;
        h_t_prev[15] = 21'b111111111101010000101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 73 timeout!");
                $fdisplay(fd_cycles, "Test Vector  73: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  73: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 73");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 74
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111100110101000;
        x_t[1] = 21'b111111111110111110000;
        x_t[2] = 21'b111111111110011011101;
        x_t[3] = 21'b000000000000010000111;
        x_t[4] = 21'b000000000000010011010;
        x_t[5] = 21'b000000000000001000100;
        x_t[6] = 21'b111111111110111110100;
        x_t[7] = 21'b111111111110011010110;
        x_t[8] = 21'b111111111110111001011;
        x_t[9] = 21'b111111111111011110110;
        x_t[10] = 21'b000000000000001111010;
        x_t[11] = 21'b000000000001000110100;
        x_t[12] = 21'b000000000001001001100;
        x_t[13] = 21'b111111111111110100011;
        x_t[14] = 21'b111111111101011101000;
        x_t[15] = 21'b111111111110100010000;
        x_t[16] = 21'b111111111111101101101;
        x_t[17] = 21'b000000000001000100000;
        x_t[18] = 21'b000000000000110010011;
        x_t[19] = 21'b000000000000110001001;
        x_t[20] = 21'b000000000000100111011;
        x_t[21] = 21'b111111111011010010110;
        x_t[22] = 21'b111111111011010010101;
        x_t[23] = 21'b111111111100000010110;
        x_t[24] = 21'b111111111010111100001;
        x_t[25] = 21'b111111111011000011010;
        x_t[26] = 21'b111111111101010010010;
        x_t[27] = 21'b111111111101010000110;
        x_t[28] = 21'b111111111100010001001;
        x_t[29] = 21'b111111111011001101000;
        x_t[30] = 21'b111111111110011100010;
        x_t[31] = 21'b111111111101110101111;
        x_t[32] = 21'b111111111101110101110;
        x_t[33] = 21'b111111111110001101111;
        x_t[34] = 21'b111111111111010011110;
        x_t[35] = 21'b111111111111010001101;
        x_t[36] = 21'b111111111110100000001;
        x_t[37] = 21'b111111111111011100010;
        x_t[38] = 21'b111111111011010101111;
        x_t[39] = 21'b111111111111011001100;
        x_t[40] = 21'b111111111011000111110;
        x_t[41] = 21'b000000000010111101110;
        x_t[42] = 21'b111111111001110111000;
        x_t[43] = 21'b111111111100110111000;
        x_t[44] = 21'b111111111101100001111;
        x_t[45] = 21'b111111111110010011010;
        x_t[46] = 21'b111111111111101101010;
        x_t[47] = 21'b111111111111110111111;
        x_t[48] = 21'b000000000001001010010;
        x_t[49] = 21'b000000000001000001001;
        x_t[50] = 21'b000000000001100010010;
        x_t[51] = 21'b000000000001100111110;
        x_t[52] = 21'b000000000000110101100;
        x_t[53] = 21'b000000000000111011101;
        x_t[54] = 21'b000000000000101001000;
        x_t[55] = 21'b000000000001100100111;
        x_t[56] = 21'b000000000001010111001;
        x_t[57] = 21'b000000000010100100000;
        x_t[58] = 21'b000000000001000101001;
        x_t[59] = 21'b000000000000101010101;
        x_t[60] = 21'b000000000001011111000;
        x_t[61] = 21'b000000000001011110100;
        x_t[62] = 21'b111111111111000100010;
        x_t[63] = 21'b111111111111001111111;
        
        h_t_prev[0] = 21'b111111111100110101000;
        h_t_prev[1] = 21'b111111111110111110000;
        h_t_prev[2] = 21'b111111111110011011101;
        h_t_prev[3] = 21'b000000000000010000111;
        h_t_prev[4] = 21'b000000000000010011010;
        h_t_prev[5] = 21'b000000000000001000100;
        h_t_prev[6] = 21'b111111111110111110100;
        h_t_prev[7] = 21'b111111111110011010110;
        h_t_prev[8] = 21'b111111111110111001011;
        h_t_prev[9] = 21'b111111111111011110110;
        h_t_prev[10] = 21'b000000000000001111010;
        h_t_prev[11] = 21'b000000000001000110100;
        h_t_prev[12] = 21'b000000000001001001100;
        h_t_prev[13] = 21'b111111111111110100011;
        h_t_prev[14] = 21'b111111111101011101000;
        h_t_prev[15] = 21'b111111111110100010000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 74 timeout!");
                $fdisplay(fd_cycles, "Test Vector  74: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  74: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 74");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 75
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111100100001010;
        x_t[1] = 21'b111111111111010001101;
        x_t[2] = 21'b111111111110100000100;
        x_t[3] = 21'b000000000000001100000;
        x_t[4] = 21'b000000000000001001001;
        x_t[5] = 21'b000000000000011110101;
        x_t[6] = 21'b111111111111010001010;
        x_t[7] = 21'b111111111111011100111;
        x_t[8] = 21'b000000000000000001101;
        x_t[9] = 21'b111111111111110010110;
        x_t[10] = 21'b111111111111110110110;
        x_t[11] = 21'b000000000001000110100;
        x_t[12] = 21'b000000000000110010001;
        x_t[13] = 21'b000000000000001000111;
        x_t[14] = 21'b111111111110111100000;
        x_t[15] = 21'b111111111111100100001;
        x_t[16] = 21'b000000000000000001011;
        x_t[17] = 21'b000000000000100001100;
        x_t[18] = 21'b111111111111111101101;
        x_t[19] = 21'b111111111111110100110;
        x_t[20] = 21'b000000000000001110010;
        x_t[21] = 21'b111111111011011011000;
        x_t[22] = 21'b111111111011101000111;
        x_t[23] = 21'b111111111100001110011;
        x_t[24] = 21'b111111111010101001111;
        x_t[25] = 21'b111111111010110000101;
        x_t[26] = 21'b111111111101001110000;
        x_t[27] = 21'b111111111101011000101;
        x_t[28] = 21'b111111111100100111001;
        x_t[29] = 21'b111111111010101111111;
        x_t[30] = 21'b111111111101011101111;
        x_t[31] = 21'b111111111101001101111;
        x_t[32] = 21'b111111111101001000010;
        x_t[33] = 21'b111111111101011111100;
        x_t[34] = 21'b111111111110100100001;
        x_t[35] = 21'b111111111110010110100;
        x_t[36] = 21'b111111111110000111011;
        x_t[37] = 21'b111111111110100111010;
        x_t[38] = 21'b111111111011111001001;
        x_t[39] = 21'b111111111101111010000;
        x_t[40] = 21'b111111111100111001111;
        x_t[41] = 21'b111111111101100010000;
        x_t[42] = 21'b111111111010111000010;
        x_t[43] = 21'b111111111011010100010;
        x_t[44] = 21'b111111111101101101000;
        x_t[45] = 21'b111111111100011111001;
        x_t[46] = 21'b111111111111101101010;
        x_t[47] = 21'b111111111111100100000;
        x_t[48] = 21'b000000000000011010101;
        x_t[49] = 21'b111111111111101001001;
        x_t[50] = 21'b111111111111001111000;
        x_t[51] = 21'b111111111111001101010;
        x_t[52] = 21'b111111111110000111100;
        x_t[53] = 21'b111111111110111011101;
        x_t[54] = 21'b111111111110110001001;
        x_t[55] = 21'b000000000000110101011;
        x_t[56] = 21'b000000000000011011000;
        x_t[57] = 21'b000000000000100100001;
        x_t[58] = 21'b111111111110111001100;
        x_t[59] = 21'b111111111111100011101;
        x_t[60] = 21'b000000000001101010100;
        x_t[61] = 21'b000000000000111001010;
        x_t[62] = 21'b111111111110100110101;
        x_t[63] = 21'b111111111111100101111;
        
        h_t_prev[0] = 21'b111111111100100001010;
        h_t_prev[1] = 21'b111111111111010001101;
        h_t_prev[2] = 21'b111111111110100000100;
        h_t_prev[3] = 21'b000000000000001100000;
        h_t_prev[4] = 21'b000000000000001001001;
        h_t_prev[5] = 21'b000000000000011110101;
        h_t_prev[6] = 21'b111111111111010001010;
        h_t_prev[7] = 21'b111111111111011100111;
        h_t_prev[8] = 21'b000000000000000001101;
        h_t_prev[9] = 21'b111111111111110010110;
        h_t_prev[10] = 21'b111111111111110110110;
        h_t_prev[11] = 21'b000000000001000110100;
        h_t_prev[12] = 21'b000000000000110010001;
        h_t_prev[13] = 21'b000000000000001000111;
        h_t_prev[14] = 21'b111111111110111100000;
        h_t_prev[15] = 21'b111111111111100100001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 75 timeout!");
                $fdisplay(fd_cycles, "Test Vector  75: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  75: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 75");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 76
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111011101011000;
        x_t[1] = 21'b111111111100111110110;
        x_t[2] = 21'b111111111100110101110;
        x_t[3] = 21'b111111111110111001111;
        x_t[4] = 21'b111111111110101110010;
        x_t[5] = 21'b111111111110010100000;
        x_t[6] = 21'b111111111101010100110;
        x_t[7] = 21'b111111111101100010110;
        x_t[8] = 21'b111111111110000101111;
        x_t[9] = 21'b111111111101110000100;
        x_t[10] = 21'b111111111101110111101;
        x_t[11] = 21'b111111111111010001010;
        x_t[12] = 21'b111111111110011001111;
        x_t[13] = 21'b111111111101001010001;
        x_t[14] = 21'b111111111101110010001;
        x_t[15] = 21'b111111111101111110011;
        x_t[16] = 21'b111111111110001010100;
        x_t[17] = 21'b111111111110001000100;
        x_t[18] = 21'b111111111101100100110;
        x_t[19] = 21'b111111111101110000111;
        x_t[20] = 21'b111111111101111110011;
        x_t[21] = 21'b111111111011010101100;
        x_t[22] = 21'b111111111011100010100;
        x_t[23] = 21'b111111111100001011011;
        x_t[24] = 21'b111111111010101100111;
        x_t[25] = 21'b111111111010110000101;
        x_t[26] = 21'b111111111101001110000;
        x_t[27] = 21'b111111111100111101001;
        x_t[28] = 21'b111111111100010001001;
        x_t[29] = 21'b111111111011001000110;
        x_t[30] = 21'b111111111101100001110;
        x_t[31] = 21'b111111111100101110111;
        x_t[32] = 21'b111111111101010001011;
        x_t[33] = 21'b111111111101110110110;
        x_t[34] = 21'b111111111110101101101;
        x_t[35] = 21'b111111111110010110100;
        x_t[36] = 21'b111111111101011111101;
        x_t[37] = 21'b111111111110000110101;
        x_t[38] = 21'b111111111101101000000;
        x_t[39] = 21'b111111111101001101111;
        x_t[40] = 21'b111111111110100001001;
        x_t[41] = 21'b111111111100001110100;
        x_t[42] = 21'b111111111101001100100;
        x_t[43] = 21'b111111111100110111000;
        x_t[44] = 21'b111111111101111101111;
        x_t[45] = 21'b111111111101011101000;
        x_t[46] = 21'b000000000000000111001;
        x_t[47] = 21'b111111111111110010111;
        x_t[48] = 21'b000000000000010001001;
        x_t[49] = 21'b111111111111001101010;
        x_t[50] = 21'b111111111110101101110;
        x_t[51] = 21'b111111111110110000010;
        x_t[52] = 21'b111111111110001100101;
        x_t[53] = 21'b111111111111101000001;
        x_t[54] = 21'b111111111111111111000;
        x_t[55] = 21'b000000000001011100010;
        x_t[56] = 21'b000000000000111101011;
        x_t[57] = 21'b000000000000011111111;
        x_t[58] = 21'b111111111111010011110;
        x_t[59] = 21'b000000000000101110101;
        x_t[60] = 21'b000000000001011111000;
        x_t[61] = 21'b000000000000110001000;
        x_t[62] = 21'b111111111110111001001;
        x_t[63] = 21'b000000000000111001100;
        
        h_t_prev[0] = 21'b111111111011101011000;
        h_t_prev[1] = 21'b111111111100111110110;
        h_t_prev[2] = 21'b111111111100110101110;
        h_t_prev[3] = 21'b111111111110111001111;
        h_t_prev[4] = 21'b111111111110101110010;
        h_t_prev[5] = 21'b111111111110010100000;
        h_t_prev[6] = 21'b111111111101010100110;
        h_t_prev[7] = 21'b111111111101100010110;
        h_t_prev[8] = 21'b111111111110000101111;
        h_t_prev[9] = 21'b111111111101110000100;
        h_t_prev[10] = 21'b111111111101110111101;
        h_t_prev[11] = 21'b111111111111010001010;
        h_t_prev[12] = 21'b111111111110011001111;
        h_t_prev[13] = 21'b111111111101001010001;
        h_t_prev[14] = 21'b111111111101110010001;
        h_t_prev[15] = 21'b111111111101111110011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 76 timeout!");
                $fdisplay(fd_cycles, "Test Vector  76: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  76: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 76");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 77
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111110001000111;
        x_t[1] = 21'b111111111111010110100;
        x_t[2] = 21'b111111111111000010100;
        x_t[3] = 21'b000000000000110111100;
        x_t[4] = 21'b000000000000110001100;
        x_t[5] = 21'b000000000000001000100;
        x_t[6] = 21'b111111111110101011111;
        x_t[7] = 21'b000000000001010111001;
        x_t[8] = 21'b000000000000110000000;
        x_t[9] = 21'b000000000000000001111;
        x_t[10] = 21'b000000000000001010011;
        x_t[11] = 21'b000000000001101010001;
        x_t[12] = 21'b000000000000100000100;
        x_t[13] = 21'b111111111111001011100;
        x_t[14] = 21'b000000000000010101101;
        x_t[15] = 21'b000000000000100110010;
        x_t[16] = 21'b000000000000010000010;
        x_t[17] = 21'b000000000000010010101;
        x_t[18] = 21'b111111111111100011010;
        x_t[19] = 21'b111111111111110100110;
        x_t[20] = 21'b000000000000100001000;
        x_t[21] = 21'b111111111100011010100;
        x_t[22] = 21'b111111111100100101001;
        x_t[23] = 21'b111111111100111001111;
        x_t[24] = 21'b111111111100010001011;
        x_t[25] = 21'b111111111100010001000;
        x_t[26] = 21'b111111111110101010111;
        x_t[27] = 21'b111111111110001111101;
        x_t[28] = 21'b111111111100110110111;
        x_t[29] = 21'b111111111101000101101;
        x_t[30] = 21'b000000000000000001110;
        x_t[31] = 21'b111111111110101111100;
        x_t[32] = 21'b111111111110111001111;
        x_t[33] = 21'b111111111111001110101;
        x_t[34] = 21'b000000000000010110011;
        x_t[35] = 21'b111111111111111001001;
        x_t[36] = 21'b111111111110111001000;
        x_t[37] = 21'b111111111111001011111;
        x_t[38] = 21'b111111111111100001001;
        x_t[39] = 21'b111111111101101011010;
        x_t[40] = 21'b000000000000001101111;
        x_t[41] = 21'b111111111101111101110;
        x_t[42] = 21'b111111111101000000101;
        x_t[43] = 21'b111111111111100110101;
        x_t[44] = 21'b111111111111111110010;
        x_t[45] = 21'b111111111110010011010;
        x_t[46] = 21'b000000000001010100111;
        x_t[47] = 21'b000000000000111101100;
        x_t[48] = 21'b000000000001011101011;
        x_t[49] = 21'b000000000000000100111;
        x_t[50] = 21'b111111111111010011110;
        x_t[51] = 21'b111111111110111110110;
        x_t[52] = 21'b111111111110010001110;
        x_t[53] = 21'b111111111111010111011;
        x_t[54] = 21'b111111111111100111001;
        x_t[55] = 21'b000000000001110001110;
        x_t[56] = 21'b000000000001001110100;
        x_t[57] = 21'b000000000000001110111;
        x_t[58] = 21'b111111111110110000111;
        x_t[59] = 21'b111111111111010011111;
        x_t[60] = 21'b000000000001101110011;
        x_t[61] = 21'b000000000001010010001;
        x_t[62] = 21'b111111111110110101011;
        x_t[63] = 21'b000000000010001101001;
        
        h_t_prev[0] = 21'b111111111110001000111;
        h_t_prev[1] = 21'b111111111111010110100;
        h_t_prev[2] = 21'b111111111111000010100;
        h_t_prev[3] = 21'b000000000000110111100;
        h_t_prev[4] = 21'b000000000000110001100;
        h_t_prev[5] = 21'b000000000000001000100;
        h_t_prev[6] = 21'b111111111110101011111;
        h_t_prev[7] = 21'b000000000001010111001;
        h_t_prev[8] = 21'b000000000000110000000;
        h_t_prev[9] = 21'b000000000000000001111;
        h_t_prev[10] = 21'b000000000000001010011;
        h_t_prev[11] = 21'b000000000001101010001;
        h_t_prev[12] = 21'b000000000000100000100;
        h_t_prev[13] = 21'b111111111111001011100;
        h_t_prev[14] = 21'b000000000000010101101;
        h_t_prev[15] = 21'b000000000000100110010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 77 timeout!");
                $fdisplay(fd_cycles, "Test Vector  77: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  77: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 77");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 78
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111110100110100;
        x_t[1] = 21'b111111111111010110100;
        x_t[2] = 21'b111111111110100000100;
        x_t[3] = 21'b111111111111111000110;
        x_t[4] = 21'b111111111111100101110;
        x_t[5] = 21'b111111111111001011100;
        x_t[6] = 21'b111111111101110011111;
        x_t[7] = 21'b000000000000011111001;
        x_t[8] = 21'b111111111111110111011;
        x_t[9] = 21'b111111111111000101110;
        x_t[10] = 21'b111111111110110111010;
        x_t[11] = 21'b111111111111101010110;
        x_t[12] = 21'b111111111110001000011;
        x_t[13] = 21'b111111111101001010001;
        x_t[14] = 21'b111111111110100001101;
        x_t[15] = 21'b111111111111000000100;
        x_t[16] = 21'b111111111110101000010;
        x_t[17] = 21'b111111111110100110001;
        x_t[18] = 21'b111111111101010101000;
        x_t[19] = 21'b111111111101001010100;
        x_t[20] = 21'b111111111101010010101;
        x_t[21] = 21'b111111111011101110011;
        x_t[22] = 21'b111111111011111011111;
        x_t[23] = 21'b111111111100000010110;
        x_t[24] = 21'b111111111011010111100;
        x_t[25] = 21'b111111111011011100001;
        x_t[26] = 21'b111111111101001110000;
        x_t[27] = 21'b111111111101000101000;
        x_t[28] = 21'b111111111100000001011;
        x_t[29] = 21'b111111111011001000110;
        x_t[30] = 21'b111111111111100110011;
        x_t[31] = 21'b111111111101000000101;
        x_t[32] = 21'b111111111101000011110;
        x_t[33] = 21'b111111111101001000011;
        x_t[34] = 21'b111111111110010101110;
        x_t[35] = 21'b111111111110000010110;
        x_t[36] = 21'b111111111101000110110;
        x_t[37] = 21'b111111111101010101101;
        x_t[38] = 21'b111111111100011100011;
        x_t[39] = 21'b111111111011101110011;
        x_t[40] = 21'b111111111100011110110;
        x_t[41] = 21'b111111111101100010000;
        x_t[42] = 21'b111111111001011001011;
        x_t[43] = 21'b111111111011101010010;
        x_t[44] = 21'b111111111101001011100;
        x_t[45] = 21'b111111111001011101110;
        x_t[46] = 21'b111111111110010000000;
        x_t[47] = 21'b111111111101101100101;
        x_t[48] = 21'b111111111110000010001;
        x_t[49] = 21'b111111111100111001000;
        x_t[50] = 21'b111111111100010101101;
        x_t[51] = 21'b111111111100000010011;
        x_t[52] = 21'b111111111011001010010;
        x_t[53] = 21'b111111111011111000110;
        x_t[54] = 21'b111111111011011111011;
        x_t[55] = 21'b111111111111001001100;
        x_t[56] = 21'b111111111110101111100;
        x_t[57] = 21'b111111111101101100111;
        x_t[58] = 21'b111111111100011000001;
        x_t[59] = 21'b111111111100100110001;
        x_t[60] = 21'b000000000000110100111;
        x_t[61] = 21'b111111111111111011010;
        x_t[62] = 21'b111111111100110000010;
        x_t[63] = 21'b000000000000110000101;
        
        h_t_prev[0] = 21'b111111111110100110100;
        h_t_prev[1] = 21'b111111111111010110100;
        h_t_prev[2] = 21'b111111111110100000100;
        h_t_prev[3] = 21'b111111111111111000110;
        h_t_prev[4] = 21'b111111111111100101110;
        h_t_prev[5] = 21'b111111111111001011100;
        h_t_prev[6] = 21'b111111111101110011111;
        h_t_prev[7] = 21'b000000000000011111001;
        h_t_prev[8] = 21'b111111111111110111011;
        h_t_prev[9] = 21'b111111111111000101110;
        h_t_prev[10] = 21'b111111111110110111010;
        h_t_prev[11] = 21'b111111111111101010110;
        h_t_prev[12] = 21'b111111111110001000011;
        h_t_prev[13] = 21'b111111111101001010001;
        h_t_prev[14] = 21'b111111111110100001101;
        h_t_prev[15] = 21'b111111111111000000100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 78 timeout!");
                $fdisplay(fd_cycles, "Test Vector  78: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  78: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 78");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 79
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111101001000110;
        x_t[1] = 21'b111111111110010010000;
        x_t[2] = 21'b111111111101100110010;
        x_t[3] = 21'b111111111110100001110;
        x_t[4] = 21'b111111111110101001001;
        x_t[5] = 21'b111111111110011001100;
        x_t[6] = 21'b111111111101110011111;
        x_t[7] = 21'b111111111101111100010;
        x_t[8] = 21'b111111111110000101111;
        x_t[9] = 21'b111111111101111010100;
        x_t[10] = 21'b111111111101101000111;
        x_t[11] = 21'b111111111110110111110;
        x_t[12] = 21'b111111111101011111011;
        x_t[13] = 21'b111111111101001010001;
        x_t[14] = 21'b111111111100111000001;
        x_t[15] = 21'b111111111101001011101;
        x_t[16] = 21'b111111111101001111000;
        x_t[17] = 21'b111111111101010111001;
        x_t[18] = 21'b111111111100110101011;
        x_t[19] = 21'b111111111100111010000;
        x_t[20] = 21'b111111111101000110001;
        x_t[21] = 21'b111111111011111001011;
        x_t[22] = 21'b111111111011111111000;
        x_t[23] = 21'b111111111100000101101;
        x_t[24] = 21'b111111111011101100110;
        x_t[25] = 21'b111111111011101000100;
        x_t[26] = 21'b111111111101110100000;
        x_t[27] = 21'b111111111101011100100;
        x_t[28] = 21'b111111111100000001011;
        x_t[29] = 21'b111111111011111110111;
        x_t[30] = 21'b111111111111001111000;
        x_t[31] = 21'b111111111101011011010;
        x_t[32] = 21'b111111111101111110110;
        x_t[33] = 21'b111111111110010010100;
        x_t[34] = 21'b111111111111000101011;
        x_t[35] = 21'b111111111110101111001;
        x_t[36] = 21'b111111111101111000011;
        x_t[37] = 21'b111111111110000110101;
        x_t[38] = 21'b111111111101011000111;
        x_t[39] = 21'b111111111110011110110;
        x_t[40] = 21'b111111111110011011110;
        x_t[41] = 21'b000000000001011100011;
        x_t[42] = 21'b111111111010001110110;
        x_t[43] = 21'b111111111001111100100;
        x_t[44] = 21'b111111111101010110110;
        x_t[45] = 21'b111111111011001010000;
        x_t[46] = 21'b111111111110101001111;
        x_t[47] = 21'b111111111101110001101;
        x_t[48] = 21'b111111111110000110111;
        x_t[49] = 21'b111111111101011110001;
        x_t[50] = 21'b111111111101011000001;
        x_t[51] = 21'b111111111101111111111;
        x_t[52] = 21'b111111111101001010001;
        x_t[53] = 21'b111111111101110011010;
        x_t[54] = 21'b111111111101010111010;
        x_t[55] = 21'b111111111111100011011;
        x_t[56] = 21'b111111111111001001011;
        x_t[57] = 21'b111111111111001010101;
        x_t[58] = 21'b111111111110101100100;
        x_t[59] = 21'b111111111110101100011;
        x_t[60] = 21'b111111111111110111100;
        x_t[61] = 21'b111111111110110100111;
        x_t[62] = 21'b111111111011111000110;
        x_t[63] = 21'b111111111111011000101;
        
        h_t_prev[0] = 21'b111111111101001000110;
        h_t_prev[1] = 21'b111111111110010010000;
        h_t_prev[2] = 21'b111111111101100110010;
        h_t_prev[3] = 21'b111111111110100001110;
        h_t_prev[4] = 21'b111111111110101001001;
        h_t_prev[5] = 21'b111111111110011001100;
        h_t_prev[6] = 21'b111111111101110011111;
        h_t_prev[7] = 21'b111111111101111100010;
        h_t_prev[8] = 21'b111111111110000101111;
        h_t_prev[9] = 21'b111111111101111010100;
        h_t_prev[10] = 21'b111111111101101000111;
        h_t_prev[11] = 21'b111111111110110111110;
        h_t_prev[12] = 21'b111111111101011111011;
        h_t_prev[13] = 21'b111111111101001010001;
        h_t_prev[14] = 21'b111111111100111000001;
        h_t_prev[15] = 21'b111111111101001011101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 79 timeout!");
                $fdisplay(fd_cycles, "Test Vector  79: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  79: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 79");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 80
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111101010111100;
        x_t[1] = 21'b111111111110101111011;
        x_t[2] = 21'b111111111110100000100;
        x_t[3] = 21'b111111111111101010010;
        x_t[4] = 21'b111111111111110100111;
        x_t[5] = 21'b000000000000000011000;
        x_t[6] = 21'b111111111110101011111;
        x_t[7] = 21'b111111111110111110011;
        x_t[8] = 21'b111111111110100100110;
        x_t[9] = 21'b111111111110100010101;
        x_t[10] = 21'b111111111110101000100;
        x_t[11] = 21'b000000000000001001011;
        x_t[12] = 21'b111111111111010100011;
        x_t[13] = 21'b111111111110111101111;
        x_t[14] = 21'b111111111101010111110;
        x_t[15] = 21'b111111111101100101000;
        x_t[16] = 21'b111111111110001111011;
        x_t[17] = 21'b111111111110001101011;
        x_t[18] = 21'b111111111110100100000;
        x_t[19] = 21'b111111111110111101110;
        x_t[20] = 21'b111111111111000011010;
        x_t[21] = 21'b111111111100000001101;
        x_t[22] = 21'b111111111011110010011;
        x_t[23] = 21'b111111111100000010110;
        x_t[24] = 21'b111111111011101111111;
        x_t[25] = 21'b111111111011110101000;
        x_t[26] = 21'b111111111101100111011;
        x_t[27] = 21'b111111111101001100110;
        x_t[28] = 21'b111111111011110111111;
        x_t[29] = 21'b111111111100011100000;
        x_t[30] = 21'b111111111110100100001;
        x_t[31] = 21'b111111111101110001011;
        x_t[32] = 21'b111111111101111010010;
        x_t[33] = 21'b111111111110010111001;
        x_t[34] = 21'b111111111111001010001;
        x_t[35] = 21'b111111111110100000011;
        x_t[36] = 21'b111111111101101110100;
        x_t[37] = 21'b111111111110001010101;
        x_t[38] = 21'b111111111101100011000;
        x_t[39] = 21'b111111111110110100110;
        x_t[40] = 21'b111111111011010010101;
        x_t[41] = 21'b111111111111010001010;
        x_t[42] = 21'b111111111001110111000;
        x_t[43] = 21'b111111111110111010110;
        x_t[44] = 21'b111111111101000110000;
        x_t[45] = 21'b111111111101100100110;
        x_t[46] = 21'b111111111110001010110;
        x_t[47] = 21'b111111111101101100101;
        x_t[48] = 21'b111111111110001011110;
        x_t[49] = 21'b111111111110010101110;
        x_t[50] = 21'b111111111110101001000;
        x_t[51] = 21'b111111111111110011111;
        x_t[52] = 21'b111111111111001111001;
        x_t[53] = 21'b111111111111101101110;
        x_t[54] = 21'b111111111111011011001;
        x_t[55] = 21'b111111111111000000111;
        x_t[56] = 21'b111111111110101011010;
        x_t[57] = 21'b000000000000001010101;
        x_t[58] = 21'b000000000000100010010;
        x_t[59] = 21'b000000000000011110111;
        x_t[60] = 21'b111111111111100000100;
        x_t[61] = 21'b111111111111010001111;
        x_t[62] = 21'b111111111101011001000;
        x_t[63] = 21'b111111111111101110101;
        
        h_t_prev[0] = 21'b111111111101010111100;
        h_t_prev[1] = 21'b111111111110101111011;
        h_t_prev[2] = 21'b111111111110100000100;
        h_t_prev[3] = 21'b111111111111101010010;
        h_t_prev[4] = 21'b111111111111110100111;
        h_t_prev[5] = 21'b000000000000000011000;
        h_t_prev[6] = 21'b111111111110101011111;
        h_t_prev[7] = 21'b111111111110111110011;
        h_t_prev[8] = 21'b111111111110100100110;
        h_t_prev[9] = 21'b111111111110100010101;
        h_t_prev[10] = 21'b111111111110101000100;
        h_t_prev[11] = 21'b000000000000001001011;
        h_t_prev[12] = 21'b111111111111010100011;
        h_t_prev[13] = 21'b111111111110111101111;
        h_t_prev[14] = 21'b111111111101010111110;
        h_t_prev[15] = 21'b111111111101100101000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 80 timeout!");
                $fdisplay(fd_cycles, "Test Vector  80: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  80: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 80");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 81
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000001110000110;
        x_t[1] = 21'b000000000001110011001;
        x_t[2] = 21'b000000000000101101011;
        x_t[3] = 21'b000000000001100011000;
        x_t[4] = 21'b000000000001111101011;
        x_t[5] = 21'b000000000000111010011;
        x_t[6] = 21'b000000000000111011000;
        x_t[7] = 21'b000000000000011010000;
        x_t[8] = 21'b000000000001001111000;
        x_t[9] = 21'b000000000001100001000;
        x_t[10] = 21'b000000000010001001101;
        x_t[11] = 21'b000000000000001110100;
        x_t[12] = 21'b000000000001011011000;
        x_t[13] = 21'b000000000010000011100;
        x_t[14] = 21'b000000000001011010001;
        x_t[15] = 21'b000000000001011110001;
        x_t[16] = 21'b000000000001100100100;
        x_t[17] = 21'b000000000001010111110;
        x_t[18] = 21'b000000000001010111010;
        x_t[19] = 21'b000000000001111110000;
        x_t[20] = 21'b000000000001000000011;
        x_t[21] = 21'b000000000000100011110;
        x_t[22] = 21'b000000000000101111101;
        x_t[23] = 21'b111111111111011111001;
        x_t[24] = 21'b111111111111010100010;
        x_t[25] = 21'b111111111111011110001;
        x_t[26] = 21'b111111111111011101101;
        x_t[27] = 21'b111111111111101010000;
        x_t[28] = 21'b000000000000011111111;
        x_t[29] = 21'b000000000000110010101;
        x_t[30] = 21'b111111111111100010100;
        x_t[31] = 21'b111111111110101111100;
        x_t[32] = 21'b111111111111100111010;
        x_t[33] = 21'b111111111111010111111;
        x_t[34] = 21'b111111111111000000101;
        x_t[35] = 21'b111111111111010110101;
        x_t[36] = 21'b111111111111011011111;
        x_t[37] = 21'b000000000000111110000;
        x_t[38] = 21'b111111111111100001001;
        x_t[39] = 21'b000000000001011101110;
        x_t[40] = 21'b111111111111111000001;
        x_t[41] = 21'b111111111101111101110;
        x_t[42] = 21'b111111111111010100111;
        x_t[43] = 21'b000000000011101101111;
        x_t[44] = 21'b111111111110001001000;
        x_t[45] = 21'b000000000010101001110;
        x_t[46] = 21'b000000000001000000001;
        x_t[47] = 21'b000000000000111000100;
        x_t[48] = 21'b000000000001000101100;
        x_t[49] = 21'b000000000001000001001;
        x_t[50] = 21'b000000000001101011110;
        x_t[51] = 21'b000000000001111011001;
        x_t[52] = 21'b000000000001101000101;
        x_t[53] = 21'b000000000001010111100;
        x_t[54] = 21'b000000000000111011000;
        x_t[55] = 21'b000000000001010011101;
        x_t[56] = 21'b000000000000111001000;
        x_t[57] = 21'b000000000010010011000;
        x_t[58] = 21'b000000000010101001100;
        x_t[59] = 21'b000000000010110100111;
        x_t[60] = 21'b000000000010110111001;
        x_t[61] = 21'b000000000100100101010;
        x_t[62] = 21'b000000000010010011011;
        x_t[63] = 21'b000000000001111011100;
        
        h_t_prev[0] = 21'b000000000001110000110;
        h_t_prev[1] = 21'b000000000001110011001;
        h_t_prev[2] = 21'b000000000000101101011;
        h_t_prev[3] = 21'b000000000001100011000;
        h_t_prev[4] = 21'b000000000001111101011;
        h_t_prev[5] = 21'b000000000000111010011;
        h_t_prev[6] = 21'b000000000000111011000;
        h_t_prev[7] = 21'b000000000000011010000;
        h_t_prev[8] = 21'b000000000001001111000;
        h_t_prev[9] = 21'b000000000001100001000;
        h_t_prev[10] = 21'b000000000010001001101;
        h_t_prev[11] = 21'b000000000000001110100;
        h_t_prev[12] = 21'b000000000001011011000;
        h_t_prev[13] = 21'b000000000010000011100;
        h_t_prev[14] = 21'b000000000001011010001;
        h_t_prev[15] = 21'b000000000001011110001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 81 timeout!");
                $fdisplay(fd_cycles, "Test Vector  81: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  81: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 81");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 82
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000000100110110;
        x_t[1] = 21'b000000000000110011100;
        x_t[2] = 21'b000000000000000110100;
        x_t[3] = 21'b000000000001001111110;
        x_t[4] = 21'b000000000001100100001;
        x_t[5] = 21'b000000000000000011000;
        x_t[6] = 21'b111111111111110000011;
        x_t[7] = 21'b111111111111010111111;
        x_t[8] = 21'b000000000000011011011;
        x_t[9] = 21'b000000000001001000000;
        x_t[10] = 21'b000000000001100111011;
        x_t[11] = 21'b000000000000011000101;
        x_t[12] = 21'b000000000000110010001;
        x_t[13] = 21'b000000000000111000101;
        x_t[14] = 21'b000000000000110000000;
        x_t[15] = 21'b000000000000011100001;
        x_t[16] = 21'b000000000000101110000;
        x_t[17] = 21'b000000000000110000010;
        x_t[18] = 21'b000000000000111100111;
        x_t[19] = 21'b000000000001010111101;
        x_t[20] = 21'b000000000000001110010;
        x_t[21] = 21'b000000000000111001111;
        x_t[22] = 21'b000000000001000101111;
        x_t[23] = 21'b000000000000000010000;
        x_t[24] = 21'b111111111111100000011;
        x_t[25] = 21'b111111111111100100010;
        x_t[26] = 21'b000000000000000011101;
        x_t[27] = 21'b000000000000000101100;
        x_t[28] = 21'b000000000000110010110;
        x_t[29] = 21'b000000000000010101100;
        x_t[30] = 21'b111111111111011110101;
        x_t[31] = 21'b111111111111000001010;
        x_t[32] = 21'b000000000000001011101;
        x_t[33] = 21'b000000000000001010110;
        x_t[34] = 21'b111111111111100110110;
        x_t[35] = 21'b111111111111100101011;
        x_t[36] = 21'b111111111111000011000;
        x_t[37] = 21'b000000000000101101110;
        x_t[38] = 21'b111111111111000111111;
        x_t[39] = 21'b111111111111111110010;
        x_t[40] = 21'b000000000000000011000;
        x_t[41] = 21'b111111111011010000000;
        x_t[42] = 21'b111111111101101010001;
        x_t[43] = 21'b000000000010000000001;
        x_t[44] = 21'b111111111101011100010;
        x_t[45] = 21'b000000000100000110101;
        x_t[46] = 21'b000000000000011011111;
        x_t[47] = 21'b000000000000011010101;
        x_t[48] = 21'b000000000000110111010;
        x_t[49] = 21'b000000000001000001001;
        x_t[50] = 21'b000000000001011000110;
        x_t[51] = 21'b000000000001111011001;
        x_t[52] = 21'b000000000001100011100;
        x_t[53] = 21'b000000000001011101000;
        x_t[54] = 21'b000000000001101010111;
        x_t[55] = 21'b000000000001001011000;
        x_t[56] = 21'b000000000000110000100;
        x_t[57] = 21'b000000000010000110010;
        x_t[58] = 21'b000000000010010011101;
        x_t[59] = 21'b000000000011000000101;
        x_t[60] = 21'b000000000010111011000;
        x_t[61] = 21'b000000000100000000000;
        x_t[62] = 21'b000000000001001101001;
        x_t[63] = 21'b000000000010001101001;
        
        h_t_prev[0] = 21'b000000000000100110110;
        h_t_prev[1] = 21'b000000000000110011100;
        h_t_prev[2] = 21'b000000000000000110100;
        h_t_prev[3] = 21'b000000000001001111110;
        h_t_prev[4] = 21'b000000000001100100001;
        h_t_prev[5] = 21'b000000000000000011000;
        h_t_prev[6] = 21'b111111111111110000011;
        h_t_prev[7] = 21'b111111111111010111111;
        h_t_prev[8] = 21'b000000000000011011011;
        h_t_prev[9] = 21'b000000000001001000000;
        h_t_prev[10] = 21'b000000000001100111011;
        h_t_prev[11] = 21'b000000000000011000101;
        h_t_prev[12] = 21'b000000000000110010001;
        h_t_prev[13] = 21'b000000000000111000101;
        h_t_prev[14] = 21'b000000000000110000000;
        h_t_prev[15] = 21'b000000000000011100001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 82 timeout!");
                $fdisplay(fd_cycles, "Test Vector  82: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  82: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 82");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 83
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111111010111110;
        x_t[1] = 21'b000000000000000010100;
        x_t[2] = 21'b000000000000000001101;
        x_t[3] = 21'b000000000001100011000;
        x_t[4] = 21'b000000000001101110001;
        x_t[5] = 21'b000000000000000011000;
        x_t[6] = 21'b111111111111010001010;
        x_t[7] = 21'b111111111101110111001;
        x_t[8] = 21'b111111111111001110000;
        x_t[9] = 21'b000000000000101001111;
        x_t[10] = 21'b000000000001111010111;
        x_t[11] = 21'b111111111111111111001;
        x_t[12] = 21'b000000000000011010101;
        x_t[13] = 21'b000000000000110001110;
        x_t[14] = 21'b111111111110110110110;
        x_t[15] = 21'b111111111111110011011;
        x_t[16] = 21'b000000000000010000010;
        x_t[17] = 21'b000000000000011100100;
        x_t[18] = 21'b000000000000011101010;
        x_t[19] = 21'b000000000000101011101;
        x_t[20] = 21'b111111111111110101010;
        x_t[21] = 21'b111111111111100111000;
        x_t[22] = 21'b111111111111101101000;
        x_t[23] = 21'b111111111110111100011;
        x_t[24] = 21'b111111111101100110101;
        x_t[25] = 21'b111111111101110001010;
        x_t[26] = 21'b111111111110100010100;
        x_t[27] = 21'b111111111110101011001;
        x_t[28] = 21'b111111111111110000101;
        x_t[29] = 21'b111111111110001100010;
        x_t[30] = 21'b111111111101001010011;
        x_t[31] = 21'b111111111101101101000;
        x_t[32] = 21'b111111111110010101100;
        x_t[33] = 21'b111111111110100101000;
        x_t[34] = 21'b111111111101111110000;
        x_t[35] = 21'b111111111101101111000;
        x_t[36] = 21'b111111111101000001110;
        x_t[37] = 21'b111111111111000011110;
        x_t[38] = 21'b111111111100111010101;
        x_t[39] = 21'b111111111111010010001;
        x_t[40] = 21'b111111111100100100001;
        x_t[41] = 21'b111111111100100011011;
        x_t[42] = 21'b111111111100010001010;
        x_t[43] = 21'b111111111111110001100;
        x_t[44] = 21'b111111111100000010111;
        x_t[45] = 21'b000000000011110111001;
        x_t[46] = 21'b111111111110111110101;
        x_t[47] = 21'b111111111111100100000;
        x_t[48] = 21'b111111111111111110000;
        x_t[49] = 21'b000000000000010010110;
        x_t[50] = 21'b000000000000010110010;
        x_t[51] = 21'b000000000000100100001;
        x_t[52] = 21'b000000000000010001101;
        x_t[53] = 21'b000000000000100101011;
        x_t[54] = 21'b000000000001101010111;
        x_t[55] = 21'b000000000001010011101;
        x_t[56] = 21'b000000000000011011000;
        x_t[57] = 21'b000000000001001010100;
        x_t[58] = 21'b000000000001010110101;
        x_t[59] = 21'b000000000010111100110;
        x_t[60] = 21'b000000000010100111111;
        x_t[61] = 21'b000000000011100011000;
        x_t[62] = 21'b000000000000010001111;
        x_t[63] = 21'b000000000010001000110;
        
        h_t_prev[0] = 21'b111111111111010111110;
        h_t_prev[1] = 21'b000000000000000010100;
        h_t_prev[2] = 21'b000000000000000001101;
        h_t_prev[3] = 21'b000000000001100011000;
        h_t_prev[4] = 21'b000000000001101110001;
        h_t_prev[5] = 21'b000000000000000011000;
        h_t_prev[6] = 21'b111111111111010001010;
        h_t_prev[7] = 21'b111111111101110111001;
        h_t_prev[8] = 21'b111111111111001110000;
        h_t_prev[9] = 21'b000000000000101001111;
        h_t_prev[10] = 21'b000000000001111010111;
        h_t_prev[11] = 21'b111111111111111111001;
        h_t_prev[12] = 21'b000000000000011010101;
        h_t_prev[13] = 21'b000000000000110001110;
        h_t_prev[14] = 21'b111111111110110110110;
        h_t_prev[15] = 21'b111111111111110011011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 83 timeout!");
                $fdisplay(fd_cycles, "Test Vector  83: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  83: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 83");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 84
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111101101011010;
        x_t[1] = 21'b111111111110011011110;
        x_t[2] = 21'b111111111110001101001;
        x_t[3] = 21'b111111111111100000100;
        x_t[4] = 21'b111111111111101111111;
        x_t[5] = 21'b111111111110000011011;
        x_t[6] = 21'b111111111101001000010;
        x_t[7] = 21'b111111111100000111001;
        x_t[8] = 21'b111111111110000000110;
        x_t[9] = 21'b111111111111001111110;
        x_t[10] = 21'b000000000000011101111;
        x_t[11] = 21'b111111111101110000100;
        x_t[12] = 21'b111111111110100101101;
        x_t[13] = 21'b111111111111101101101;
        x_t[14] = 21'b111111111110110110110;
        x_t[15] = 21'b111111111111100100001;
        x_t[16] = 21'b111111111111011001110;
        x_t[17] = 21'b111111111111010010100;
        x_t[18] = 21'b111111111110101110100;
        x_t[19] = 21'b111111111110111101110;
        x_t[20] = 21'b111111111110010111011;
        x_t[21] = 21'b111111111111010000111;
        x_t[22] = 21'b111111111111000011110;
        x_t[23] = 21'b111111111110000101010;
        x_t[24] = 21'b111111111101100011100;
        x_t[25] = 21'b111111111101011110101;
        x_t[26] = 21'b111111111101110100000;
        x_t[27] = 21'b111111111101101000011;
        x_t[28] = 21'b111111111110101011011;
        x_t[29] = 21'b111111111110011100111;
        x_t[30] = 21'b111111111101010110000;
        x_t[31] = 21'b111111111100101010011;
        x_t[32] = 21'b111111111110000011011;
        x_t[33] = 21'b111111111101110010001;
        x_t[34] = 21'b111111111101000100111;
        x_t[35] = 21'b111111111101010110011;
        x_t[36] = 21'b111111111100010000000;
        x_t[37] = 21'b111111111110001110110;
        x_t[38] = 21'b111111111101111100010;
        x_t[39] = 21'b000000000000010100010;
        x_t[40] = 21'b111111111111010111100;
        x_t[41] = 21'b111111111111100110001;
        x_t[42] = 21'b111111111110001101110;
        x_t[43] = 21'b111111111101100010111;
        x_t[44] = 21'b111111111101010001001;
        x_t[45] = 21'b000000000001110011101;
        x_t[46] = 21'b000000000000010001100;
        x_t[47] = 21'b000000000000001011110;
        x_t[48] = 21'b111111111111100001100;
        x_t[49] = 21'b111111111111110111000;
        x_t[50] = 21'b111111111111000101100;
        x_t[51] = 21'b111111111110111110110;
        x_t[52] = 21'b111111111110100001001;
        x_t[53] = 21'b111111111110111011101;
        x_t[54] = 21'b000000000000110101000;
        x_t[55] = 21'b000000000001101101100;
        x_t[56] = 21'b000000000000010010011;
        x_t[57] = 21'b111111111111110101010;
        x_t[58] = 21'b000000000000010101001;
        x_t[59] = 21'b000000000011000000101;
        x_t[60] = 21'b000000000010100111111;
        x_t[61] = 21'b000000000011010010011;
        x_t[62] = 21'b111111111111111111011;
        x_t[63] = 21'b000000000010000100010;
        
        h_t_prev[0] = 21'b111111111101101011010;
        h_t_prev[1] = 21'b111111111110011011110;
        h_t_prev[2] = 21'b111111111110001101001;
        h_t_prev[3] = 21'b111111111111100000100;
        h_t_prev[4] = 21'b111111111111101111111;
        h_t_prev[5] = 21'b111111111110000011011;
        h_t_prev[6] = 21'b111111111101001000010;
        h_t_prev[7] = 21'b111111111100000111001;
        h_t_prev[8] = 21'b111111111110000000110;
        h_t_prev[9] = 21'b111111111111001111110;
        h_t_prev[10] = 21'b000000000000011101111;
        h_t_prev[11] = 21'b111111111101110000100;
        h_t_prev[12] = 21'b111111111110100101101;
        h_t_prev[13] = 21'b111111111111101101101;
        h_t_prev[14] = 21'b111111111110110110110;
        h_t_prev[15] = 21'b111111111111100100001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 84 timeout!");
                $fdisplay(fd_cycles, "Test Vector  84: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  84: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 84");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 85
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111110100110100;
        x_t[1] = 21'b111111111111001100110;
        x_t[2] = 21'b111111111110000011011;
        x_t[3] = 21'b111111111110110000010;
        x_t[4] = 21'b111111111110110011010;
        x_t[5] = 21'b111111111101010111000;
        x_t[6] = 21'b111111111101010100110;
        x_t[7] = 21'b111111111101011101110;
        x_t[8] = 21'b111111111110100100110;
        x_t[9] = 21'b111111111110111011101;
        x_t[10] = 21'b111111111111011110011;
        x_t[11] = 21'b111111111101000010101;
        x_t[12] = 21'b111111111101011001100;
        x_t[13] = 21'b111111111111001011100;
        x_t[14] = 21'b111111111111010110011;
        x_t[15] = 21'b111111111111101001010;
        x_t[16] = 21'b111111111110110111001;
        x_t[17] = 21'b111111111110001000100;
        x_t[18] = 21'b111111111101000101001;
        x_t[19] = 21'b111111111101010000000;
        x_t[20] = 21'b111111111100100110110;
        x_t[21] = 21'b111111111110110010100;
        x_t[22] = 21'b111111111110010100001;
        x_t[23] = 21'b111111111101100101011;
        x_t[24] = 21'b111111111100111111000;
        x_t[25] = 21'b111111111100111111101;
        x_t[26] = 21'b111111111101000001011;
        x_t[27] = 21'b111111111101001000111;
        x_t[28] = 21'b111111111110011011101;
        x_t[29] = 21'b111111111101011010011;
        x_t[30] = 21'b111111111100110010111;
        x_t[31] = 21'b111111111100011101001;
        x_t[32] = 21'b111111111101101000001;
        x_t[33] = 21'b111111111101000011110;
        x_t[34] = 21'b111111111100010101010;
        x_t[35] = 21'b111111111100101001111;
        x_t[36] = 21'b111111111011111100001;
        x_t[37] = 21'b111111111101101110001;
        x_t[38] = 21'b111111111101001110111;
        x_t[39] = 21'b111111111110110100110;
        x_t[40] = 21'b111111111101101010110;
        x_t[41] = 21'b111111111100100011011;
        x_t[42] = 21'b111111111100110100110;
        x_t[43] = 21'b000000000010000000001;
        x_t[44] = 21'b111111111101010110110;
        x_t[45] = 21'b000000000001000101010;
        x_t[46] = 21'b000000000000010001100;
        x_t[47] = 21'b000000000000000001110;
        x_t[48] = 21'b111111111111000000001;
        x_t[49] = 21'b111111111111010110101;
        x_t[50] = 21'b111111111110000111110;
        x_t[51] = 21'b111111111101111111111;
        x_t[52] = 21'b111111111101100011110;
        x_t[53] = 21'b111111111110011111110;
        x_t[54] = 21'b000000000000101001000;
        x_t[55] = 21'b000000000000111001110;
        x_t[56] = 21'b111111111111101011110;
        x_t[57] = 21'b111111111110101100110;
        x_t[58] = 21'b111111111111110010010;
        x_t[59] = 21'b000000000011010000100;
        x_t[60] = 21'b000000000010010100101;
        x_t[61] = 21'b000000000010111001101;
        x_t[62] = 21'b000000000000011101000;
        x_t[63] = 21'b000000000010000100010;
        
        h_t_prev[0] = 21'b111111111110100110100;
        h_t_prev[1] = 21'b111111111111001100110;
        h_t_prev[2] = 21'b111111111110000011011;
        h_t_prev[3] = 21'b111111111110110000010;
        h_t_prev[4] = 21'b111111111110110011010;
        h_t_prev[5] = 21'b111111111101010111000;
        h_t_prev[6] = 21'b111111111101010100110;
        h_t_prev[7] = 21'b111111111101011101110;
        h_t_prev[8] = 21'b111111111110100100110;
        h_t_prev[9] = 21'b111111111110111011101;
        h_t_prev[10] = 21'b111111111111011110011;
        h_t_prev[11] = 21'b111111111101000010101;
        h_t_prev[12] = 21'b111111111101011001100;
        h_t_prev[13] = 21'b111111111111001011100;
        h_t_prev[14] = 21'b111111111111010110011;
        h_t_prev[15] = 21'b111111111111101001010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 85 timeout!");
                $fdisplay(fd_cycles, "Test Vector  85: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  85: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 85");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 86
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111110100110100;
        x_t[1] = 21'b111111111111010001101;
        x_t[2] = 21'b111111111110010110111;
        x_t[3] = 21'b111111111110101011011;
        x_t[4] = 21'b111111111111001100100;
        x_t[5] = 21'b111111111110000011011;
        x_t[6] = 21'b111111111101100111011;
        x_t[7] = 21'b111111111110010101101;
        x_t[8] = 21'b111111111111010011010;
        x_t[9] = 21'b111111111111011110110;
        x_t[10] = 21'b111111111111101101000;
        x_t[11] = 21'b111111111101100110010;
        x_t[12] = 21'b111111111101111100101;
        x_t[13] = 21'b111111111111001011100;
        x_t[14] = 21'b000000000000010000011;
        x_t[15] = 21'b000000000000011100001;
        x_t[16] = 21'b111111111111010100110;
        x_t[17] = 21'b111111111110100001001;
        x_t[18] = 21'b111111111101011111100;
        x_t[19] = 21'b111111111101101011011;
        x_t[20] = 21'b111111111100111111110;
        x_t[21] = 21'b111111111111011110101;
        x_t[22] = 21'b111111111110110011111;
        x_t[23] = 21'b111111111101101110000;
        x_t[24] = 21'b111111111101101111110;
        x_t[25] = 21'b111111111101101110001;
        x_t[26] = 21'b111111111101110100000;
        x_t[27] = 21'b111111111101101100010;
        x_t[28] = 21'b111111111110011000100;
        x_t[29] = 21'b111111111110101101101;
        x_t[30] = 21'b111111111101110101010;
        x_t[31] = 21'b111111111101101101000;
        x_t[32] = 21'b111111111110101100010;
        x_t[33] = 21'b111111111110001101111;
        x_t[34] = 21'b111111111101101010111;
        x_t[35] = 21'b111111111110000010110;
        x_t[36] = 21'b111111111101010101101;
        x_t[37] = 21'b111111111110011111000;
        x_t[38] = 21'b111111111110100100100;
        x_t[39] = 21'b111111111111111110010;
        x_t[40] = 21'b111111111111101101010;
        x_t[41] = 21'b111111111011111001101;
        x_t[42] = 21'b111111111111110010100;
        x_t[43] = 21'b000000000010000000001;
        x_t[44] = 21'b111111111111001100000;
        x_t[45] = 21'b000000000010010010101;
        x_t[46] = 21'b000000000001000101010;
        x_t[47] = 21'b000000000000101001101;
        x_t[48] = 21'b111111111111101011000;
        x_t[49] = 21'b111111111111100100100;
        x_t[50] = 21'b111111111110010001010;
        x_t[51] = 21'b111111111110000100110;
        x_t[52] = 21'b111111111101110011001;
        x_t[53] = 21'b111111111110110110000;
        x_t[54] = 21'b000000000000010001000;
        x_t[55] = 21'b000000000000110001001;
        x_t[56] = 21'b111111111111100011001;
        x_t[57] = 21'b111111111110011011110;
        x_t[58] = 21'b111111111111011100100;
        x_t[59] = 21'b000000000010010101010;
        x_t[60] = 21'b000000000001111101101;
        x_t[61] = 21'b000000000010001100001;
        x_t[62] = 21'b000000000000100100011;
        x_t[63] = 21'b000000000001100101100;
        
        h_t_prev[0] = 21'b111111111110100110100;
        h_t_prev[1] = 21'b111111111111010001101;
        h_t_prev[2] = 21'b111111111110010110111;
        h_t_prev[3] = 21'b111111111110101011011;
        h_t_prev[4] = 21'b111111111111001100100;
        h_t_prev[5] = 21'b111111111110000011011;
        h_t_prev[6] = 21'b111111111101100111011;
        h_t_prev[7] = 21'b111111111110010101101;
        h_t_prev[8] = 21'b111111111111010011010;
        h_t_prev[9] = 21'b111111111111011110110;
        h_t_prev[10] = 21'b111111111111101101000;
        h_t_prev[11] = 21'b111111111101100110010;
        h_t_prev[12] = 21'b111111111101111100101;
        h_t_prev[13] = 21'b111111111111001011100;
        h_t_prev[14] = 21'b000000000000010000011;
        h_t_prev[15] = 21'b000000000000011100001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 86 timeout!");
                $fdisplay(fd_cycles, "Test Vector  86: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  86: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 86");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 87
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000000001001001;
        x_t[1] = 21'b000000000000010110001;
        x_t[2] = 21'b111111111111010001001;
        x_t[3] = 21'b111111111111010110111;
        x_t[4] = 21'b000000000000001110010;
        x_t[5] = 21'b111111111111101100110;
        x_t[6] = 21'b111111111111110110100;
        x_t[7] = 21'b111111111111010111111;
        x_t[8] = 21'b000000000000000001101;
        x_t[9] = 21'b000000000000010000111;
        x_t[10] = 21'b000000000000100010111;
        x_t[11] = 21'b111111111110011110011;
        x_t[12] = 21'b111111111111110111100;
        x_t[13] = 21'b000000000001000110010;
        x_t[14] = 21'b000000000001001010011;
        x_t[15] = 21'b000000000000110101100;
        x_t[16] = 21'b111111111111111100100;
        x_t[17] = 21'b111111111111001000101;
        x_t[18] = 21'b111111111110101110100;
        x_t[19] = 21'b111111111111001000110;
        x_t[20] = 21'b111111111110101010001;
        x_t[21] = 21'b000000000000110111001;
        x_t[22] = 21'b000000000000011001100;
        x_t[23] = 21'b111111111111010000101;
        x_t[24] = 21'b111111111111001110001;
        x_t[25] = 21'b111111111111001011011;
        x_t[26] = 21'b111111111110110011011;
        x_t[27] = 21'b111111111111010110011;
        x_t[28] = 21'b111111111111111010001;
        x_t[29] = 21'b000000000000100110010;
        x_t[30] = 21'b111111111111011010110;
        x_t[31] = 21'b111111111110011001010;
        x_t[32] = 21'b111111111111010000101;
        x_t[33] = 21'b111111111110101001101;
        x_t[34] = 21'b111111111110011010100;
        x_t[35] = 21'b111111111110111101111;
        x_t[36] = 21'b111111111111000011000;
        x_t[37] = 21'b111111111111111000110;
        x_t[38] = 21'b000000000000001001011;
        x_t[39] = 21'b000000000010101110101;
        x_t[40] = 21'b000000000010000000000;
        x_t[41] = 21'b000000000000100100110;
        x_t[42] = 21'b000000000000111001101;
        x_t[43] = 21'b000000000010001011001;
        x_t[44] = 21'b111111111111110011001;
        x_t[45] = 21'b000000000011001000110;
        x_t[46] = 21'b000000000001100100011;
        x_t[47] = 21'b000000000001010110011;
        x_t[48] = 21'b000000000000001100011;
        x_t[49] = 21'b111111111111111011101;
        x_t[50] = 21'b111111111110110111010;
        x_t[51] = 21'b111111111110001110011;
        x_t[52] = 21'b111111111110001100101;
        x_t[53] = 21'b111111111111010001111;
        x_t[54] = 21'b111111111111111001000;
        x_t[55] = 21'b000000000001001011000;
        x_t[56] = 21'b000000000000010010011;
        x_t[57] = 21'b111111111110100100010;
        x_t[58] = 21'b111111111110110000111;
        x_t[59] = 21'b000000000000101110101;
        x_t[60] = 21'b000000000001001011111;
        x_t[61] = 21'b000000000000101000110;
        x_t[62] = 21'b111111111111000100010;
        x_t[63] = 21'b111111111111111011111;
        
        h_t_prev[0] = 21'b000000000000001001001;
        h_t_prev[1] = 21'b000000000000010110001;
        h_t_prev[2] = 21'b111111111111010001001;
        h_t_prev[3] = 21'b111111111111010110111;
        h_t_prev[4] = 21'b000000000000001110010;
        h_t_prev[5] = 21'b111111111111101100110;
        h_t_prev[6] = 21'b111111111111110110100;
        h_t_prev[7] = 21'b111111111111010111111;
        h_t_prev[8] = 21'b000000000000000001101;
        h_t_prev[9] = 21'b000000000000010000111;
        h_t_prev[10] = 21'b000000000000100010111;
        h_t_prev[11] = 21'b111111111110011110011;
        h_t_prev[12] = 21'b111111111111110111100;
        h_t_prev[13] = 21'b000000000001000110010;
        h_t_prev[14] = 21'b000000000001001010011;
        h_t_prev[15] = 21'b000000000000110101100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 87 timeout!");
                $fdisplay(fd_cycles, "Test Vector  87: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  87: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 87");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 88
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000000111111011;
        x_t[1] = 21'b000000000001000010001;
        x_t[2] = 21'b111111111111110111111;
        x_t[3] = 21'b111111111111111101100;
        x_t[4] = 21'b000000000000100010011;
        x_t[5] = 21'b000000000000000011000;
        x_t[6] = 21'b000000000000000011000;
        x_t[7] = 21'b000000000000011111001;
        x_t[8] = 21'b000000000000111010011;
        x_t[9] = 21'b000000000001001101000;
        x_t[10] = 21'b000000000010000100101;
        x_t[11] = 21'b111111111111010110011;
        x_t[12] = 21'b000000000000110111111;
        x_t[13] = 21'b000000000001101111001;
        x_t[14] = 21'b000000000010100100000;
        x_t[15] = 21'b000000000001111100110;
        x_t[16] = 21'b000000000001000001111;
        x_t[17] = 21'b000000000000010010101;
        x_t[18] = 21'b111111111111110011001;
        x_t[19] = 21'b000000000000010000001;
        x_t[20] = 21'b111111111111101111000;
        x_t[21] = 21'b111111111111110100110;
        x_t[22] = 21'b000000000000000011010;
        x_t[23] = 21'b111111111111000010001;
        x_t[24] = 21'b111111111110101111101;
        x_t[25] = 21'b111111111110101001010;
        x_t[26] = 21'b111111111110001001001;
        x_t[27] = 21'b111111111110111110110;
        x_t[28] = 21'b111111111111111101010;
        x_t[29] = 21'b000000000000000000110;
        x_t[30] = 21'b111111111110100100001;
        x_t[31] = 21'b111111111110000111100;
        x_t[32] = 21'b111111111111000011000;
        x_t[33] = 21'b111111111110001101111;
        x_t[34] = 21'b111111111101100110001;
        x_t[35] = 21'b111111111110000111101;
        x_t[36] = 21'b111111111101111101011;
        x_t[37] = 21'b111111111110001110110;
        x_t[38] = 21'b111111111111111111011;
        x_t[39] = 21'b000000000001010110011;
        x_t[40] = 21'b000000000011000001001;
        x_t[41] = 21'b111111111101101111111;
        x_t[42] = 21'b111111111110000111110;
        x_t[43] = 21'b000000000011101101111;
        x_t[44] = 21'b000000000000100101011;
        x_t[45] = 21'b000000000011011000010;
        x_t[46] = 21'b000000000011100101111;
        x_t[47] = 21'b000000000011001101110;
        x_t[48] = 21'b000000000001100110111;
        x_t[49] = 21'b000000000001101010111;
        x_t[50] = 21'b000000000000001100110;
        x_t[51] = 21'b111111111110101011011;
        x_t[52] = 21'b111111111110100001001;
        x_t[53] = 21'b111111111111010001111;
        x_t[54] = 21'b111111111111011011001;
        x_t[55] = 21'b000000000010010000000;
        x_t[56] = 21'b000000000010000010001;
        x_t[57] = 21'b111111111111001110111;
        x_t[58] = 21'b111111111101101011000;
        x_t[59] = 21'b111111111111000000001;
        x_t[60] = 21'b000000000001000100001;
        x_t[61] = 21'b111111111111001001101;
        x_t[62] = 21'b111111111100100101001;
        x_t[63] = 21'b111111111110101100101;
        
        h_t_prev[0] = 21'b000000000000111111011;
        h_t_prev[1] = 21'b000000000001000010001;
        h_t_prev[2] = 21'b111111111111110111111;
        h_t_prev[3] = 21'b111111111111111101100;
        h_t_prev[4] = 21'b000000000000100010011;
        h_t_prev[5] = 21'b000000000000000011000;
        h_t_prev[6] = 21'b000000000000000011000;
        h_t_prev[7] = 21'b000000000000011111001;
        h_t_prev[8] = 21'b000000000000111010011;
        h_t_prev[9] = 21'b000000000001001101000;
        h_t_prev[10] = 21'b000000000010000100101;
        h_t_prev[11] = 21'b111111111111010110011;
        h_t_prev[12] = 21'b000000000000110111111;
        h_t_prev[13] = 21'b000000000001101111001;
        h_t_prev[14] = 21'b000000000010100100000;
        h_t_prev[15] = 21'b000000000001111100110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 88 timeout!");
                $fdisplay(fd_cycles, "Test Vector  88: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  88: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 88");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 89
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000001011000001;
        x_t[1] = 21'b000000000001000111001;
        x_t[2] = 21'b000000000000001011011;
        x_t[3] = 21'b000000000000101101111;
        x_t[4] = 21'b000000000001001010111;
        x_t[5] = 21'b111111111111111101011;
        x_t[6] = 21'b111111111110100101101;
        x_t[7] = 21'b000000000001000010110;
        x_t[8] = 21'b000000000000110101010;
        x_t[9] = 21'b000000000001011100000;
        x_t[10] = 21'b000000000010101011111;
        x_t[11] = 21'b111111111111111111001;
        x_t[12] = 21'b000000000001010101010;
        x_t[13] = 21'b000000000001110101111;
        x_t[14] = 21'b000000000010110011111;
        x_t[15] = 21'b000000000001110111101;
        x_t[16] = 21'b000000000001011111101;
        x_t[17] = 21'b000000000001000100000;
        x_t[18] = 21'b000000000000001101011;
        x_t[19] = 21'b000000000000011011001;
        x_t[20] = 21'b111111111111110101010;
        x_t[21] = 21'b111111111111011011111;
        x_t[22] = 21'b111111111111101001111;
        x_t[23] = 21'b111111111110100101001;
        x_t[24] = 21'b111111111110101001101;
        x_t[25] = 21'b111111111110100011000;
        x_t[26] = 21'b111111111110011010000;
        x_t[27] = 21'b111111111110011111011;
        x_t[28] = 21'b111111111111010001001;
        x_t[29] = 21'b000000000000000000110;
        x_t[30] = 21'b111111111110010100100;
        x_t[31] = 21'b111111111110010000011;
        x_t[32] = 21'b111111111111110000011;
        x_t[33] = 21'b111111111111000000110;
        x_t[34] = 21'b111111111110000111100;
        x_t[35] = 21'b111111111110111001000;
        x_t[36] = 21'b111111111101110011100;
        x_t[37] = 21'b111111111101100001111;
        x_t[38] = 21'b000000000000100010101;
        x_t[39] = 21'b000000000000000101101;
        x_t[40] = 21'b000000000001001111000;
        x_t[41] = 21'b111111111011010000000;
        x_t[42] = 21'b111111111110011001101;
        x_t[43] = 21'b000000000010000000001;
        x_t[44] = 21'b111111111110110101101;
        x_t[45] = 21'b000000000001100100001;
        x_t[46] = 21'b000000000001001111101;
        x_t[47] = 21'b000000000001101111010;
        x_t[48] = 21'b000000000000110010100;
        x_t[49] = 21'b000000000001001010011;
        x_t[50] = 21'b111111111111110000010;
        x_t[51] = 21'b111111111101010100100;
        x_t[52] = 21'b111111111101001111010;
        x_t[53] = 21'b111111111100111011100;
        x_t[54] = 21'b111111111100100111010;
        x_t[55] = 21'b000000000000010111001;
        x_t[56] = 21'b000000000000101100001;
        x_t[57] = 21'b111111111101101100111;
        x_t[58] = 21'b111111111010100010011;
        x_t[59] = 21'b111111111010010100001;
        x_t[60] = 21'b111111111111111111001;
        x_t[61] = 21'b111111111100110100101;
        x_t[62] = 21'b111111111000110001001;
        x_t[63] = 21'b111111111100010111000;
        
        h_t_prev[0] = 21'b000000000001011000001;
        h_t_prev[1] = 21'b000000000001000111001;
        h_t_prev[2] = 21'b000000000000001011011;
        h_t_prev[3] = 21'b000000000000101101111;
        h_t_prev[4] = 21'b000000000001001010111;
        h_t_prev[5] = 21'b111111111111111101011;
        h_t_prev[6] = 21'b111111111110100101101;
        h_t_prev[7] = 21'b000000000001000010110;
        h_t_prev[8] = 21'b000000000000110101010;
        h_t_prev[9] = 21'b000000000001011100000;
        h_t_prev[10] = 21'b000000000010101011111;
        h_t_prev[11] = 21'b111111111111111111001;
        h_t_prev[12] = 21'b000000000001010101010;
        h_t_prev[13] = 21'b000000000001110101111;
        h_t_prev[14] = 21'b000000000010110011111;
        h_t_prev[15] = 21'b000000000001110111101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 89 timeout!");
                $fdisplay(fd_cycles, "Test Vector  89: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  89: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 89");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 90
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000001110000110;
        x_t[1] = 21'b000000000001101110010;
        x_t[2] = 21'b000000000001001010100;
        x_t[3] = 21'b000000000001111011010;
        x_t[4] = 21'b000000000010100101110;
        x_t[5] = 21'b000000000001011011110;
        x_t[6] = 21'b000000000000000011000;
        x_t[7] = 21'b000000000000000000100;
        x_t[8] = 21'b000000000000100101110;
        x_t[9] = 21'b000000000001111010001;
        x_t[10] = 21'b000000000011011100110;
        x_t[11] = 21'b000000000001100101001;
        x_t[12] = 21'b000000000001110010100;
        x_t[13] = 21'b000000000001101111001;
        x_t[14] = 21'b000000000000100000001;
        x_t[15] = 21'b000000000000111010101;
        x_t[16] = 21'b000000000001010000110;
        x_t[17] = 21'b000000000001001101111;
        x_t[18] = 21'b000000000000011000000;
        x_t[19] = 21'b111111111111111010010;
        x_t[20] = 21'b111111111110111101000;
        x_t[21] = 21'b000000000000011011100;
        x_t[22] = 21'b000000000000101001010;
        x_t[23] = 21'b111111111111110000100;
        x_t[24] = 21'b111111111111000101000;
        x_t[25] = 21'b111111111111000010001;
        x_t[26] = 21'b000000000000000011101;
        x_t[27] = 21'b000000000000001101011;
        x_t[28] = 21'b000000000000101100100;
        x_t[29] = 21'b111111111111011011011;
        x_t[30] = 21'b111111111111001111000;
        x_t[31] = 21'b111111111111110110100;
        x_t[32] = 21'b000000000000111101101;
        x_t[33] = 21'b000000000000111101101;
        x_t[34] = 21'b000000000000000011011;
        x_t[35] = 21'b000000000000011011110;
        x_t[36] = 21'b000000000000010010100;
        x_t[37] = 21'b000000000000011101011;
        x_t[38] = 21'b111111111111110000010;
        x_t[39] = 21'b000000000010111101011;
        x_t[40] = 21'b111111111111110010101;
        x_t[41] = 21'b111111111100010101100;
        x_t[42] = 21'b111111111100110100110;
        x_t[43] = 21'b000000000000000111100;
        x_t[44] = 21'b111111111100111010110;
        x_t[45] = 21'b000000000000100110010;
        x_t[46] = 21'b111111111110010101001;
        x_t[47] = 21'b111111111111010000001;
        x_t[48] = 21'b111111111110110110101;
        x_t[49] = 21'b111111111111110111000;
        x_t[50] = 21'b111111111111000101100;
        x_t[51] = 21'b111111111100000111001;
        x_t[52] = 21'b111111111011111000011;
        x_t[53] = 21'b111111111010110000011;
        x_t[54] = 21'b111111111001111111100;
        x_t[55] = 21'b111111111101110111100;
        x_t[56] = 21'b111111111110010001100;
        x_t[57] = 21'b111111111100000110100;
        x_t[58] = 21'b111111111000010110110;
        x_t[59] = 21'b111111110110100011011;
        x_t[60] = 21'b111111111101011010010;
        x_t[61] = 21'b111111111001011101011;
        x_t[62] = 21'b111111110100011000000;
        x_t[63] = 21'b111111111000101101110;
        
        h_t_prev[0] = 21'b000000000001110000110;
        h_t_prev[1] = 21'b000000000001101110010;
        h_t_prev[2] = 21'b000000000001001010100;
        h_t_prev[3] = 21'b000000000001111011010;
        h_t_prev[4] = 21'b000000000010100101110;
        h_t_prev[5] = 21'b000000000001011011110;
        h_t_prev[6] = 21'b000000000000000011000;
        h_t_prev[7] = 21'b000000000000000000100;
        h_t_prev[8] = 21'b000000000000100101110;
        h_t_prev[9] = 21'b000000000001111010001;
        h_t_prev[10] = 21'b000000000011011100110;
        h_t_prev[11] = 21'b000000000001100101001;
        h_t_prev[12] = 21'b000000000001110010100;
        h_t_prev[13] = 21'b000000000001101111001;
        h_t_prev[14] = 21'b000000000000100000001;
        h_t_prev[15] = 21'b000000000000111010101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 90 timeout!");
                $fdisplay(fd_cycles, "Test Vector  90: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  90: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 90");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 91
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000001000100011;
        x_t[1] = 21'b000000000010010000100;
        x_t[2] = 21'b000000000010101011101;
        x_t[3] = 21'b000000000011100101101;
        x_t[4] = 21'b000000000011100111011;
        x_t[5] = 21'b000000000010001000001;
        x_t[6] = 21'b000000000001011010001;
        x_t[7] = 21'b000000000000000000100;
        x_t[8] = 21'b000000000000111111100;
        x_t[9] = 21'b000000000011000000010;
        x_t[10] = 21'b000000000100101111111;
        x_t[11] = 21'b000000000001111001100;
        x_t[12] = 21'b000000000001100000111;
        x_t[13] = 21'b000000000001010011111;
        x_t[14] = 21'b111111111111010110011;
        x_t[15] = 21'b000000000000111111101;
        x_t[16] = 21'b000000000001011111101;
        x_t[17] = 21'b000000000001100001101;
        x_t[18] = 21'b000000000000100010100;
        x_t[19] = 21'b111111111111100100010;
        x_t[20] = 21'b111111111110001010111;
        x_t[21] = 21'b000000000000110111001;
        x_t[22] = 21'b000000000001000010110;
        x_t[23] = 21'b000000000000010011011;
        x_t[24] = 21'b111111111111010111010;
        x_t[25] = 21'b111111111111010100110;
        x_t[26] = 21'b000000000000110110011;
        x_t[27] = 21'b000000000000110000110;
        x_t[28] = 21'b000000000001010010010;
        x_t[29] = 21'b111111111111011011011;
        x_t[30] = 21'b111111111111111001111;
        x_t[31] = 21'b000000000000101011101;
        x_t[32] = 21'b000000000010000001110;
        x_t[33] = 21'b000000000010000111101;
        x_t[34] = 21'b000000000001001111100;
        x_t[35] = 21'b000000000001001101000;
        x_t[36] = 21'b000000000000101011011;
        x_t[37] = 21'b000000000000001001000;
        x_t[38] = 21'b111111111111001100111;
        x_t[39] = 21'b000000000011000100101;
        x_t[40] = 21'b111111111110110001100;
        x_t[41] = 21'b111111111111101101001;
        x_t[42] = 21'b111111111110110111010;
        x_t[43] = 21'b000000000011101101111;
        x_t[44] = 21'b111111111110100100111;
        x_t[45] = 21'b000000000000010110110;
        x_t[46] = 21'b111111111110110100010;
        x_t[47] = 21'b111111111111100100000;
        x_t[48] = 21'b111111111111001110011;
        x_t[49] = 21'b000000000000110111111;
        x_t[50] = 21'b000000000000011111110;
        x_t[51] = 21'b111111111101110001011;
        x_t[52] = 21'b111111111101010100011;
        x_t[53] = 21'b111111111100010100101;
        x_t[54] = 21'b111111111011010011011;
        x_t[55] = 21'b111111111110001101001;
        x_t[56] = 21'b111111111110101111100;
        x_t[57] = 21'b111111111101111001101;
        x_t[58] = 21'b111111111010011001101;
        x_t[59] = 21'b111111111000111001011;
        x_t[60] = 21'b111111111011101111000;
        x_t[61] = 21'b111111111000000010011;
        x_t[62] = 21'b111111110010110111110;
        x_t[63] = 21'b111111110111110000010;
        
        h_t_prev[0] = 21'b000000000001000100011;
        h_t_prev[1] = 21'b000000000010010000100;
        h_t_prev[2] = 21'b000000000010101011101;
        h_t_prev[3] = 21'b000000000011100101101;
        h_t_prev[4] = 21'b000000000011100111011;
        h_t_prev[5] = 21'b000000000010001000001;
        h_t_prev[6] = 21'b000000000001011010001;
        h_t_prev[7] = 21'b000000000000000000100;
        h_t_prev[8] = 21'b000000000000111111100;
        h_t_prev[9] = 21'b000000000011000000010;
        h_t_prev[10] = 21'b000000000100101111111;
        h_t_prev[11] = 21'b000000000001111001100;
        h_t_prev[12] = 21'b000000000001100000111;
        h_t_prev[13] = 21'b000000000001010011111;
        h_t_prev[14] = 21'b111111111111010110011;
        h_t_prev[15] = 21'b000000000000111111101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 91 timeout!");
                $fdisplay(fd_cycles, "Test Vector  91: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  91: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 91");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 92
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000001110000110;
        x_t[1] = 21'b000000000011010101000;
        x_t[2] = 21'b000000000011110100011;
        x_t[3] = 21'b000000000100100100011;
        x_t[4] = 21'b000000000100001010110;
        x_t[5] = 21'b000000000010011110010;
        x_t[6] = 21'b000000000001011010001;
        x_t[7] = 21'b000000000000001010110;
        x_t[8] = 21'b000000000010101011111;
        x_t[9] = 21'b000000000100101110100;
        x_t[10] = 21'b000000000110001100111;
        x_t[11] = 21'b000000000010011000000;
        x_t[12] = 21'b000000000010000100000;
        x_t[13] = 21'b000000000010101100011;
        x_t[14] = 21'b000000000000110101010;
        x_t[15] = 21'b000000000010101111100;
        x_t[16] = 21'b000000000011100101100;
        x_t[17] = 21'b000000000011011101000;
        x_t[18] = 21'b000000000010000001011;
        x_t[19] = 21'b000000000000110110101;
        x_t[20] = 21'b111111111111010110000;
        x_t[21] = 21'b000000000001011011000;
        x_t[22] = 21'b000000000001000101111;
        x_t[23] = 21'b111111111111110011100;
        x_t[24] = 21'b000000000000101001100;
        x_t[25] = 21'b000000000000100010100;
        x_t[26] = 21'b000000000000110010001;
        x_t[27] = 21'b000000000000011001010;
        x_t[28] = 21'b000000000000101100100;
        x_t[29] = 21'b000000000010010010011;
        x_t[30] = 21'b111111111111100110011;
        x_t[31] = 21'b000000000000011110011;
        x_t[32] = 21'b000000000010001010111;
        x_t[33] = 21'b000000000001111001110;
        x_t[34] = 21'b000000000001010100011;
        x_t[35] = 21'b000000000001010110111;
        x_t[36] = 21'b000000000000001101100;
        x_t[37] = 21'b111111111110100111010;
        x_t[38] = 21'b000000000001110011010;
        x_t[39] = 21'b000000000011000100101;
        x_t[40] = 21'b000000000010100110000;
        x_t[41] = 21'b111111111111011111001;
        x_t[42] = 21'b000000000010000110110;
        x_t[43] = 21'b000000000000111110011;
        x_t[44] = 21'b000000000000110000100;
        x_t[45] = 21'b000000000000010110110;
        x_t[46] = 21'b000000000000100110010;
        x_t[47] = 21'b000000000001001100011;
        x_t[48] = 21'b000000000000100100001;
        x_t[49] = 21'b000000000010011101110;
        x_t[50] = 21'b000000000010100100110;
        x_t[51] = 21'b111111111111111101100;
        x_t[52] = 21'b111111111111011001011;
        x_t[53] = 21'b111111111101111110011;
        x_t[54] = 21'b111111111100011011010;
        x_t[55] = 21'b111111111111001001100;
        x_t[56] = 21'b000000000000000001001;
        x_t[57] = 21'b000000000000001010101;
        x_t[58] = 21'b111111111101001000001;
        x_t[59] = 21'b111111111011100011000;
        x_t[60] = 21'b111111111100001001110;
        x_t[61] = 21'b111111111001100101101;
        x_t[62] = 21'b111111110100110101100;
        x_t[63] = 21'b111111110111110100101;
        
        h_t_prev[0] = 21'b000000000001110000110;
        h_t_prev[1] = 21'b000000000011010101000;
        h_t_prev[2] = 21'b000000000011110100011;
        h_t_prev[3] = 21'b000000000100100100011;
        h_t_prev[4] = 21'b000000000100001010110;
        h_t_prev[5] = 21'b000000000010011110010;
        h_t_prev[6] = 21'b000000000001011010001;
        h_t_prev[7] = 21'b000000000000001010110;
        h_t_prev[8] = 21'b000000000010101011111;
        h_t_prev[9] = 21'b000000000100101110100;
        h_t_prev[10] = 21'b000000000110001100111;
        h_t_prev[11] = 21'b000000000010011000000;
        h_t_prev[12] = 21'b000000000010000100000;
        h_t_prev[13] = 21'b000000000010101100011;
        h_t_prev[14] = 21'b000000000000110101010;
        h_t_prev[15] = 21'b000000000010101111100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 92 timeout!");
                $fdisplay(fd_cycles, "Test Vector  92: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  92: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 92");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 93
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000011010011011;
        x_t[1] = 21'b000000000100101101001;
        x_t[2] = 21'b000000000100111000011;
        x_t[3] = 21'b000000000101011001101;
        x_t[4] = 21'b000000000100111000010;
        x_t[5] = 21'b000000000011011011010;
        x_t[6] = 21'b000000000010010010001;
        x_t[7] = 21'b000000000010101101101;
        x_t[8] = 21'b000000000100110111001;
        x_t[9] = 21'b000000000110101011110;
        x_t[10] = 21'b000000001000001100001;
        x_t[11] = 21'b000000000100110000111;
        x_t[12] = 21'b000000000011100111100;
        x_t[13] = 21'b000000000011100010111;
        x_t[14] = 21'b000000000011111101101;
        x_t[15] = 21'b000000000101101011110;
        x_t[16] = 21'b000000000110010111111;
        x_t[17] = 21'b000000000110001001110;
        x_t[18] = 21'b000000000100111001111;
        x_t[19] = 21'b000000000011110001011;
        x_t[20] = 21'b000000000001011111101;
        x_t[21] = 21'b000000000010010101000;
        x_t[22] = 21'b000000000010000010001;
        x_t[23] = 21'b000000000000110011010;
        x_t[24] = 21'b000000000001100000010;
        x_t[25] = 21'b000000000001011010011;
        x_t[26] = 21'b000000000001110101110;
        x_t[27] = 21'b000000000001110111100;
        x_t[28] = 21'b000000000001111000000;
        x_t[29] = 21'b000000000011000100010;
        x_t[30] = 21'b000000000000101000110;
        x_t[31] = 21'b000000000010001000111;
        x_t[32] = 21'b000000000011011100101;
        x_t[33] = 21'b000000000011010001101;
        x_t[34] = 21'b000000000010100101010;
        x_t[35] = 21'b000000000010110100101;
        x_t[36] = 21'b000000000010000100110;
        x_t[37] = 21'b000000000000001001000;
        x_t[38] = 21'b000000000011100111010;
        x_t[39] = 21'b000000000100000110110;
        x_t[40] = 21'b000000000101101111001;
        x_t[41] = 21'b000000000000010110110;
        x_t[42] = 21'b000000000010001100101;
        x_t[43] = 21'b111111111111000101101;
        x_t[44] = 21'b000000000011111001101;
        x_t[45] = 21'b000000000011001000110;
        x_t[46] = 21'b000000000011100000110;
        x_t[47] = 21'b000000000100011000010;
        x_t[48] = 21'b000000000011100111100;
        x_t[49] = 21'b000000000101010010100;
        x_t[50] = 21'b000000000101100010111;
        x_t[51] = 21'b000000000011111101100;
        x_t[52] = 21'b000000000011011001010;
        x_t[53] = 21'b000000000001110011011;
        x_t[54] = 21'b000000000000010111000;
        x_t[55] = 21'b000000000001110001110;
        x_t[56] = 21'b000000000010100100100;
        x_t[57] = 21'b000000000011001010011;
        x_t[58] = 21'b000000000001010010010;
        x_t[59] = 21'b111111111111100111101;
        x_t[60] = 21'b111111111110110110010;
        x_t[61] = 21'b111111111101010101110;
        x_t[62] = 21'b111111111001110000000;
        x_t[63] = 21'b111111111001111000101;
        
        h_t_prev[0] = 21'b000000000011010011011;
        h_t_prev[1] = 21'b000000000100101101001;
        h_t_prev[2] = 21'b000000000100111000011;
        h_t_prev[3] = 21'b000000000101011001101;
        h_t_prev[4] = 21'b000000000100111000010;
        h_t_prev[5] = 21'b000000000011011011010;
        h_t_prev[6] = 21'b000000000010010010001;
        h_t_prev[7] = 21'b000000000010101101101;
        h_t_prev[8] = 21'b000000000100110111001;
        h_t_prev[9] = 21'b000000000110101011110;
        h_t_prev[10] = 21'b000000001000001100001;
        h_t_prev[11] = 21'b000000000100110000111;
        h_t_prev[12] = 21'b000000000011100111100;
        h_t_prev[13] = 21'b000000000011100010111;
        h_t_prev[14] = 21'b000000000011111101101;
        h_t_prev[15] = 21'b000000000101101011110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 93 timeout!");
                $fdisplay(fd_cycles, "Test Vector  93: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  93: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 93");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 94
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000100100010010;
        x_t[1] = 21'b000000000101111011011;
        x_t[2] = 21'b000000000101110111100;
        x_t[3] = 21'b000000000110000101001;
        x_t[4] = 21'b000000000101101111111;
        x_t[5] = 21'b000000000100001101010;
        x_t[6] = 21'b000000000011000011111;
        x_t[7] = 21'b000000000100001001010;
        x_t[8] = 21'b000000000101111111010;
        x_t[9] = 21'b000000000111000100111;
        x_t[10] = 21'b000000001000000111001;
        x_t[11] = 21'b000000000101101110000;
        x_t[12] = 21'b000000000100111111011;
        x_t[13] = 21'b000000000100110100110;
        x_t[14] = 21'b000000000100111100111;
        x_t[15] = 21'b000000000110001010010;
        x_t[16] = 21'b000000000110101011110;
        x_t[17] = 21'b000000000101111111111;
        x_t[18] = 21'b000000000101100100000;
        x_t[19] = 21'b000000000101010100010;
        x_t[20] = 21'b000000000011010000010;
        x_t[21] = 21'b000000000001100110000;
        x_t[22] = 21'b000000000001001100010;
        x_t[23] = 21'b111111111111100111111;
        x_t[24] = 21'b000000000000010001001;
        x_t[25] = 21'b000000000000001111110;
        x_t[26] = 21'b000000000000111010100;
        x_t[27] = 21'b000000000000011101001;
        x_t[28] = 21'b111111111111110000101;
        x_t[29] = 21'b000000000001100000011;
        x_t[30] = 21'b000000000000000001110;
        x_t[31] = 21'b000000000000110100100;
        x_t[32] = 21'b000000000010010011111;
        x_t[33] = 21'b000000000001111001110;
        x_t[34] = 21'b000000000000111100100;
        x_t[35] = 21'b000000000001001000001;
        x_t[36] = 21'b111111111111101010110;
        x_t[37] = 21'b111111111110011111000;
        x_t[38] = 21'b000000000010010001100;
        x_t[39] = 21'b000000000010100111010;
        x_t[40] = 21'b000000000011100111010;
        x_t[41] = 21'b111111111110111100011;
        x_t[42] = 21'b000000000000001010010;
        x_t[43] = 21'b111111111011110101010;
        x_t[44] = 21'b000000000001110011101;
        x_t[45] = 21'b000000000010010010101;
        x_t[46] = 21'b000000000010110010001;
        x_t[47] = 21'b000000000011011100101;
        x_t[48] = 21'b000000000010100000000;
        x_t[49] = 21'b000000000100000011110;
        x_t[50] = 21'b000000000011110101100;
        x_t[51] = 21'b000000000011101111000;
        x_t[52] = 21'b000000000011001111000;
        x_t[53] = 21'b000000000010000100000;
        x_t[54] = 21'b000000000000100011000;
        x_t[55] = 21'b000000000001100000100;
        x_t[56] = 21'b000000000001110101010;
        x_t[57] = 21'b000000000010111101101;
        x_t[58] = 21'b000000000010001111010;
        x_t[59] = 21'b000000000001001110010;
        x_t[60] = 21'b000000000001010011100;
        x_t[61] = 21'b000000000000100100101;
        x_t[62] = 21'b111111111110010000100;
        x_t[63] = 21'b111111111100010111000;
        
        h_t_prev[0] = 21'b000000000100100010010;
        h_t_prev[1] = 21'b000000000101111011011;
        h_t_prev[2] = 21'b000000000101110111100;
        h_t_prev[3] = 21'b000000000110000101001;
        h_t_prev[4] = 21'b000000000101101111111;
        h_t_prev[5] = 21'b000000000100001101010;
        h_t_prev[6] = 21'b000000000011000011111;
        h_t_prev[7] = 21'b000000000100001001010;
        h_t_prev[8] = 21'b000000000101111111010;
        h_t_prev[9] = 21'b000000000111000100111;
        h_t_prev[10] = 21'b000000001000000111001;
        h_t_prev[11] = 21'b000000000101101110000;
        h_t_prev[12] = 21'b000000000100111111011;
        h_t_prev[13] = 21'b000000000100110100110;
        h_t_prev[14] = 21'b000000000100111100111;
        h_t_prev[15] = 21'b000000000110001010010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 94 timeout!");
                $fdisplay(fd_cycles, "Test Vector  94: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  94: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 94");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 95
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000010001110011;
        x_t[1] = 21'b000000000011010000001;
        x_t[2] = 21'b000000000010110000100;
        x_t[3] = 21'b000000000010100110110;
        x_t[4] = 21'b000000000010000111100;
        x_t[5] = 21'b000000000000011001001;
        x_t[6] = 21'b111111111110011111011;
        x_t[7] = 21'b000000000001111010110;
        x_t[8] = 21'b000000000011101001110;
        x_t[9] = 21'b000000000011111100011;
        x_t[10] = 21'b000000000100111001110;
        x_t[11] = 21'b000000000010101100011;
        x_t[12] = 21'b000000000010100001010;
        x_t[13] = 21'b000000000001101000010;
        x_t[14] = 21'b000000000010111110011;
        x_t[15] = 21'b000000000100000110000;
        x_t[16] = 21'b000000000100011100000;
        x_t[17] = 21'b000000000011110000110;
        x_t[18] = 21'b000000000011111010101;
        x_t[19] = 21'b000000000011110110111;
        x_t[20] = 21'b000000000010000101001;
        x_t[21] = 21'b111111111111011001001;
        x_t[22] = 21'b111111111111001101010;
        x_t[23] = 21'b111111111110001011000;
        x_t[24] = 21'b111111111110001110010;
        x_t[25] = 21'b111111111110010011100;
        x_t[26] = 21'b111111111110010001101;
        x_t[27] = 21'b111111111110001011110;
        x_t[28] = 21'b111111111111100000111;
        x_t[29] = 21'b111111111111100011101;
        x_t[30] = 21'b111111111110001100101;
        x_t[31] = 21'b111111111101111010010;
        x_t[32] = 21'b111111111111110100111;
        x_t[33] = 21'b111111111110110111100;
        x_t[34] = 21'b111111111101111001010;
        x_t[35] = 21'b111111111110011011011;
        x_t[36] = 21'b111111111100110111111;
        x_t[37] = 21'b111111111101001101100;
        x_t[38] = 21'b111111111111111111011;
        x_t[39] = 21'b111111111111111110010;
        x_t[40] = 21'b000000000000111001011;
        x_t[41] = 21'b111111111010111011001;
        x_t[42] = 21'b000000000000000100010;
        x_t[43] = 21'b000000000010101100000;
        x_t[44] = 21'b000000000000111011110;
        x_t[45] = 21'b000000000011010000100;
        x_t[46] = 21'b000000000011011011100;
        x_t[47] = 21'b000000000011100001101;
        x_t[48] = 21'b000000000011000001011;
        x_t[49] = 21'b000000000100100100001;
        x_t[50] = 21'b000000000100011011100;
        x_t[51] = 21'b000000000100111100010;
        x_t[52] = 21'b000000000100100101111;
        x_t[53] = 21'b000000000011111110100;
        x_t[54] = 21'b000000000011000100110;
        x_t[55] = 21'b000000000011001000001;
        x_t[56] = 21'b000000000011100100111;
        x_t[57] = 21'b000000000100111101100;
        x_t[58] = 21'b000000000100110101000;
        x_t[59] = 21'b000000000100101011010;
        x_t[60] = 21'b000000000011011001101;
        x_t[61] = 21'b000000000011110011100;
        x_t[62] = 21'b000000000001101010101;
        x_t[63] = 21'b111111111111110011001;
        
        h_t_prev[0] = 21'b000000000010001110011;
        h_t_prev[1] = 21'b000000000011010000001;
        h_t_prev[2] = 21'b000000000010110000100;
        h_t_prev[3] = 21'b000000000010100110110;
        h_t_prev[4] = 21'b000000000010000111100;
        h_t_prev[5] = 21'b000000000000011001001;
        h_t_prev[6] = 21'b111111111110011111011;
        h_t_prev[7] = 21'b000000000001111010110;
        h_t_prev[8] = 21'b000000000011101001110;
        h_t_prev[9] = 21'b000000000011111100011;
        h_t_prev[10] = 21'b000000000100111001110;
        h_t_prev[11] = 21'b000000000010101100011;
        h_t_prev[12] = 21'b000000000010100001010;
        h_t_prev[13] = 21'b000000000001101000010;
        h_t_prev[14] = 21'b000000000010111110011;
        h_t_prev[15] = 21'b000000000100000110000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 95 timeout!");
                $fdisplay(fd_cycles, "Test Vector  95: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  95: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 95");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 96
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000001000100011;
        x_t[1] = 21'b000000000001111100111;
        x_t[2] = 21'b000000000001011001000;
        x_t[3] = 21'b000000000001010100100;
        x_t[4] = 21'b000000000000110001100;
        x_t[5] = 21'b111111111111001011100;
        x_t[6] = 21'b111111111101101101101;
        x_t[7] = 21'b000000000001000111111;
        x_t[8] = 21'b000000000010011100011;
        x_t[9] = 21'b000000000011001111010;
        x_t[10] = 21'b000000000100011100011;
        x_t[11] = 21'b000000000010011000000;
        x_t[12] = 21'b000000000010001111110;
        x_t[13] = 21'b000000000001010011111;
        x_t[14] = 21'b000000000010100100000;
        x_t[15] = 21'b000000000011101100101;
        x_t[16] = 21'b000000000011111110010;
        x_t[17] = 21'b000000000100001001011;
        x_t[18] = 21'b000000000100010101000;
        x_t[19] = 21'b000000000100100010110;
        x_t[20] = 21'b000000000010110111010;
        x_t[21] = 21'b111111111110111010110;
        x_t[22] = 21'b111111111110011101110;
        x_t[23] = 21'b111111111101100010011;
        x_t[24] = 21'b111111111101111000111;
        x_t[25] = 21'b111111111101111101110;
        x_t[26] = 21'b111111111101011010101;
        x_t[27] = 21'b111111111101100000100;
        x_t[28] = 21'b111111111111010100010;
        x_t[29] = 21'b111111111111100111110;
        x_t[30] = 21'b111111111110001000110;
        x_t[31] = 21'b111111111101101101000;
        x_t[32] = 21'b111111111111001100000;
        x_t[33] = 21'b111111111110100000011;
        x_t[34] = 21'b111111111101010111111;
        x_t[35] = 21'b111111111101101010000;
        x_t[36] = 21'b111111111100110010111;
        x_t[37] = 21'b111111111100111001001;
        x_t[38] = 21'b111111111111110101010;
        x_t[39] = 21'b111111111110110100110;
        x_t[40] = 21'b000000000000111110110;
        x_t[41] = 21'b111111111001110101100;
        x_t[42] = 21'b000000000000111111101;
        x_t[43] = 21'b000000000011101101111;
        x_t[44] = 21'b111111111111101000000;
        x_t[45] = 21'b000000000101000100100;
        x_t[46] = 21'b000000000010001101111;
        x_t[47] = 21'b000000000011001000110;
        x_t[48] = 21'b000000000010101110011;
        x_t[49] = 21'b000000000100101101100;
        x_t[50] = 21'b000000000100111100110;
        x_t[51] = 21'b000000000101100111110;
        x_t[52] = 21'b000000000101001001110;
        x_t[53] = 21'b000000000100111011110;
        x_t[54] = 21'b000000000100110000101;
        x_t[55] = 21'b000000000011101010101;
        x_t[56] = 21'b000000000011110001110;
        x_t[57] = 21'b000000000101111101100;
        x_t[58] = 21'b000000000101101101110;
        x_t[59] = 21'b000000000101111110001;
        x_t[60] = 21'b000000000101000101000;
        x_t[61] = 21'b000000000110011001001;
        x_t[62] = 21'b000000000011111010111;
        x_t[63] = 21'b000000000011001010110;
        
        h_t_prev[0] = 21'b000000000001000100011;
        h_t_prev[1] = 21'b000000000001111100111;
        h_t_prev[2] = 21'b000000000001011001000;
        h_t_prev[3] = 21'b000000000001010100100;
        h_t_prev[4] = 21'b000000000000110001100;
        h_t_prev[5] = 21'b111111111111001011100;
        h_t_prev[6] = 21'b111111111101101101101;
        h_t_prev[7] = 21'b000000000001000111111;
        h_t_prev[8] = 21'b000000000010011100011;
        h_t_prev[9] = 21'b000000000011001111010;
        h_t_prev[10] = 21'b000000000100011100011;
        h_t_prev[11] = 21'b000000000010011000000;
        h_t_prev[12] = 21'b000000000010001111110;
        h_t_prev[13] = 21'b000000000001010011111;
        h_t_prev[14] = 21'b000000000010100100000;
        h_t_prev[15] = 21'b000000000011101100101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 96 timeout!");
                $fdisplay(fd_cycles, "Test Vector  96: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  96: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 96");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 97
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111111000100001;
        x_t[1] = 21'b111111111111000111111;
        x_t[2] = 21'b111111111101111001101;
        x_t[3] = 21'b111111111110100110100;
        x_t[4] = 21'b111111111110111101011;
        x_t[5] = 21'b111111111110011111001;
        x_t[6] = 21'b111111111111001011000;
        x_t[7] = 21'b111111111111111011100;
        x_t[8] = 21'b111111111110010000001;
        x_t[9] = 21'b111111111101010111100;
        x_t[10] = 21'b111111111101101101110;
        x_t[11] = 21'b111111111101100110010;
        x_t[12] = 21'b111111111110111101000;
        x_t[13] = 21'b000000000000101011000;
        x_t[14] = 21'b111111111110010001110;
        x_t[15] = 21'b111111111110010111111;
        x_t[16] = 21'b111111111101110001101;
        x_t[17] = 21'b111111111101011100001;
        x_t[18] = 21'b111111111110100100000;
        x_t[19] = 21'b111111111110000110111;
        x_t[20] = 21'b000000000000101101101;
        x_t[21] = 21'b000000000001100000100;
        x_t[22] = 21'b000000000001011111010;
        x_t[23] = 21'b000000000000111001001;
        x_t[24] = 21'b000000000000111011110;
        x_t[25] = 21'b000000000000110101001;
        x_t[26] = 21'b000000000000011000110;
        x_t[27] = 21'b111111111111011010010;
        x_t[28] = 21'b111111111110111011001;
        x_t[29] = 21'b000000000000001101010;
        x_t[30] = 21'b000000000001000000001;
        x_t[31] = 21'b111111111111100100110;
        x_t[32] = 21'b000000000000010000001;
        x_t[33] = 21'b111111111111010011010;
        x_t[34] = 21'b111111111111001111000;
        x_t[35] = 21'b111111111111100000100;
        x_t[36] = 21'b111111111111000011000;
        x_t[37] = 21'b111111111111001011111;
        x_t[38] = 21'b111111111111111111011;
        x_t[39] = 21'b000000000010010001010;
        x_t[40] = 21'b111111111111110010101;
        x_t[41] = 21'b000000000110000111011;
        x_t[42] = 21'b111111111111001111000;
        x_t[43] = 21'b000000000010000000001;
        x_t[44] = 21'b111111111110000011011;
        x_t[45] = 21'b000000000010101001110;
        x_t[46] = 21'b111111111100111101001;
        x_t[47] = 21'b111111111110010100011;
        x_t[48] = 21'b111111111110011010000;
        x_t[49] = 21'b111111111110101000010;
        x_t[50] = 21'b111111111110010110000;
        x_t[51] = 21'b111111111110110101000;
        x_t[52] = 21'b111111111110111010110;
        x_t[53] = 21'b111111111111110011010;
        x_t[54] = 21'b000000000000101111000;
        x_t[55] = 21'b111111111101010000101;
        x_t[56] = 21'b111111111110100111000;
        x_t[57] = 21'b111111111111000010001;
        x_t[58] = 21'b111111111111001111011;
        x_t[59] = 21'b111111111111001000000;
        x_t[60] = 21'b111111111111001001100;
        x_t[61] = 21'b111111111110100000010;
        x_t[62] = 21'b111111111110100110101;
        x_t[63] = 21'b000000000000001101100;
        
        h_t_prev[0] = 21'b111111111111000100001;
        h_t_prev[1] = 21'b111111111111000111111;
        h_t_prev[2] = 21'b111111111101111001101;
        h_t_prev[3] = 21'b111111111110100110100;
        h_t_prev[4] = 21'b111111111110111101011;
        h_t_prev[5] = 21'b111111111110011111001;
        h_t_prev[6] = 21'b111111111111001011000;
        h_t_prev[7] = 21'b111111111111111011100;
        h_t_prev[8] = 21'b111111111110010000001;
        h_t_prev[9] = 21'b111111111101010111100;
        h_t_prev[10] = 21'b111111111101101101110;
        h_t_prev[11] = 21'b111111111101100110010;
        h_t_prev[12] = 21'b111111111110111101000;
        h_t_prev[13] = 21'b000000000000101011000;
        h_t_prev[14] = 21'b111111111110010001110;
        h_t_prev[15] = 21'b111111111110010111111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 97 timeout!");
                $fdisplay(fd_cycles, "Test Vector  97: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  97: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 97");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 98
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b000000000000000100010;
        x_t[1] = 21'b111111111111111101101;
        x_t[2] = 21'b111111111110101010010;
        x_t[3] = 21'b111111111111100101011;
        x_t[4] = 21'b111111111111100000110;
        x_t[5] = 21'b111111111110111010111;
        x_t[6] = 21'b111111111111010001010;
        x_t[7] = 21'b000000000000011010000;
        x_t[8] = 21'b111111111110011111101;
        x_t[9] = 21'b111111111101110000100;
        x_t[10] = 21'b111111111110011001111;
        x_t[11] = 21'b111111111110011001010;
        x_t[12] = 21'b111111111111001110101;
        x_t[13] = 21'b000000000001011010101;
        x_t[14] = 21'b111111111110010111000;
        x_t[15] = 21'b111111111110000011100;
        x_t[16] = 21'b111111111101101100110;
        x_t[17] = 21'b111111111101101111111;
        x_t[18] = 21'b111111111110101001010;
        x_t[19] = 21'b111111111101110110011;
        x_t[20] = 21'b000000000000010100100;
        x_t[21] = 21'b000000000001100110000;
        x_t[22] = 21'b000000000001011000111;
        x_t[23] = 21'b000000000000110011010;
        x_t[24] = 21'b000000000000111110110;
        x_t[25] = 21'b000000000000111011010;
        x_t[26] = 21'b000000000000001100001;
        x_t[27] = 21'b111111111111100010001;
        x_t[28] = 21'b111111111110101011011;
        x_t[29] = 21'b000000000000001101010;
        x_t[30] = 21'b000000000001000000001;
        x_t[31] = 21'b111111111111110010000;
        x_t[32] = 21'b000000000000010000001;
        x_t[33] = 21'b111111111111001010000;
        x_t[34] = 21'b111111111111000101011;
        x_t[35] = 21'b111111111111000111110;
        x_t[36] = 21'b111111111110110100000;
        x_t[37] = 21'b111111111110100011001;
        x_t[38] = 21'b111111111111110101010;
        x_t[39] = 21'b000000000001000111110;
        x_t[40] = 21'b111111111110110110111;
        x_t[41] = 21'b000000000000101011101;
        x_t[42] = 21'b111111111110011001101;
        x_t[43] = 21'b000000000001001001011;
        x_t[44] = 21'b111111111101000000011;
        x_t[45] = 21'b000000000001001100111;
        x_t[46] = 21'b111111111100001001010;
        x_t[47] = 21'b111111111101010011110;
        x_t[48] = 21'b111111111101010111010;
        x_t[49] = 21'b111111111101110000101;
        x_t[50] = 21'b111111111101101011001;
        x_t[51] = 21'b111111111101111111111;
        x_t[52] = 21'b111111111110000010100;
        x_t[53] = 21'b111111111110011111110;
        x_t[54] = 21'b111111111110110111001;
        x_t[55] = 21'b111111111011111010011;
        x_t[56] = 21'b111111111101010001000;
        x_t[57] = 21'b111111111101111001101;
        x_t[58] = 21'b111111111110011011000;
        x_t[59] = 21'b111111111110100000100;
        x_t[60] = 21'b111111111110001100001;
        x_t[61] = 21'b111111111101111111001;
        x_t[62] = 21'b111111111110011111010;
        x_t[63] = 21'b111111111111101010010;
        
        h_t_prev[0] = 21'b000000000000000100010;
        h_t_prev[1] = 21'b111111111111111101101;
        h_t_prev[2] = 21'b111111111110101010010;
        h_t_prev[3] = 21'b111111111111100101011;
        h_t_prev[4] = 21'b111111111111100000110;
        h_t_prev[5] = 21'b111111111110111010111;
        h_t_prev[6] = 21'b111111111111010001010;
        h_t_prev[7] = 21'b000000000000011010000;
        h_t_prev[8] = 21'b111111111110011111101;
        h_t_prev[9] = 21'b111111111101110000100;
        h_t_prev[10] = 21'b111111111110011001111;
        h_t_prev[11] = 21'b111111111110011001010;
        h_t_prev[12] = 21'b111111111111001110101;
        h_t_prev[13] = 21'b000000000001011010101;
        h_t_prev[14] = 21'b111111111110010111000;
        h_t_prev[15] = 21'b111111111110000011100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 98 timeout!");
                $fdisplay(fd_cycles, "Test Vector  98: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  98: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 98");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 99
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111110111010010;
        x_t[1] = 21'b111111111110100101100;
        x_t[2] = 21'b111111111101011100100;
        x_t[3] = 21'b111111111110011100111;
        x_t[4] = 21'b111111111110010101000;
        x_t[5] = 21'b111111111101101101001;
        x_t[6] = 21'b111111111101101101101;
        x_t[7] = 21'b111111111110101010000;
        x_t[8] = 21'b111111111100101001000;
        x_t[9] = 21'b111111111100000010010;
        x_t[10] = 21'b111111111100101110010;
        x_t[11] = 21'b111111111100011110111;
        x_t[12] = 21'b111111111100111100010;
        x_t[13] = 21'b111111111110001110010;
        x_t[14] = 21'b111111111100101101101;
        x_t[15] = 21'b111111111011111010010;
        x_t[16] = 21'b111111111011100001111;
        x_t[17] = 21'b111111111011111001011;
        x_t[18] = 21'b111111111100011011000;
        x_t[19] = 21'b111111111011001100001;
        x_t[20] = 21'b111111111100101101000;
        x_t[21] = 21'b000000000001001010011;
        x_t[22] = 21'b000000000000110110000;
        x_t[23] = 21'b000000000000010110010;
        x_t[24] = 21'b000000000000001011000;
        x_t[25] = 21'b000000000000000110100;
        x_t[26] = 21'b111111111111001100110;
        x_t[27] = 21'b111111111110101011001;
        x_t[28] = 21'b111111111101111100001;
        x_t[29] = 21'b111111111111011011011;
        x_t[30] = 21'b000000000000000101101;
        x_t[31] = 21'b111111111110101011000;
        x_t[32] = 21'b111111111110110101011;
        x_t[33] = 21'b111111111101110110110;
        x_t[34] = 21'b111111111110000010110;
        x_t[35] = 21'b111111111110000111101;
        x_t[36] = 21'b111111111101011111101;
        x_t[37] = 21'b111111111101011101110;
        x_t[38] = 21'b111111111111000010110;
        x_t[39] = 21'b111111111110010000000;
        x_t[40] = 21'b111111111110000110000;
        x_t[41] = 21'b111111111100010101100;
        x_t[42] = 21'b111111111101110000001;
        x_t[43] = 21'b111111111110101111110;
        x_t[44] = 21'b111111111100001110001;
        x_t[45] = 21'b111111111100000111111;
        x_t[46] = 21'b111111111011001011001;
        x_t[47] = 21'b111111111011100001011;
        x_t[48] = 21'b111111111011001101001;
        x_t[49] = 21'b111111111011001001111;
        x_t[50] = 21'b111111111011000100111;
        x_t[51] = 21'b111111111011000011101;
        x_t[52] = 21'b111111111010101011101;
        x_t[53] = 21'b111111111010011010001;
        x_t[54] = 21'b111111111001101101100;
        x_t[55] = 21'b111111111010010111001;
        x_t[56] = 21'b111111111011010000001;
        x_t[57] = 21'b111111111011100000001;
        x_t[58] = 21'b111111111011011111100;
        x_t[59] = 21'b111111111011001011011;
        x_t[60] = 21'b111111111100111011101;
        x_t[61] = 21'b111111111100011011110;
        x_t[62] = 21'b111111111101000110100;
        x_t[63] = 21'b111111111110000000101;
        
        h_t_prev[0] = 21'b111111111110111010010;
        h_t_prev[1] = 21'b111111111110100101100;
        h_t_prev[2] = 21'b111111111101011100100;
        h_t_prev[3] = 21'b111111111110011100111;
        h_t_prev[4] = 21'b111111111110010101000;
        h_t_prev[5] = 21'b111111111101101101001;
        h_t_prev[6] = 21'b111111111101101101101;
        h_t_prev[7] = 21'b111111111110101010000;
        h_t_prev[8] = 21'b111111111100101001000;
        h_t_prev[9] = 21'b111111111100000010010;
        h_t_prev[10] = 21'b111111111100101110010;
        h_t_prev[11] = 21'b111111111100011110111;
        h_t_prev[12] = 21'b111111111100111100010;
        h_t_prev[13] = 21'b111111111110001110010;
        h_t_prev[14] = 21'b111111111100101101101;
        h_t_prev[15] = 21'b111111111011111010010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 99 timeout!");
                $fdisplay(fd_cycles, "Test Vector  99: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  99: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 99");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 100
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 21'b111111111110111010010;
        x_t[1] = 21'b111111111110010010000;
        x_t[2] = 21'b111111111100101100000;
        x_t[3] = 21'b111111111101110110010;
        x_t[4] = 21'b111111111101110110101;
        x_t[5] = 21'b111111111101001011111;
        x_t[6] = 21'b111111111101100001010;
        x_t[7] = 21'b111111111111001000101;
        x_t[8] = 21'b111111111011110101100;
        x_t[9] = 21'b111111111011000001001;
        x_t[10] = 21'b111111111011010110001;
        x_t[11] = 21'b111111111011000011010;
        x_t[12] = 21'b111111111011000111001;
        x_t[13] = 21'b111111111100010011101;
        x_t[14] = 21'b111111111100111000001;
        x_t[15] = 21'b111111111011010110101;
        x_t[16] = 21'b111111111010010010101;
        x_t[17] = 21'b111111111010010110101;
        x_t[18] = 21'b111111111010111100001;
        x_t[19] = 21'b111111111001001000011;
        x_t[20] = 21'b111111111010010000101;
        x_t[21] = 21'b000000000010001010000;
        x_t[22] = 21'b000000000010010010000;
        x_t[23] = 21'b000000000001100100101;
        x_t[24] = 21'b000000000001011010010;
        x_t[25] = 21'b000000000001001110000;
        x_t[26] = 21'b000000000000110010001;
        x_t[27] = 21'b000000000000001001100;
        x_t[28] = 21'b111111111111001010111;
        x_t[29] = 21'b000000000001001011101;
        x_t[30] = 21'b000000000001000100001;
        x_t[31] = 21'b111111111111101101101;
        x_t[32] = 21'b111111111111110000011;
        x_t[33] = 21'b111111111111010111111;
        x_t[34] = 21'b111111111111101011100;
        x_t[35] = 21'b111111111111101010011;
        x_t[36] = 21'b111111111111011011111;
        x_t[37] = 21'b111111111111010000000;
        x_t[38] = 21'b000000000000101100110;
        x_t[39] = 21'b111111111111101000010;
        x_t[40] = 21'b000000000000011000110;
        x_t[41] = 21'b111111111111000011011;
        x_t[42] = 21'b000000000000011100000;
        x_t[43] = 21'b111111111011010100010;
        x_t[44] = 21'b111111111101001011100;
        x_t[45] = 21'b111111111000011111110;
        x_t[46] = 21'b111111111011101010001;
        x_t[47] = 21'b111111111011011100011;
        x_t[48] = 21'b111111111010110101010;
        x_t[49] = 21'b111111111010010010010;
        x_t[50] = 21'b111111111010000010011;
        x_t[51] = 21'b111111111001110110010;
        x_t[52] = 21'b111111111001110011011;
        x_t[53] = 21'b111111111001000001000;
        x_t[54] = 21'b111111111000010011101;
        x_t[55] = 21'b111111111001111000111;
        x_t[56] = 21'b111111111010001111101;
        x_t[57] = 21'b111111111010100000010;
        x_t[58] = 21'b111111111010010101010;
        x_t[59] = 21'b111111111001111100011;
        x_t[60] = 21'b111111111011101111000;
        x_t[61] = 21'b111111111011000000110;
        x_t[62] = 21'b111111111011101101110;
        x_t[63] = 21'b111111111101010100101;
        
        h_t_prev[0] = 21'b111111111110111010010;
        h_t_prev[1] = 21'b111111111110010010000;
        h_t_prev[2] = 21'b111111111100101100000;
        h_t_prev[3] = 21'b111111111101110110010;
        h_t_prev[4] = 21'b111111111101110110101;
        h_t_prev[5] = 21'b111111111101001011111;
        h_t_prev[6] = 21'b111111111101100001010;
        h_t_prev[7] = 21'b111111111111001000101;
        h_t_prev[8] = 21'b111111111011110101100;
        h_t_prev[9] = 21'b111111111011000001001;
        h_t_prev[10] = 21'b111111111011010110001;
        h_t_prev[11] = 21'b111111111011000011010;
        h_t_prev[12] = 21'b111111111011000111001;
        h_t_prev[13] = 21'b111111111100010011101;
        h_t_prev[14] = 21'b111111111100111000001;
        h_t_prev[15] = 21'b111111111011010110101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 100 timeout!");
                $fdisplay(fd_cycles, "Test Vector 100: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector 100: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b %021b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 100");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Write summary to cycles file
    $fdisplay(fd_cycles, "");
    $fdisplay(fd_cycles, "==========================================================");
    $fdisplay(fd_cycles, "SUMMARY");
    $fdisplay(fd_cycles, "==========================================================");
    $fdisplay(fd_cycles, "Total Test Vectors: %0d", 100);
    $fdisplay(fd_cycles, "Total Cycles:       %0d", total_cycles);
    $fdisplay(fd_cycles, "Average Cycles:     %.2f", real'(total_cycles) / 100);
    $fdisplay(fd_cycles, "Total Time:         %.2f us @ 100MHz", total_cycles * 0.01);
    $fdisplay(fd_cycles, "Average Time:       %.2f us @ 100MHz", (total_cycles * 0.01) / 100);
    $fdisplay(fd_cycles, "Throughput:         %.2f computations/ms @ 100MHz", 100000.0 / (real'(total_cycles) / 100));
    $fdisplay(fd_cycles, "==========================================================");
    
    $fclose(fd_output);
    $fclose(fd_cycles);
    
    $display("");
    $display("==========================================================");
    $display("Simulation Complete");
    $display("==========================================================");
    $display("Test Vectors:   %0d", 100);
    $display("Total Cycles:   %0d", total_cycles);
    $display("Average Cycles: %.2f", real'(total_cycles) / 100);
    $display("==========================================================");
    $display("Output file:    output_d64_h16_dw21_fb11_np1.txt");
    $display("Cycles file:    cycles_d64_h16_dw21_fb11_np1.txt");
    $display("==========================================================");
    
    $finish;
end

endmodule