
`timescale 1ns / 1ps
// GRU Cell Implementation (Fixed-Point Qm.f)
// d = 256 (input features), h = 8 (hidden units)
// WIDTH = INT_WIDTH + FRAC_WIDTH

module gru #(
    parameter int INT_WIDTH  = 4,
    parameter int FRAC_WIDTH = 5,
    parameter int WIDTH      = INT_WIDTH + FRAC_WIDTH
)(
    input  logic                     clk,
    input  logic                     reset,

    // Inputs (d=256)
        input  logic signed [WIDTH-1:0]  x_0,
    input  logic signed [WIDTH-1:0]  x_1,
    input  logic signed [WIDTH-1:0]  x_2,
    input  logic signed [WIDTH-1:0]  x_3,
    input  logic signed [WIDTH-1:0]  x_4,
    input  logic signed [WIDTH-1:0]  x_5,
    input  logic signed [WIDTH-1:0]  x_6,
    input  logic signed [WIDTH-1:0]  x_7,
    input  logic signed [WIDTH-1:0]  x_8,
    input  logic signed [WIDTH-1:0]  x_9,
    input  logic signed [WIDTH-1:0]  x_10,
    input  logic signed [WIDTH-1:0]  x_11,
    input  logic signed [WIDTH-1:0]  x_12,
    input  logic signed [WIDTH-1:0]  x_13,
    input  logic signed [WIDTH-1:0]  x_14,
    input  logic signed [WIDTH-1:0]  x_15,
    input  logic signed [WIDTH-1:0]  x_16,
    input  logic signed [WIDTH-1:0]  x_17,
    input  logic signed [WIDTH-1:0]  x_18,
    input  logic signed [WIDTH-1:0]  x_19,
    input  logic signed [WIDTH-1:0]  x_20,
    input  logic signed [WIDTH-1:0]  x_21,
    input  logic signed [WIDTH-1:0]  x_22,
    input  logic signed [WIDTH-1:0]  x_23,
    input  logic signed [WIDTH-1:0]  x_24,
    input  logic signed [WIDTH-1:0]  x_25,
    input  logic signed [WIDTH-1:0]  x_26,
    input  logic signed [WIDTH-1:0]  x_27,
    input  logic signed [WIDTH-1:0]  x_28,
    input  logic signed [WIDTH-1:0]  x_29,
    input  logic signed [WIDTH-1:0]  x_30,
    input  logic signed [WIDTH-1:0]  x_31,
    input  logic signed [WIDTH-1:0]  x_32,
    input  logic signed [WIDTH-1:0]  x_33,
    input  logic signed [WIDTH-1:0]  x_34,
    input  logic signed [WIDTH-1:0]  x_35,
    input  logic signed [WIDTH-1:0]  x_36,
    input  logic signed [WIDTH-1:0]  x_37,
    input  logic signed [WIDTH-1:0]  x_38,
    input  logic signed [WIDTH-1:0]  x_39,
    input  logic signed [WIDTH-1:0]  x_40,
    input  logic signed [WIDTH-1:0]  x_41,
    input  logic signed [WIDTH-1:0]  x_42,
    input  logic signed [WIDTH-1:0]  x_43,
    input  logic signed [WIDTH-1:0]  x_44,
    input  logic signed [WIDTH-1:0]  x_45,
    input  logic signed [WIDTH-1:0]  x_46,
    input  logic signed [WIDTH-1:0]  x_47,
    input  logic signed [WIDTH-1:0]  x_48,
    input  logic signed [WIDTH-1:0]  x_49,
    input  logic signed [WIDTH-1:0]  x_50,
    input  logic signed [WIDTH-1:0]  x_51,
    input  logic signed [WIDTH-1:0]  x_52,
    input  logic signed [WIDTH-1:0]  x_53,
    input  logic signed [WIDTH-1:0]  x_54,
    input  logic signed [WIDTH-1:0]  x_55,
    input  logic signed [WIDTH-1:0]  x_56,
    input  logic signed [WIDTH-1:0]  x_57,
    input  logic signed [WIDTH-1:0]  x_58,
    input  logic signed [WIDTH-1:0]  x_59,
    input  logic signed [WIDTH-1:0]  x_60,
    input  logic signed [WIDTH-1:0]  x_61,
    input  logic signed [WIDTH-1:0]  x_62,
    input  logic signed [WIDTH-1:0]  x_63,
    input  logic signed [WIDTH-1:0]  x_64,
    input  logic signed [WIDTH-1:0]  x_65,
    input  logic signed [WIDTH-1:0]  x_66,
    input  logic signed [WIDTH-1:0]  x_67,
    input  logic signed [WIDTH-1:0]  x_68,
    input  logic signed [WIDTH-1:0]  x_69,
    input  logic signed [WIDTH-1:0]  x_70,
    input  logic signed [WIDTH-1:0]  x_71,
    input  logic signed [WIDTH-1:0]  x_72,
    input  logic signed [WIDTH-1:0]  x_73,
    input  logic signed [WIDTH-1:0]  x_74,
    input  logic signed [WIDTH-1:0]  x_75,
    input  logic signed [WIDTH-1:0]  x_76,
    input  logic signed [WIDTH-1:0]  x_77,
    input  logic signed [WIDTH-1:0]  x_78,
    input  logic signed [WIDTH-1:0]  x_79,
    input  logic signed [WIDTH-1:0]  x_80,
    input  logic signed [WIDTH-1:0]  x_81,
    input  logic signed [WIDTH-1:0]  x_82,
    input  logic signed [WIDTH-1:0]  x_83,
    input  logic signed [WIDTH-1:0]  x_84,
    input  logic signed [WIDTH-1:0]  x_85,
    input  logic signed [WIDTH-1:0]  x_86,
    input  logic signed [WIDTH-1:0]  x_87,
    input  logic signed [WIDTH-1:0]  x_88,
    input  logic signed [WIDTH-1:0]  x_89,
    input  logic signed [WIDTH-1:0]  x_90,
    input  logic signed [WIDTH-1:0]  x_91,
    input  logic signed [WIDTH-1:0]  x_92,
    input  logic signed [WIDTH-1:0]  x_93,
    input  logic signed [WIDTH-1:0]  x_94,
    input  logic signed [WIDTH-1:0]  x_95,
    input  logic signed [WIDTH-1:0]  x_96,
    input  logic signed [WIDTH-1:0]  x_97,
    input  logic signed [WIDTH-1:0]  x_98,
    input  logic signed [WIDTH-1:0]  x_99,
    input  logic signed [WIDTH-1:0]  x_100,
    input  logic signed [WIDTH-1:0]  x_101,
    input  logic signed [WIDTH-1:0]  x_102,
    input  logic signed [WIDTH-1:0]  x_103,
    input  logic signed [WIDTH-1:0]  x_104,
    input  logic signed [WIDTH-1:0]  x_105,
    input  logic signed [WIDTH-1:0]  x_106,
    input  logic signed [WIDTH-1:0]  x_107,
    input  logic signed [WIDTH-1:0]  x_108,
    input  logic signed [WIDTH-1:0]  x_109,
    input  logic signed [WIDTH-1:0]  x_110,
    input  logic signed [WIDTH-1:0]  x_111,
    input  logic signed [WIDTH-1:0]  x_112,
    input  logic signed [WIDTH-1:0]  x_113,
    input  logic signed [WIDTH-1:0]  x_114,
    input  logic signed [WIDTH-1:0]  x_115,
    input  logic signed [WIDTH-1:0]  x_116,
    input  logic signed [WIDTH-1:0]  x_117,
    input  logic signed [WIDTH-1:0]  x_118,
    input  logic signed [WIDTH-1:0]  x_119,
    input  logic signed [WIDTH-1:0]  x_120,
    input  logic signed [WIDTH-1:0]  x_121,
    input  logic signed [WIDTH-1:0]  x_122,
    input  logic signed [WIDTH-1:0]  x_123,
    input  logic signed [WIDTH-1:0]  x_124,
    input  logic signed [WIDTH-1:0]  x_125,
    input  logic signed [WIDTH-1:0]  x_126,
    input  logic signed [WIDTH-1:0]  x_127,
    input  logic signed [WIDTH-1:0]  x_128,
    input  logic signed [WIDTH-1:0]  x_129,
    input  logic signed [WIDTH-1:0]  x_130,
    input  logic signed [WIDTH-1:0]  x_131,
    input  logic signed [WIDTH-1:0]  x_132,
    input  logic signed [WIDTH-1:0]  x_133,
    input  logic signed [WIDTH-1:0]  x_134,
    input  logic signed [WIDTH-1:0]  x_135,
    input  logic signed [WIDTH-1:0]  x_136,
    input  logic signed [WIDTH-1:0]  x_137,
    input  logic signed [WIDTH-1:0]  x_138,
    input  logic signed [WIDTH-1:0]  x_139,
    input  logic signed [WIDTH-1:0]  x_140,
    input  logic signed [WIDTH-1:0]  x_141,
    input  logic signed [WIDTH-1:0]  x_142,
    input  logic signed [WIDTH-1:0]  x_143,
    input  logic signed [WIDTH-1:0]  x_144,
    input  logic signed [WIDTH-1:0]  x_145,
    input  logic signed [WIDTH-1:0]  x_146,
    input  logic signed [WIDTH-1:0]  x_147,
    input  logic signed [WIDTH-1:0]  x_148,
    input  logic signed [WIDTH-1:0]  x_149,
    input  logic signed [WIDTH-1:0]  x_150,
    input  logic signed [WIDTH-1:0]  x_151,
    input  logic signed [WIDTH-1:0]  x_152,
    input  logic signed [WIDTH-1:0]  x_153,
    input  logic signed [WIDTH-1:0]  x_154,
    input  logic signed [WIDTH-1:0]  x_155,
    input  logic signed [WIDTH-1:0]  x_156,
    input  logic signed [WIDTH-1:0]  x_157,
    input  logic signed [WIDTH-1:0]  x_158,
    input  logic signed [WIDTH-1:0]  x_159,
    input  logic signed [WIDTH-1:0]  x_160,
    input  logic signed [WIDTH-1:0]  x_161,
    input  logic signed [WIDTH-1:0]  x_162,
    input  logic signed [WIDTH-1:0]  x_163,
    input  logic signed [WIDTH-1:0]  x_164,
    input  logic signed [WIDTH-1:0]  x_165,
    input  logic signed [WIDTH-1:0]  x_166,
    input  logic signed [WIDTH-1:0]  x_167,
    input  logic signed [WIDTH-1:0]  x_168,
    input  logic signed [WIDTH-1:0]  x_169,
    input  logic signed [WIDTH-1:0]  x_170,
    input  logic signed [WIDTH-1:0]  x_171,
    input  logic signed [WIDTH-1:0]  x_172,
    input  logic signed [WIDTH-1:0]  x_173,
    input  logic signed [WIDTH-1:0]  x_174,
    input  logic signed [WIDTH-1:0]  x_175,
    input  logic signed [WIDTH-1:0]  x_176,
    input  logic signed [WIDTH-1:0]  x_177,
    input  logic signed [WIDTH-1:0]  x_178,
    input  logic signed [WIDTH-1:0]  x_179,
    input  logic signed [WIDTH-1:0]  x_180,
    input  logic signed [WIDTH-1:0]  x_181,
    input  logic signed [WIDTH-1:0]  x_182,
    input  logic signed [WIDTH-1:0]  x_183,
    input  logic signed [WIDTH-1:0]  x_184,
    input  logic signed [WIDTH-1:0]  x_185,
    input  logic signed [WIDTH-1:0]  x_186,
    input  logic signed [WIDTH-1:0]  x_187,
    input  logic signed [WIDTH-1:0]  x_188,
    input  logic signed [WIDTH-1:0]  x_189,
    input  logic signed [WIDTH-1:0]  x_190,
    input  logic signed [WIDTH-1:0]  x_191,
    input  logic signed [WIDTH-1:0]  x_192,
    input  logic signed [WIDTH-1:0]  x_193,
    input  logic signed [WIDTH-1:0]  x_194,
    input  logic signed [WIDTH-1:0]  x_195,
    input  logic signed [WIDTH-1:0]  x_196,
    input  logic signed [WIDTH-1:0]  x_197,
    input  logic signed [WIDTH-1:0]  x_198,
    input  logic signed [WIDTH-1:0]  x_199,
    input  logic signed [WIDTH-1:0]  x_200,
    input  logic signed [WIDTH-1:0]  x_201,
    input  logic signed [WIDTH-1:0]  x_202,
    input  logic signed [WIDTH-1:0]  x_203,
    input  logic signed [WIDTH-1:0]  x_204,
    input  logic signed [WIDTH-1:0]  x_205,
    input  logic signed [WIDTH-1:0]  x_206,
    input  logic signed [WIDTH-1:0]  x_207,
    input  logic signed [WIDTH-1:0]  x_208,
    input  logic signed [WIDTH-1:0]  x_209,
    input  logic signed [WIDTH-1:0]  x_210,
    input  logic signed [WIDTH-1:0]  x_211,
    input  logic signed [WIDTH-1:0]  x_212,
    input  logic signed [WIDTH-1:0]  x_213,
    input  logic signed [WIDTH-1:0]  x_214,
    input  logic signed [WIDTH-1:0]  x_215,
    input  logic signed [WIDTH-1:0]  x_216,
    input  logic signed [WIDTH-1:0]  x_217,
    input  logic signed [WIDTH-1:0]  x_218,
    input  logic signed [WIDTH-1:0]  x_219,
    input  logic signed [WIDTH-1:0]  x_220,
    input  logic signed [WIDTH-1:0]  x_221,
    input  logic signed [WIDTH-1:0]  x_222,
    input  logic signed [WIDTH-1:0]  x_223,
    input  logic signed [WIDTH-1:0]  x_224,
    input  logic signed [WIDTH-1:0]  x_225,
    input  logic signed [WIDTH-1:0]  x_226,
    input  logic signed [WIDTH-1:0]  x_227,
    input  logic signed [WIDTH-1:0]  x_228,
    input  logic signed [WIDTH-1:0]  x_229,
    input  logic signed [WIDTH-1:0]  x_230,
    input  logic signed [WIDTH-1:0]  x_231,
    input  logic signed [WIDTH-1:0]  x_232,
    input  logic signed [WIDTH-1:0]  x_233,
    input  logic signed [WIDTH-1:0]  x_234,
    input  logic signed [WIDTH-1:0]  x_235,
    input  logic signed [WIDTH-1:0]  x_236,
    input  logic signed [WIDTH-1:0]  x_237,
    input  logic signed [WIDTH-1:0]  x_238,
    input  logic signed [WIDTH-1:0]  x_239,
    input  logic signed [WIDTH-1:0]  x_240,
    input  logic signed [WIDTH-1:0]  x_241,
    input  logic signed [WIDTH-1:0]  x_242,
    input  logic signed [WIDTH-1:0]  x_243,
    input  logic signed [WIDTH-1:0]  x_244,
    input  logic signed [WIDTH-1:0]  x_245,
    input  logic signed [WIDTH-1:0]  x_246,
    input  logic signed [WIDTH-1:0]  x_247,
    input  logic signed [WIDTH-1:0]  x_248,
    input  logic signed [WIDTH-1:0]  x_249,
    input  logic signed [WIDTH-1:0]  x_250,
    input  logic signed [WIDTH-1:0]  x_251,
    input  logic signed [WIDTH-1:0]  x_252,
    input  logic signed [WIDTH-1:0]  x_253,
    input  logic signed [WIDTH-1:0]  x_254,
    input  logic signed [WIDTH-1:0]  x_255,

    // Previous hidden state (h=8)
        input  logic signed [WIDTH-1:0]  h_0,
    input  logic signed [WIDTH-1:0]  h_1,
    input  logic signed [WIDTH-1:0]  h_2,
    input  logic signed [WIDTH-1:0]  h_3,
    input  logic signed [WIDTH-1:0]  h_4,
    input  logic signed [WIDTH-1:0]  h_5,
    input  logic signed [WIDTH-1:0]  h_6,
    input  logic signed [WIDTH-1:0]  h_7,

    // Input weights (h×d for each gate)
    input  logic signed [WIDTH-1:0]  w_ir_0_0, w_ir_0_1, w_ir_0_2, w_ir_0_3, w_ir_0_4, w_ir_0_5, w_ir_0_6, w_ir_0_7, w_ir_0_8, w_ir_0_9, w_ir_0_10, w_ir_0_11, w_ir_0_12, w_ir_0_13, w_ir_0_14, w_ir_0_15, w_ir_0_16, w_ir_0_17, w_ir_0_18, w_ir_0_19, w_ir_0_20, w_ir_0_21, w_ir_0_22, w_ir_0_23, w_ir_0_24, w_ir_0_25, w_ir_0_26, w_ir_0_27, w_ir_0_28, w_ir_0_29, w_ir_0_30, w_ir_0_31, w_ir_0_32, w_ir_0_33, w_ir_0_34, w_ir_0_35, w_ir_0_36, w_ir_0_37, w_ir_0_38, w_ir_0_39, w_ir_0_40, w_ir_0_41, w_ir_0_42, w_ir_0_43, w_ir_0_44, w_ir_0_45, w_ir_0_46, w_ir_0_47, w_ir_0_48, w_ir_0_49, w_ir_0_50, w_ir_0_51, w_ir_0_52, w_ir_0_53, w_ir_0_54, w_ir_0_55, w_ir_0_56, w_ir_0_57, w_ir_0_58, w_ir_0_59, w_ir_0_60, w_ir_0_61, w_ir_0_62, w_ir_0_63, w_ir_0_64, w_ir_0_65, w_ir_0_66, w_ir_0_67, w_ir_0_68, w_ir_0_69, w_ir_0_70, w_ir_0_71, w_ir_0_72, w_ir_0_73, w_ir_0_74, w_ir_0_75, w_ir_0_76, w_ir_0_77, w_ir_0_78, w_ir_0_79, w_ir_0_80, w_ir_0_81, w_ir_0_82, w_ir_0_83, w_ir_0_84, w_ir_0_85, w_ir_0_86, w_ir_0_87, w_ir_0_88, w_ir_0_89, w_ir_0_90, w_ir_0_91, w_ir_0_92, w_ir_0_93, w_ir_0_94, w_ir_0_95, w_ir_0_96, w_ir_0_97, w_ir_0_98, w_ir_0_99, w_ir_0_100, w_ir_0_101, w_ir_0_102, w_ir_0_103, w_ir_0_104, w_ir_0_105, w_ir_0_106, w_ir_0_107, w_ir_0_108, w_ir_0_109, w_ir_0_110, w_ir_0_111, w_ir_0_112, w_ir_0_113, w_ir_0_114, w_ir_0_115, w_ir_0_116, w_ir_0_117, w_ir_0_118, w_ir_0_119, w_ir_0_120, w_ir_0_121, w_ir_0_122, w_ir_0_123, w_ir_0_124, w_ir_0_125, w_ir_0_126, w_ir_0_127, w_ir_0_128, w_ir_0_129, w_ir_0_130, w_ir_0_131, w_ir_0_132, w_ir_0_133, w_ir_0_134, w_ir_0_135, w_ir_0_136, w_ir_0_137, w_ir_0_138, w_ir_0_139, w_ir_0_140, w_ir_0_141, w_ir_0_142, w_ir_0_143, w_ir_0_144, w_ir_0_145, w_ir_0_146, w_ir_0_147, w_ir_0_148, w_ir_0_149, w_ir_0_150, w_ir_0_151, w_ir_0_152, w_ir_0_153, w_ir_0_154, w_ir_0_155, w_ir_0_156, w_ir_0_157, w_ir_0_158, w_ir_0_159, w_ir_0_160, w_ir_0_161, w_ir_0_162, w_ir_0_163, w_ir_0_164, w_ir_0_165, w_ir_0_166, w_ir_0_167, w_ir_0_168, w_ir_0_169, w_ir_0_170, w_ir_0_171, w_ir_0_172, w_ir_0_173, w_ir_0_174, w_ir_0_175, w_ir_0_176, w_ir_0_177, w_ir_0_178, w_ir_0_179, w_ir_0_180, w_ir_0_181, w_ir_0_182, w_ir_0_183, w_ir_0_184, w_ir_0_185, w_ir_0_186, w_ir_0_187, w_ir_0_188, w_ir_0_189, w_ir_0_190, w_ir_0_191, w_ir_0_192, w_ir_0_193, w_ir_0_194, w_ir_0_195, w_ir_0_196, w_ir_0_197, w_ir_0_198, w_ir_0_199, w_ir_0_200, w_ir_0_201, w_ir_0_202, w_ir_0_203, w_ir_0_204, w_ir_0_205, w_ir_0_206, w_ir_0_207, w_ir_0_208, w_ir_0_209, w_ir_0_210, w_ir_0_211, w_ir_0_212, w_ir_0_213, w_ir_0_214, w_ir_0_215, w_ir_0_216, w_ir_0_217, w_ir_0_218, w_ir_0_219, w_ir_0_220, w_ir_0_221, w_ir_0_222, w_ir_0_223, w_ir_0_224, w_ir_0_225, w_ir_0_226, w_ir_0_227, w_ir_0_228, w_ir_0_229, w_ir_0_230, w_ir_0_231, w_ir_0_232, w_ir_0_233, w_ir_0_234, w_ir_0_235, w_ir_0_236, w_ir_0_237, w_ir_0_238, w_ir_0_239, w_ir_0_240, w_ir_0_241, w_ir_0_242, w_ir_0_243, w_ir_0_244, w_ir_0_245, w_ir_0_246, w_ir_0_247, w_ir_0_248, w_ir_0_249, w_ir_0_250, w_ir_0_251, w_ir_0_252, w_ir_0_253, w_ir_0_254, w_ir_0_255, w_ir_1_0, w_ir_1_1, w_ir_1_2, w_ir_1_3, w_ir_1_4, w_ir_1_5, w_ir_1_6, w_ir_1_7, w_ir_1_8, w_ir_1_9, w_ir_1_10, w_ir_1_11, w_ir_1_12, w_ir_1_13, w_ir_1_14, w_ir_1_15, w_ir_1_16, w_ir_1_17, w_ir_1_18, w_ir_1_19, w_ir_1_20, w_ir_1_21, w_ir_1_22, w_ir_1_23, w_ir_1_24, w_ir_1_25, w_ir_1_26, w_ir_1_27, w_ir_1_28, w_ir_1_29, w_ir_1_30, w_ir_1_31, w_ir_1_32, w_ir_1_33, w_ir_1_34, w_ir_1_35, w_ir_1_36, w_ir_1_37, w_ir_1_38, w_ir_1_39, w_ir_1_40, w_ir_1_41, w_ir_1_42, w_ir_1_43, w_ir_1_44, w_ir_1_45, w_ir_1_46, w_ir_1_47, w_ir_1_48, w_ir_1_49, w_ir_1_50, w_ir_1_51, w_ir_1_52, w_ir_1_53, w_ir_1_54, w_ir_1_55, w_ir_1_56, w_ir_1_57, w_ir_1_58, w_ir_1_59, w_ir_1_60, w_ir_1_61, w_ir_1_62, w_ir_1_63, w_ir_1_64, w_ir_1_65, w_ir_1_66, w_ir_1_67, w_ir_1_68, w_ir_1_69, w_ir_1_70, w_ir_1_71, w_ir_1_72, w_ir_1_73, w_ir_1_74, w_ir_1_75, w_ir_1_76, w_ir_1_77, w_ir_1_78, w_ir_1_79, w_ir_1_80, w_ir_1_81, w_ir_1_82, w_ir_1_83, w_ir_1_84, w_ir_1_85, w_ir_1_86, w_ir_1_87, w_ir_1_88, w_ir_1_89, w_ir_1_90, w_ir_1_91, w_ir_1_92, w_ir_1_93, w_ir_1_94, w_ir_1_95, w_ir_1_96, w_ir_1_97, w_ir_1_98, w_ir_1_99, w_ir_1_100, w_ir_1_101, w_ir_1_102, w_ir_1_103, w_ir_1_104, w_ir_1_105, w_ir_1_106, w_ir_1_107, w_ir_1_108, w_ir_1_109, w_ir_1_110, w_ir_1_111, w_ir_1_112, w_ir_1_113, w_ir_1_114, w_ir_1_115, w_ir_1_116, w_ir_1_117, w_ir_1_118, w_ir_1_119, w_ir_1_120, w_ir_1_121, w_ir_1_122, w_ir_1_123, w_ir_1_124, w_ir_1_125, w_ir_1_126, w_ir_1_127, w_ir_1_128, w_ir_1_129, w_ir_1_130, w_ir_1_131, w_ir_1_132, w_ir_1_133, w_ir_1_134, w_ir_1_135, w_ir_1_136, w_ir_1_137, w_ir_1_138, w_ir_1_139, w_ir_1_140, w_ir_1_141, w_ir_1_142, w_ir_1_143, w_ir_1_144, w_ir_1_145, w_ir_1_146, w_ir_1_147, w_ir_1_148, w_ir_1_149, w_ir_1_150, w_ir_1_151, w_ir_1_152, w_ir_1_153, w_ir_1_154, w_ir_1_155, w_ir_1_156, w_ir_1_157, w_ir_1_158, w_ir_1_159, w_ir_1_160, w_ir_1_161, w_ir_1_162, w_ir_1_163, w_ir_1_164, w_ir_1_165, w_ir_1_166, w_ir_1_167, w_ir_1_168, w_ir_1_169, w_ir_1_170, w_ir_1_171, w_ir_1_172, w_ir_1_173, w_ir_1_174, w_ir_1_175, w_ir_1_176, w_ir_1_177, w_ir_1_178, w_ir_1_179, w_ir_1_180, w_ir_1_181, w_ir_1_182, w_ir_1_183, w_ir_1_184, w_ir_1_185, w_ir_1_186, w_ir_1_187, w_ir_1_188, w_ir_1_189, w_ir_1_190, w_ir_1_191, w_ir_1_192, w_ir_1_193, w_ir_1_194, w_ir_1_195, w_ir_1_196, w_ir_1_197, w_ir_1_198, w_ir_1_199, w_ir_1_200, w_ir_1_201, w_ir_1_202, w_ir_1_203, w_ir_1_204, w_ir_1_205, w_ir_1_206, w_ir_1_207, w_ir_1_208, w_ir_1_209, w_ir_1_210, w_ir_1_211, w_ir_1_212, w_ir_1_213, w_ir_1_214, w_ir_1_215, w_ir_1_216, w_ir_1_217, w_ir_1_218, w_ir_1_219, w_ir_1_220, w_ir_1_221, w_ir_1_222, w_ir_1_223, w_ir_1_224, w_ir_1_225, w_ir_1_226, w_ir_1_227, w_ir_1_228, w_ir_1_229, w_ir_1_230, w_ir_1_231, w_ir_1_232, w_ir_1_233, w_ir_1_234, w_ir_1_235, w_ir_1_236, w_ir_1_237, w_ir_1_238, w_ir_1_239, w_ir_1_240, w_ir_1_241, w_ir_1_242, w_ir_1_243, w_ir_1_244, w_ir_1_245, w_ir_1_246, w_ir_1_247, w_ir_1_248, w_ir_1_249, w_ir_1_250, w_ir_1_251, w_ir_1_252, w_ir_1_253, w_ir_1_254, w_ir_1_255, w_ir_2_0, w_ir_2_1, w_ir_2_2, w_ir_2_3, w_ir_2_4, w_ir_2_5, w_ir_2_6, w_ir_2_7, w_ir_2_8, w_ir_2_9, w_ir_2_10, w_ir_2_11, w_ir_2_12, w_ir_2_13, w_ir_2_14, w_ir_2_15, w_ir_2_16, w_ir_2_17, w_ir_2_18, w_ir_2_19, w_ir_2_20, w_ir_2_21, w_ir_2_22, w_ir_2_23, w_ir_2_24, w_ir_2_25, w_ir_2_26, w_ir_2_27, w_ir_2_28, w_ir_2_29, w_ir_2_30, w_ir_2_31, w_ir_2_32, w_ir_2_33, w_ir_2_34, w_ir_2_35, w_ir_2_36, w_ir_2_37, w_ir_2_38, w_ir_2_39, w_ir_2_40, w_ir_2_41, w_ir_2_42, w_ir_2_43, w_ir_2_44, w_ir_2_45, w_ir_2_46, w_ir_2_47, w_ir_2_48, w_ir_2_49, w_ir_2_50, w_ir_2_51, w_ir_2_52, w_ir_2_53, w_ir_2_54, w_ir_2_55, w_ir_2_56, w_ir_2_57, w_ir_2_58, w_ir_2_59, w_ir_2_60, w_ir_2_61, w_ir_2_62, w_ir_2_63, w_ir_2_64, w_ir_2_65, w_ir_2_66, w_ir_2_67, w_ir_2_68, w_ir_2_69, w_ir_2_70, w_ir_2_71, w_ir_2_72, w_ir_2_73, w_ir_2_74, w_ir_2_75, w_ir_2_76, w_ir_2_77, w_ir_2_78, w_ir_2_79, w_ir_2_80, w_ir_2_81, w_ir_2_82, w_ir_2_83, w_ir_2_84, w_ir_2_85, w_ir_2_86, w_ir_2_87, w_ir_2_88, w_ir_2_89, w_ir_2_90, w_ir_2_91, w_ir_2_92, w_ir_2_93, w_ir_2_94, w_ir_2_95, w_ir_2_96, w_ir_2_97, w_ir_2_98, w_ir_2_99, w_ir_2_100, w_ir_2_101, w_ir_2_102, w_ir_2_103, w_ir_2_104, w_ir_2_105, w_ir_2_106, w_ir_2_107, w_ir_2_108, w_ir_2_109, w_ir_2_110, w_ir_2_111, w_ir_2_112, w_ir_2_113, w_ir_2_114, w_ir_2_115, w_ir_2_116, w_ir_2_117, w_ir_2_118, w_ir_2_119, w_ir_2_120, w_ir_2_121, w_ir_2_122, w_ir_2_123, w_ir_2_124, w_ir_2_125, w_ir_2_126, w_ir_2_127, w_ir_2_128, w_ir_2_129, w_ir_2_130, w_ir_2_131, w_ir_2_132, w_ir_2_133, w_ir_2_134, w_ir_2_135, w_ir_2_136, w_ir_2_137, w_ir_2_138, w_ir_2_139, w_ir_2_140, w_ir_2_141, w_ir_2_142, w_ir_2_143, w_ir_2_144, w_ir_2_145, w_ir_2_146, w_ir_2_147, w_ir_2_148, w_ir_2_149, w_ir_2_150, w_ir_2_151, w_ir_2_152, w_ir_2_153, w_ir_2_154, w_ir_2_155, w_ir_2_156, w_ir_2_157, w_ir_2_158, w_ir_2_159, w_ir_2_160, w_ir_2_161, w_ir_2_162, w_ir_2_163, w_ir_2_164, w_ir_2_165, w_ir_2_166, w_ir_2_167, w_ir_2_168, w_ir_2_169, w_ir_2_170, w_ir_2_171, w_ir_2_172, w_ir_2_173, w_ir_2_174, w_ir_2_175, w_ir_2_176, w_ir_2_177, w_ir_2_178, w_ir_2_179, w_ir_2_180, w_ir_2_181, w_ir_2_182, w_ir_2_183, w_ir_2_184, w_ir_2_185, w_ir_2_186, w_ir_2_187, w_ir_2_188, w_ir_2_189, w_ir_2_190, w_ir_2_191, w_ir_2_192, w_ir_2_193, w_ir_2_194, w_ir_2_195, w_ir_2_196, w_ir_2_197, w_ir_2_198, w_ir_2_199, w_ir_2_200, w_ir_2_201, w_ir_2_202, w_ir_2_203, w_ir_2_204, w_ir_2_205, w_ir_2_206, w_ir_2_207, w_ir_2_208, w_ir_2_209, w_ir_2_210, w_ir_2_211, w_ir_2_212, w_ir_2_213, w_ir_2_214, w_ir_2_215, w_ir_2_216, w_ir_2_217, w_ir_2_218, w_ir_2_219, w_ir_2_220, w_ir_2_221, w_ir_2_222, w_ir_2_223, w_ir_2_224, w_ir_2_225, w_ir_2_226, w_ir_2_227, w_ir_2_228, w_ir_2_229, w_ir_2_230, w_ir_2_231, w_ir_2_232, w_ir_2_233, w_ir_2_234, w_ir_2_235, w_ir_2_236, w_ir_2_237, w_ir_2_238, w_ir_2_239, w_ir_2_240, w_ir_2_241, w_ir_2_242, w_ir_2_243, w_ir_2_244, w_ir_2_245, w_ir_2_246, w_ir_2_247, w_ir_2_248, w_ir_2_249, w_ir_2_250, w_ir_2_251, w_ir_2_252, w_ir_2_253, w_ir_2_254, w_ir_2_255, w_ir_3_0, w_ir_3_1, w_ir_3_2, w_ir_3_3, w_ir_3_4, w_ir_3_5, w_ir_3_6, w_ir_3_7, w_ir_3_8, w_ir_3_9, w_ir_3_10, w_ir_3_11, w_ir_3_12, w_ir_3_13, w_ir_3_14, w_ir_3_15, w_ir_3_16, w_ir_3_17, w_ir_3_18, w_ir_3_19, w_ir_3_20, w_ir_3_21, w_ir_3_22, w_ir_3_23, w_ir_3_24, w_ir_3_25, w_ir_3_26, w_ir_3_27, w_ir_3_28, w_ir_3_29, w_ir_3_30, w_ir_3_31, w_ir_3_32, w_ir_3_33, w_ir_3_34, w_ir_3_35, w_ir_3_36, w_ir_3_37, w_ir_3_38, w_ir_3_39, w_ir_3_40, w_ir_3_41, w_ir_3_42, w_ir_3_43, w_ir_3_44, w_ir_3_45, w_ir_3_46, w_ir_3_47, w_ir_3_48, w_ir_3_49, w_ir_3_50, w_ir_3_51, w_ir_3_52, w_ir_3_53, w_ir_3_54, w_ir_3_55, w_ir_3_56, w_ir_3_57, w_ir_3_58, w_ir_3_59, w_ir_3_60, w_ir_3_61, w_ir_3_62, w_ir_3_63, w_ir_3_64, w_ir_3_65, w_ir_3_66, w_ir_3_67, w_ir_3_68, w_ir_3_69, w_ir_3_70, w_ir_3_71, w_ir_3_72, w_ir_3_73, w_ir_3_74, w_ir_3_75, w_ir_3_76, w_ir_3_77, w_ir_3_78, w_ir_3_79, w_ir_3_80, w_ir_3_81, w_ir_3_82, w_ir_3_83, w_ir_3_84, w_ir_3_85, w_ir_3_86, w_ir_3_87, w_ir_3_88, w_ir_3_89, w_ir_3_90, w_ir_3_91, w_ir_3_92, w_ir_3_93, w_ir_3_94, w_ir_3_95, w_ir_3_96, w_ir_3_97, w_ir_3_98, w_ir_3_99, w_ir_3_100, w_ir_3_101, w_ir_3_102, w_ir_3_103, w_ir_3_104, w_ir_3_105, w_ir_3_106, w_ir_3_107, w_ir_3_108, w_ir_3_109, w_ir_3_110, w_ir_3_111, w_ir_3_112, w_ir_3_113, w_ir_3_114, w_ir_3_115, w_ir_3_116, w_ir_3_117, w_ir_3_118, w_ir_3_119, w_ir_3_120, w_ir_3_121, w_ir_3_122, w_ir_3_123, w_ir_3_124, w_ir_3_125, w_ir_3_126, w_ir_3_127, w_ir_3_128, w_ir_3_129, w_ir_3_130, w_ir_3_131, w_ir_3_132, w_ir_3_133, w_ir_3_134, w_ir_3_135, w_ir_3_136, w_ir_3_137, w_ir_3_138, w_ir_3_139, w_ir_3_140, w_ir_3_141, w_ir_3_142, w_ir_3_143, w_ir_3_144, w_ir_3_145, w_ir_3_146, w_ir_3_147, w_ir_3_148, w_ir_3_149, w_ir_3_150, w_ir_3_151, w_ir_3_152, w_ir_3_153, w_ir_3_154, w_ir_3_155, w_ir_3_156, w_ir_3_157, w_ir_3_158, w_ir_3_159, w_ir_3_160, w_ir_3_161, w_ir_3_162, w_ir_3_163, w_ir_3_164, w_ir_3_165, w_ir_3_166, w_ir_3_167, w_ir_3_168, w_ir_3_169, w_ir_3_170, w_ir_3_171, w_ir_3_172, w_ir_3_173, w_ir_3_174, w_ir_3_175, w_ir_3_176, w_ir_3_177, w_ir_3_178, w_ir_3_179, w_ir_3_180, w_ir_3_181, w_ir_3_182, w_ir_3_183, w_ir_3_184, w_ir_3_185, w_ir_3_186, w_ir_3_187, w_ir_3_188, w_ir_3_189, w_ir_3_190, w_ir_3_191, w_ir_3_192, w_ir_3_193, w_ir_3_194, w_ir_3_195, w_ir_3_196, w_ir_3_197, w_ir_3_198, w_ir_3_199, w_ir_3_200, w_ir_3_201, w_ir_3_202, w_ir_3_203, w_ir_3_204, w_ir_3_205, w_ir_3_206, w_ir_3_207, w_ir_3_208, w_ir_3_209, w_ir_3_210, w_ir_3_211, w_ir_3_212, w_ir_3_213, w_ir_3_214, w_ir_3_215, w_ir_3_216, w_ir_3_217, w_ir_3_218, w_ir_3_219, w_ir_3_220, w_ir_3_221, w_ir_3_222, w_ir_3_223, w_ir_3_224, w_ir_3_225, w_ir_3_226, w_ir_3_227, w_ir_3_228, w_ir_3_229, w_ir_3_230, w_ir_3_231, w_ir_3_232, w_ir_3_233, w_ir_3_234, w_ir_3_235, w_ir_3_236, w_ir_3_237, w_ir_3_238, w_ir_3_239, w_ir_3_240, w_ir_3_241, w_ir_3_242, w_ir_3_243, w_ir_3_244, w_ir_3_245, w_ir_3_246, w_ir_3_247, w_ir_3_248, w_ir_3_249, w_ir_3_250, w_ir_3_251, w_ir_3_252, w_ir_3_253, w_ir_3_254, w_ir_3_255, w_ir_4_0, w_ir_4_1, w_ir_4_2, w_ir_4_3, w_ir_4_4, w_ir_4_5, w_ir_4_6, w_ir_4_7, w_ir_4_8, w_ir_4_9, w_ir_4_10, w_ir_4_11, w_ir_4_12, w_ir_4_13, w_ir_4_14, w_ir_4_15, w_ir_4_16, w_ir_4_17, w_ir_4_18, w_ir_4_19, w_ir_4_20, w_ir_4_21, w_ir_4_22, w_ir_4_23, w_ir_4_24, w_ir_4_25, w_ir_4_26, w_ir_4_27, w_ir_4_28, w_ir_4_29, w_ir_4_30, w_ir_4_31, w_ir_4_32, w_ir_4_33, w_ir_4_34, w_ir_4_35, w_ir_4_36, w_ir_4_37, w_ir_4_38, w_ir_4_39, w_ir_4_40, w_ir_4_41, w_ir_4_42, w_ir_4_43, w_ir_4_44, w_ir_4_45, w_ir_4_46, w_ir_4_47, w_ir_4_48, w_ir_4_49, w_ir_4_50, w_ir_4_51, w_ir_4_52, w_ir_4_53, w_ir_4_54, w_ir_4_55, w_ir_4_56, w_ir_4_57, w_ir_4_58, w_ir_4_59, w_ir_4_60, w_ir_4_61, w_ir_4_62, w_ir_4_63, w_ir_4_64, w_ir_4_65, w_ir_4_66, w_ir_4_67, w_ir_4_68, w_ir_4_69, w_ir_4_70, w_ir_4_71, w_ir_4_72, w_ir_4_73, w_ir_4_74, w_ir_4_75, w_ir_4_76, w_ir_4_77, w_ir_4_78, w_ir_4_79, w_ir_4_80, w_ir_4_81, w_ir_4_82, w_ir_4_83, w_ir_4_84, w_ir_4_85, w_ir_4_86, w_ir_4_87, w_ir_4_88, w_ir_4_89, w_ir_4_90, w_ir_4_91, w_ir_4_92, w_ir_4_93, w_ir_4_94, w_ir_4_95, w_ir_4_96, w_ir_4_97, w_ir_4_98, w_ir_4_99, w_ir_4_100, w_ir_4_101, w_ir_4_102, w_ir_4_103, w_ir_4_104, w_ir_4_105, w_ir_4_106, w_ir_4_107, w_ir_4_108, w_ir_4_109, w_ir_4_110, w_ir_4_111, w_ir_4_112, w_ir_4_113, w_ir_4_114, w_ir_4_115, w_ir_4_116, w_ir_4_117, w_ir_4_118, w_ir_4_119, w_ir_4_120, w_ir_4_121, w_ir_4_122, w_ir_4_123, w_ir_4_124, w_ir_4_125, w_ir_4_126, w_ir_4_127, w_ir_4_128, w_ir_4_129, w_ir_4_130, w_ir_4_131, w_ir_4_132, w_ir_4_133, w_ir_4_134, w_ir_4_135, w_ir_4_136, w_ir_4_137, w_ir_4_138, w_ir_4_139, w_ir_4_140, w_ir_4_141, w_ir_4_142, w_ir_4_143, w_ir_4_144, w_ir_4_145, w_ir_4_146, w_ir_4_147, w_ir_4_148, w_ir_4_149, w_ir_4_150, w_ir_4_151, w_ir_4_152, w_ir_4_153, w_ir_4_154, w_ir_4_155, w_ir_4_156, w_ir_4_157, w_ir_4_158, w_ir_4_159, w_ir_4_160, w_ir_4_161, w_ir_4_162, w_ir_4_163, w_ir_4_164, w_ir_4_165, w_ir_4_166, w_ir_4_167, w_ir_4_168, w_ir_4_169, w_ir_4_170, w_ir_4_171, w_ir_4_172, w_ir_4_173, w_ir_4_174, w_ir_4_175, w_ir_4_176, w_ir_4_177, w_ir_4_178, w_ir_4_179, w_ir_4_180, w_ir_4_181, w_ir_4_182, w_ir_4_183, w_ir_4_184, w_ir_4_185, w_ir_4_186, w_ir_4_187, w_ir_4_188, w_ir_4_189, w_ir_4_190, w_ir_4_191, w_ir_4_192, w_ir_4_193, w_ir_4_194, w_ir_4_195, w_ir_4_196, w_ir_4_197, w_ir_4_198, w_ir_4_199, w_ir_4_200, w_ir_4_201, w_ir_4_202, w_ir_4_203, w_ir_4_204, w_ir_4_205, w_ir_4_206, w_ir_4_207, w_ir_4_208, w_ir_4_209, w_ir_4_210, w_ir_4_211, w_ir_4_212, w_ir_4_213, w_ir_4_214, w_ir_4_215, w_ir_4_216, w_ir_4_217, w_ir_4_218, w_ir_4_219, w_ir_4_220, w_ir_4_221, w_ir_4_222, w_ir_4_223, w_ir_4_224, w_ir_4_225, w_ir_4_226, w_ir_4_227, w_ir_4_228, w_ir_4_229, w_ir_4_230, w_ir_4_231, w_ir_4_232, w_ir_4_233, w_ir_4_234, w_ir_4_235, w_ir_4_236, w_ir_4_237, w_ir_4_238, w_ir_4_239, w_ir_4_240, w_ir_4_241, w_ir_4_242, w_ir_4_243, w_ir_4_244, w_ir_4_245, w_ir_4_246, w_ir_4_247, w_ir_4_248, w_ir_4_249, w_ir_4_250, w_ir_4_251, w_ir_4_252, w_ir_4_253, w_ir_4_254, w_ir_4_255, w_ir_5_0, w_ir_5_1, w_ir_5_2, w_ir_5_3, w_ir_5_4, w_ir_5_5, w_ir_5_6, w_ir_5_7, w_ir_5_8, w_ir_5_9, w_ir_5_10, w_ir_5_11, w_ir_5_12, w_ir_5_13, w_ir_5_14, w_ir_5_15, w_ir_5_16, w_ir_5_17, w_ir_5_18, w_ir_5_19, w_ir_5_20, w_ir_5_21, w_ir_5_22, w_ir_5_23, w_ir_5_24, w_ir_5_25, w_ir_5_26, w_ir_5_27, w_ir_5_28, w_ir_5_29, w_ir_5_30, w_ir_5_31, w_ir_5_32, w_ir_5_33, w_ir_5_34, w_ir_5_35, w_ir_5_36, w_ir_5_37, w_ir_5_38, w_ir_5_39, w_ir_5_40, w_ir_5_41, w_ir_5_42, w_ir_5_43, w_ir_5_44, w_ir_5_45, w_ir_5_46, w_ir_5_47, w_ir_5_48, w_ir_5_49, w_ir_5_50, w_ir_5_51, w_ir_5_52, w_ir_5_53, w_ir_5_54, w_ir_5_55, w_ir_5_56, w_ir_5_57, w_ir_5_58, w_ir_5_59, w_ir_5_60, w_ir_5_61, w_ir_5_62, w_ir_5_63, w_ir_5_64, w_ir_5_65, w_ir_5_66, w_ir_5_67, w_ir_5_68, w_ir_5_69, w_ir_5_70, w_ir_5_71, w_ir_5_72, w_ir_5_73, w_ir_5_74, w_ir_5_75, w_ir_5_76, w_ir_5_77, w_ir_5_78, w_ir_5_79, w_ir_5_80, w_ir_5_81, w_ir_5_82, w_ir_5_83, w_ir_5_84, w_ir_5_85, w_ir_5_86, w_ir_5_87, w_ir_5_88, w_ir_5_89, w_ir_5_90, w_ir_5_91, w_ir_5_92, w_ir_5_93, w_ir_5_94, w_ir_5_95, w_ir_5_96, w_ir_5_97, w_ir_5_98, w_ir_5_99, w_ir_5_100, w_ir_5_101, w_ir_5_102, w_ir_5_103, w_ir_5_104, w_ir_5_105, w_ir_5_106, w_ir_5_107, w_ir_5_108, w_ir_5_109, w_ir_5_110, w_ir_5_111, w_ir_5_112, w_ir_5_113, w_ir_5_114, w_ir_5_115, w_ir_5_116, w_ir_5_117, w_ir_5_118, w_ir_5_119, w_ir_5_120, w_ir_5_121, w_ir_5_122, w_ir_5_123, w_ir_5_124, w_ir_5_125, w_ir_5_126, w_ir_5_127, w_ir_5_128, w_ir_5_129, w_ir_5_130, w_ir_5_131, w_ir_5_132, w_ir_5_133, w_ir_5_134, w_ir_5_135, w_ir_5_136, w_ir_5_137, w_ir_5_138, w_ir_5_139, w_ir_5_140, w_ir_5_141, w_ir_5_142, w_ir_5_143, w_ir_5_144, w_ir_5_145, w_ir_5_146, w_ir_5_147, w_ir_5_148, w_ir_5_149, w_ir_5_150, w_ir_5_151, w_ir_5_152, w_ir_5_153, w_ir_5_154, w_ir_5_155, w_ir_5_156, w_ir_5_157, w_ir_5_158, w_ir_5_159, w_ir_5_160, w_ir_5_161, w_ir_5_162, w_ir_5_163, w_ir_5_164, w_ir_5_165, w_ir_5_166, w_ir_5_167, w_ir_5_168, w_ir_5_169, w_ir_5_170, w_ir_5_171, w_ir_5_172, w_ir_5_173, w_ir_5_174, w_ir_5_175, w_ir_5_176, w_ir_5_177, w_ir_5_178, w_ir_5_179, w_ir_5_180, w_ir_5_181, w_ir_5_182, w_ir_5_183, w_ir_5_184, w_ir_5_185, w_ir_5_186, w_ir_5_187, w_ir_5_188, w_ir_5_189, w_ir_5_190, w_ir_5_191, w_ir_5_192, w_ir_5_193, w_ir_5_194, w_ir_5_195, w_ir_5_196, w_ir_5_197, w_ir_5_198, w_ir_5_199, w_ir_5_200, w_ir_5_201, w_ir_5_202, w_ir_5_203, w_ir_5_204, w_ir_5_205, w_ir_5_206, w_ir_5_207, w_ir_5_208, w_ir_5_209, w_ir_5_210, w_ir_5_211, w_ir_5_212, w_ir_5_213, w_ir_5_214, w_ir_5_215, w_ir_5_216, w_ir_5_217, w_ir_5_218, w_ir_5_219, w_ir_5_220, w_ir_5_221, w_ir_5_222, w_ir_5_223, w_ir_5_224, w_ir_5_225, w_ir_5_226, w_ir_5_227, w_ir_5_228, w_ir_5_229, w_ir_5_230, w_ir_5_231, w_ir_5_232, w_ir_5_233, w_ir_5_234, w_ir_5_235, w_ir_5_236, w_ir_5_237, w_ir_5_238, w_ir_5_239, w_ir_5_240, w_ir_5_241, w_ir_5_242, w_ir_5_243, w_ir_5_244, w_ir_5_245, w_ir_5_246, w_ir_5_247, w_ir_5_248, w_ir_5_249, w_ir_5_250, w_ir_5_251, w_ir_5_252, w_ir_5_253, w_ir_5_254, w_ir_5_255, w_ir_6_0, w_ir_6_1, w_ir_6_2, w_ir_6_3, w_ir_6_4, w_ir_6_5, w_ir_6_6, w_ir_6_7, w_ir_6_8, w_ir_6_9, w_ir_6_10, w_ir_6_11, w_ir_6_12, w_ir_6_13, w_ir_6_14, w_ir_6_15, w_ir_6_16, w_ir_6_17, w_ir_6_18, w_ir_6_19, w_ir_6_20, w_ir_6_21, w_ir_6_22, w_ir_6_23, w_ir_6_24, w_ir_6_25, w_ir_6_26, w_ir_6_27, w_ir_6_28, w_ir_6_29, w_ir_6_30, w_ir_6_31, w_ir_6_32, w_ir_6_33, w_ir_6_34, w_ir_6_35, w_ir_6_36, w_ir_6_37, w_ir_6_38, w_ir_6_39, w_ir_6_40, w_ir_6_41, w_ir_6_42, w_ir_6_43, w_ir_6_44, w_ir_6_45, w_ir_6_46, w_ir_6_47, w_ir_6_48, w_ir_6_49, w_ir_6_50, w_ir_6_51, w_ir_6_52, w_ir_6_53, w_ir_6_54, w_ir_6_55, w_ir_6_56, w_ir_6_57, w_ir_6_58, w_ir_6_59, w_ir_6_60, w_ir_6_61, w_ir_6_62, w_ir_6_63, w_ir_6_64, w_ir_6_65, w_ir_6_66, w_ir_6_67, w_ir_6_68, w_ir_6_69, w_ir_6_70, w_ir_6_71, w_ir_6_72, w_ir_6_73, w_ir_6_74, w_ir_6_75, w_ir_6_76, w_ir_6_77, w_ir_6_78, w_ir_6_79, w_ir_6_80, w_ir_6_81, w_ir_6_82, w_ir_6_83, w_ir_6_84, w_ir_6_85, w_ir_6_86, w_ir_6_87, w_ir_6_88, w_ir_6_89, w_ir_6_90, w_ir_6_91, w_ir_6_92, w_ir_6_93, w_ir_6_94, w_ir_6_95, w_ir_6_96, w_ir_6_97, w_ir_6_98, w_ir_6_99, w_ir_6_100, w_ir_6_101, w_ir_6_102, w_ir_6_103, w_ir_6_104, w_ir_6_105, w_ir_6_106, w_ir_6_107, w_ir_6_108, w_ir_6_109, w_ir_6_110, w_ir_6_111, w_ir_6_112, w_ir_6_113, w_ir_6_114, w_ir_6_115, w_ir_6_116, w_ir_6_117, w_ir_6_118, w_ir_6_119, w_ir_6_120, w_ir_6_121, w_ir_6_122, w_ir_6_123, w_ir_6_124, w_ir_6_125, w_ir_6_126, w_ir_6_127, w_ir_6_128, w_ir_6_129, w_ir_6_130, w_ir_6_131, w_ir_6_132, w_ir_6_133, w_ir_6_134, w_ir_6_135, w_ir_6_136, w_ir_6_137, w_ir_6_138, w_ir_6_139, w_ir_6_140, w_ir_6_141, w_ir_6_142, w_ir_6_143, w_ir_6_144, w_ir_6_145, w_ir_6_146, w_ir_6_147, w_ir_6_148, w_ir_6_149, w_ir_6_150, w_ir_6_151, w_ir_6_152, w_ir_6_153, w_ir_6_154, w_ir_6_155, w_ir_6_156, w_ir_6_157, w_ir_6_158, w_ir_6_159, w_ir_6_160, w_ir_6_161, w_ir_6_162, w_ir_6_163, w_ir_6_164, w_ir_6_165, w_ir_6_166, w_ir_6_167, w_ir_6_168, w_ir_6_169, w_ir_6_170, w_ir_6_171, w_ir_6_172, w_ir_6_173, w_ir_6_174, w_ir_6_175, w_ir_6_176, w_ir_6_177, w_ir_6_178, w_ir_6_179, w_ir_6_180, w_ir_6_181, w_ir_6_182, w_ir_6_183, w_ir_6_184, w_ir_6_185, w_ir_6_186, w_ir_6_187, w_ir_6_188, w_ir_6_189, w_ir_6_190, w_ir_6_191, w_ir_6_192, w_ir_6_193, w_ir_6_194, w_ir_6_195, w_ir_6_196, w_ir_6_197, w_ir_6_198, w_ir_6_199, w_ir_6_200, w_ir_6_201, w_ir_6_202, w_ir_6_203, w_ir_6_204, w_ir_6_205, w_ir_6_206, w_ir_6_207, w_ir_6_208, w_ir_6_209, w_ir_6_210, w_ir_6_211, w_ir_6_212, w_ir_6_213, w_ir_6_214, w_ir_6_215, w_ir_6_216, w_ir_6_217, w_ir_6_218, w_ir_6_219, w_ir_6_220, w_ir_6_221, w_ir_6_222, w_ir_6_223, w_ir_6_224, w_ir_6_225, w_ir_6_226, w_ir_6_227, w_ir_6_228, w_ir_6_229, w_ir_6_230, w_ir_6_231, w_ir_6_232, w_ir_6_233, w_ir_6_234, w_ir_6_235, w_ir_6_236, w_ir_6_237, w_ir_6_238, w_ir_6_239, w_ir_6_240, w_ir_6_241, w_ir_6_242, w_ir_6_243, w_ir_6_244, w_ir_6_245, w_ir_6_246, w_ir_6_247, w_ir_6_248, w_ir_6_249, w_ir_6_250, w_ir_6_251, w_ir_6_252, w_ir_6_253, w_ir_6_254, w_ir_6_255, w_ir_7_0, w_ir_7_1, w_ir_7_2, w_ir_7_3, w_ir_7_4, w_ir_7_5, w_ir_7_6, w_ir_7_7, w_ir_7_8, w_ir_7_9, w_ir_7_10, w_ir_7_11, w_ir_7_12, w_ir_7_13, w_ir_7_14, w_ir_7_15, w_ir_7_16, w_ir_7_17, w_ir_7_18, w_ir_7_19, w_ir_7_20, w_ir_7_21, w_ir_7_22, w_ir_7_23, w_ir_7_24, w_ir_7_25, w_ir_7_26, w_ir_7_27, w_ir_7_28, w_ir_7_29, w_ir_7_30, w_ir_7_31, w_ir_7_32, w_ir_7_33, w_ir_7_34, w_ir_7_35, w_ir_7_36, w_ir_7_37, w_ir_7_38, w_ir_7_39, w_ir_7_40, w_ir_7_41, w_ir_7_42, w_ir_7_43, w_ir_7_44, w_ir_7_45, w_ir_7_46, w_ir_7_47, w_ir_7_48, w_ir_7_49, w_ir_7_50, w_ir_7_51, w_ir_7_52, w_ir_7_53, w_ir_7_54, w_ir_7_55, w_ir_7_56, w_ir_7_57, w_ir_7_58, w_ir_7_59, w_ir_7_60, w_ir_7_61, w_ir_7_62, w_ir_7_63, w_ir_7_64, w_ir_7_65, w_ir_7_66, w_ir_7_67, w_ir_7_68, w_ir_7_69, w_ir_7_70, w_ir_7_71, w_ir_7_72, w_ir_7_73, w_ir_7_74, w_ir_7_75, w_ir_7_76, w_ir_7_77, w_ir_7_78, w_ir_7_79, w_ir_7_80, w_ir_7_81, w_ir_7_82, w_ir_7_83, w_ir_7_84, w_ir_7_85, w_ir_7_86, w_ir_7_87, w_ir_7_88, w_ir_7_89, w_ir_7_90, w_ir_7_91, w_ir_7_92, w_ir_7_93, w_ir_7_94, w_ir_7_95, w_ir_7_96, w_ir_7_97, w_ir_7_98, w_ir_7_99, w_ir_7_100, w_ir_7_101, w_ir_7_102, w_ir_7_103, w_ir_7_104, w_ir_7_105, w_ir_7_106, w_ir_7_107, w_ir_7_108, w_ir_7_109, w_ir_7_110, w_ir_7_111, w_ir_7_112, w_ir_7_113, w_ir_7_114, w_ir_7_115, w_ir_7_116, w_ir_7_117, w_ir_7_118, w_ir_7_119, w_ir_7_120, w_ir_7_121, w_ir_7_122, w_ir_7_123, w_ir_7_124, w_ir_7_125, w_ir_7_126, w_ir_7_127, w_ir_7_128, w_ir_7_129, w_ir_7_130, w_ir_7_131, w_ir_7_132, w_ir_7_133, w_ir_7_134, w_ir_7_135, w_ir_7_136, w_ir_7_137, w_ir_7_138, w_ir_7_139, w_ir_7_140, w_ir_7_141, w_ir_7_142, w_ir_7_143, w_ir_7_144, w_ir_7_145, w_ir_7_146, w_ir_7_147, w_ir_7_148, w_ir_7_149, w_ir_7_150, w_ir_7_151, w_ir_7_152, w_ir_7_153, w_ir_7_154, w_ir_7_155, w_ir_7_156, w_ir_7_157, w_ir_7_158, w_ir_7_159, w_ir_7_160, w_ir_7_161, w_ir_7_162, w_ir_7_163, w_ir_7_164, w_ir_7_165, w_ir_7_166, w_ir_7_167, w_ir_7_168, w_ir_7_169, w_ir_7_170, w_ir_7_171, w_ir_7_172, w_ir_7_173, w_ir_7_174, w_ir_7_175, w_ir_7_176, w_ir_7_177, w_ir_7_178, w_ir_7_179, w_ir_7_180, w_ir_7_181, w_ir_7_182, w_ir_7_183, w_ir_7_184, w_ir_7_185, w_ir_7_186, w_ir_7_187, w_ir_7_188, w_ir_7_189, w_ir_7_190, w_ir_7_191, w_ir_7_192, w_ir_7_193, w_ir_7_194, w_ir_7_195, w_ir_7_196, w_ir_7_197, w_ir_7_198, w_ir_7_199, w_ir_7_200, w_ir_7_201, w_ir_7_202, w_ir_7_203, w_ir_7_204, w_ir_7_205, w_ir_7_206, w_ir_7_207, w_ir_7_208, w_ir_7_209, w_ir_7_210, w_ir_7_211, w_ir_7_212, w_ir_7_213, w_ir_7_214, w_ir_7_215, w_ir_7_216, w_ir_7_217, w_ir_7_218, w_ir_7_219, w_ir_7_220, w_ir_7_221, w_ir_7_222, w_ir_7_223, w_ir_7_224, w_ir_7_225, w_ir_7_226, w_ir_7_227, w_ir_7_228, w_ir_7_229, w_ir_7_230, w_ir_7_231, w_ir_7_232, w_ir_7_233, w_ir_7_234, w_ir_7_235, w_ir_7_236, w_ir_7_237, w_ir_7_238, w_ir_7_239, w_ir_7_240, w_ir_7_241, w_ir_7_242, w_ir_7_243, w_ir_7_244, w_ir_7_245, w_ir_7_246, w_ir_7_247, w_ir_7_248, w_ir_7_249, w_ir_7_250, w_ir_7_251, w_ir_7_252, w_ir_7_253, w_ir_7_254, w_ir_7_255,
    input  logic signed [WIDTH-1:0]  w_iz_0_0, w_iz_0_1, w_iz_0_2, w_iz_0_3, w_iz_0_4, w_iz_0_5, w_iz_0_6, w_iz_0_7, w_iz_0_8, w_iz_0_9, w_iz_0_10, w_iz_0_11, w_iz_0_12, w_iz_0_13, w_iz_0_14, w_iz_0_15, w_iz_0_16, w_iz_0_17, w_iz_0_18, w_iz_0_19, w_iz_0_20, w_iz_0_21, w_iz_0_22, w_iz_0_23, w_iz_0_24, w_iz_0_25, w_iz_0_26, w_iz_0_27, w_iz_0_28, w_iz_0_29, w_iz_0_30, w_iz_0_31, w_iz_0_32, w_iz_0_33, w_iz_0_34, w_iz_0_35, w_iz_0_36, w_iz_0_37, w_iz_0_38, w_iz_0_39, w_iz_0_40, w_iz_0_41, w_iz_0_42, w_iz_0_43, w_iz_0_44, w_iz_0_45, w_iz_0_46, w_iz_0_47, w_iz_0_48, w_iz_0_49, w_iz_0_50, w_iz_0_51, w_iz_0_52, w_iz_0_53, w_iz_0_54, w_iz_0_55, w_iz_0_56, w_iz_0_57, w_iz_0_58, w_iz_0_59, w_iz_0_60, w_iz_0_61, w_iz_0_62, w_iz_0_63, w_iz_0_64, w_iz_0_65, w_iz_0_66, w_iz_0_67, w_iz_0_68, w_iz_0_69, w_iz_0_70, w_iz_0_71, w_iz_0_72, w_iz_0_73, w_iz_0_74, w_iz_0_75, w_iz_0_76, w_iz_0_77, w_iz_0_78, w_iz_0_79, w_iz_0_80, w_iz_0_81, w_iz_0_82, w_iz_0_83, w_iz_0_84, w_iz_0_85, w_iz_0_86, w_iz_0_87, w_iz_0_88, w_iz_0_89, w_iz_0_90, w_iz_0_91, w_iz_0_92, w_iz_0_93, w_iz_0_94, w_iz_0_95, w_iz_0_96, w_iz_0_97, w_iz_0_98, w_iz_0_99, w_iz_0_100, w_iz_0_101, w_iz_0_102, w_iz_0_103, w_iz_0_104, w_iz_0_105, w_iz_0_106, w_iz_0_107, w_iz_0_108, w_iz_0_109, w_iz_0_110, w_iz_0_111, w_iz_0_112, w_iz_0_113, w_iz_0_114, w_iz_0_115, w_iz_0_116, w_iz_0_117, w_iz_0_118, w_iz_0_119, w_iz_0_120, w_iz_0_121, w_iz_0_122, w_iz_0_123, w_iz_0_124, w_iz_0_125, w_iz_0_126, w_iz_0_127, w_iz_0_128, w_iz_0_129, w_iz_0_130, w_iz_0_131, w_iz_0_132, w_iz_0_133, w_iz_0_134, w_iz_0_135, w_iz_0_136, w_iz_0_137, w_iz_0_138, w_iz_0_139, w_iz_0_140, w_iz_0_141, w_iz_0_142, w_iz_0_143, w_iz_0_144, w_iz_0_145, w_iz_0_146, w_iz_0_147, w_iz_0_148, w_iz_0_149, w_iz_0_150, w_iz_0_151, w_iz_0_152, w_iz_0_153, w_iz_0_154, w_iz_0_155, w_iz_0_156, w_iz_0_157, w_iz_0_158, w_iz_0_159, w_iz_0_160, w_iz_0_161, w_iz_0_162, w_iz_0_163, w_iz_0_164, w_iz_0_165, w_iz_0_166, w_iz_0_167, w_iz_0_168, w_iz_0_169, w_iz_0_170, w_iz_0_171, w_iz_0_172, w_iz_0_173, w_iz_0_174, w_iz_0_175, w_iz_0_176, w_iz_0_177, w_iz_0_178, w_iz_0_179, w_iz_0_180, w_iz_0_181, w_iz_0_182, w_iz_0_183, w_iz_0_184, w_iz_0_185, w_iz_0_186, w_iz_0_187, w_iz_0_188, w_iz_0_189, w_iz_0_190, w_iz_0_191, w_iz_0_192, w_iz_0_193, w_iz_0_194, w_iz_0_195, w_iz_0_196, w_iz_0_197, w_iz_0_198, w_iz_0_199, w_iz_0_200, w_iz_0_201, w_iz_0_202, w_iz_0_203, w_iz_0_204, w_iz_0_205, w_iz_0_206, w_iz_0_207, w_iz_0_208, w_iz_0_209, w_iz_0_210, w_iz_0_211, w_iz_0_212, w_iz_0_213, w_iz_0_214, w_iz_0_215, w_iz_0_216, w_iz_0_217, w_iz_0_218, w_iz_0_219, w_iz_0_220, w_iz_0_221, w_iz_0_222, w_iz_0_223, w_iz_0_224, w_iz_0_225, w_iz_0_226, w_iz_0_227, w_iz_0_228, w_iz_0_229, w_iz_0_230, w_iz_0_231, w_iz_0_232, w_iz_0_233, w_iz_0_234, w_iz_0_235, w_iz_0_236, w_iz_0_237, w_iz_0_238, w_iz_0_239, w_iz_0_240, w_iz_0_241, w_iz_0_242, w_iz_0_243, w_iz_0_244, w_iz_0_245, w_iz_0_246, w_iz_0_247, w_iz_0_248, w_iz_0_249, w_iz_0_250, w_iz_0_251, w_iz_0_252, w_iz_0_253, w_iz_0_254, w_iz_0_255, w_iz_1_0, w_iz_1_1, w_iz_1_2, w_iz_1_3, w_iz_1_4, w_iz_1_5, w_iz_1_6, w_iz_1_7, w_iz_1_8, w_iz_1_9, w_iz_1_10, w_iz_1_11, w_iz_1_12, w_iz_1_13, w_iz_1_14, w_iz_1_15, w_iz_1_16, w_iz_1_17, w_iz_1_18, w_iz_1_19, w_iz_1_20, w_iz_1_21, w_iz_1_22, w_iz_1_23, w_iz_1_24, w_iz_1_25, w_iz_1_26, w_iz_1_27, w_iz_1_28, w_iz_1_29, w_iz_1_30, w_iz_1_31, w_iz_1_32, w_iz_1_33, w_iz_1_34, w_iz_1_35, w_iz_1_36, w_iz_1_37, w_iz_1_38, w_iz_1_39, w_iz_1_40, w_iz_1_41, w_iz_1_42, w_iz_1_43, w_iz_1_44, w_iz_1_45, w_iz_1_46, w_iz_1_47, w_iz_1_48, w_iz_1_49, w_iz_1_50, w_iz_1_51, w_iz_1_52, w_iz_1_53, w_iz_1_54, w_iz_1_55, w_iz_1_56, w_iz_1_57, w_iz_1_58, w_iz_1_59, w_iz_1_60, w_iz_1_61, w_iz_1_62, w_iz_1_63, w_iz_1_64, w_iz_1_65, w_iz_1_66, w_iz_1_67, w_iz_1_68, w_iz_1_69, w_iz_1_70, w_iz_1_71, w_iz_1_72, w_iz_1_73, w_iz_1_74, w_iz_1_75, w_iz_1_76, w_iz_1_77, w_iz_1_78, w_iz_1_79, w_iz_1_80, w_iz_1_81, w_iz_1_82, w_iz_1_83, w_iz_1_84, w_iz_1_85, w_iz_1_86, w_iz_1_87, w_iz_1_88, w_iz_1_89, w_iz_1_90, w_iz_1_91, w_iz_1_92, w_iz_1_93, w_iz_1_94, w_iz_1_95, w_iz_1_96, w_iz_1_97, w_iz_1_98, w_iz_1_99, w_iz_1_100, w_iz_1_101, w_iz_1_102, w_iz_1_103, w_iz_1_104, w_iz_1_105, w_iz_1_106, w_iz_1_107, w_iz_1_108, w_iz_1_109, w_iz_1_110, w_iz_1_111, w_iz_1_112, w_iz_1_113, w_iz_1_114, w_iz_1_115, w_iz_1_116, w_iz_1_117, w_iz_1_118, w_iz_1_119, w_iz_1_120, w_iz_1_121, w_iz_1_122, w_iz_1_123, w_iz_1_124, w_iz_1_125, w_iz_1_126, w_iz_1_127, w_iz_1_128, w_iz_1_129, w_iz_1_130, w_iz_1_131, w_iz_1_132, w_iz_1_133, w_iz_1_134, w_iz_1_135, w_iz_1_136, w_iz_1_137, w_iz_1_138, w_iz_1_139, w_iz_1_140, w_iz_1_141, w_iz_1_142, w_iz_1_143, w_iz_1_144, w_iz_1_145, w_iz_1_146, w_iz_1_147, w_iz_1_148, w_iz_1_149, w_iz_1_150, w_iz_1_151, w_iz_1_152, w_iz_1_153, w_iz_1_154, w_iz_1_155, w_iz_1_156, w_iz_1_157, w_iz_1_158, w_iz_1_159, w_iz_1_160, w_iz_1_161, w_iz_1_162, w_iz_1_163, w_iz_1_164, w_iz_1_165, w_iz_1_166, w_iz_1_167, w_iz_1_168, w_iz_1_169, w_iz_1_170, w_iz_1_171, w_iz_1_172, w_iz_1_173, w_iz_1_174, w_iz_1_175, w_iz_1_176, w_iz_1_177, w_iz_1_178, w_iz_1_179, w_iz_1_180, w_iz_1_181, w_iz_1_182, w_iz_1_183, w_iz_1_184, w_iz_1_185, w_iz_1_186, w_iz_1_187, w_iz_1_188, w_iz_1_189, w_iz_1_190, w_iz_1_191, w_iz_1_192, w_iz_1_193, w_iz_1_194, w_iz_1_195, w_iz_1_196, w_iz_1_197, w_iz_1_198, w_iz_1_199, w_iz_1_200, w_iz_1_201, w_iz_1_202, w_iz_1_203, w_iz_1_204, w_iz_1_205, w_iz_1_206, w_iz_1_207, w_iz_1_208, w_iz_1_209, w_iz_1_210, w_iz_1_211, w_iz_1_212, w_iz_1_213, w_iz_1_214, w_iz_1_215, w_iz_1_216, w_iz_1_217, w_iz_1_218, w_iz_1_219, w_iz_1_220, w_iz_1_221, w_iz_1_222, w_iz_1_223, w_iz_1_224, w_iz_1_225, w_iz_1_226, w_iz_1_227, w_iz_1_228, w_iz_1_229, w_iz_1_230, w_iz_1_231, w_iz_1_232, w_iz_1_233, w_iz_1_234, w_iz_1_235, w_iz_1_236, w_iz_1_237, w_iz_1_238, w_iz_1_239, w_iz_1_240, w_iz_1_241, w_iz_1_242, w_iz_1_243, w_iz_1_244, w_iz_1_245, w_iz_1_246, w_iz_1_247, w_iz_1_248, w_iz_1_249, w_iz_1_250, w_iz_1_251, w_iz_1_252, w_iz_1_253, w_iz_1_254, w_iz_1_255, w_iz_2_0, w_iz_2_1, w_iz_2_2, w_iz_2_3, w_iz_2_4, w_iz_2_5, w_iz_2_6, w_iz_2_7, w_iz_2_8, w_iz_2_9, w_iz_2_10, w_iz_2_11, w_iz_2_12, w_iz_2_13, w_iz_2_14, w_iz_2_15, w_iz_2_16, w_iz_2_17, w_iz_2_18, w_iz_2_19, w_iz_2_20, w_iz_2_21, w_iz_2_22, w_iz_2_23, w_iz_2_24, w_iz_2_25, w_iz_2_26, w_iz_2_27, w_iz_2_28, w_iz_2_29, w_iz_2_30, w_iz_2_31, w_iz_2_32, w_iz_2_33, w_iz_2_34, w_iz_2_35, w_iz_2_36, w_iz_2_37, w_iz_2_38, w_iz_2_39, w_iz_2_40, w_iz_2_41, w_iz_2_42, w_iz_2_43, w_iz_2_44, w_iz_2_45, w_iz_2_46, w_iz_2_47, w_iz_2_48, w_iz_2_49, w_iz_2_50, w_iz_2_51, w_iz_2_52, w_iz_2_53, w_iz_2_54, w_iz_2_55, w_iz_2_56, w_iz_2_57, w_iz_2_58, w_iz_2_59, w_iz_2_60, w_iz_2_61, w_iz_2_62, w_iz_2_63, w_iz_2_64, w_iz_2_65, w_iz_2_66, w_iz_2_67, w_iz_2_68, w_iz_2_69, w_iz_2_70, w_iz_2_71, w_iz_2_72, w_iz_2_73, w_iz_2_74, w_iz_2_75, w_iz_2_76, w_iz_2_77, w_iz_2_78, w_iz_2_79, w_iz_2_80, w_iz_2_81, w_iz_2_82, w_iz_2_83, w_iz_2_84, w_iz_2_85, w_iz_2_86, w_iz_2_87, w_iz_2_88, w_iz_2_89, w_iz_2_90, w_iz_2_91, w_iz_2_92, w_iz_2_93, w_iz_2_94, w_iz_2_95, w_iz_2_96, w_iz_2_97, w_iz_2_98, w_iz_2_99, w_iz_2_100, w_iz_2_101, w_iz_2_102, w_iz_2_103, w_iz_2_104, w_iz_2_105, w_iz_2_106, w_iz_2_107, w_iz_2_108, w_iz_2_109, w_iz_2_110, w_iz_2_111, w_iz_2_112, w_iz_2_113, w_iz_2_114, w_iz_2_115, w_iz_2_116, w_iz_2_117, w_iz_2_118, w_iz_2_119, w_iz_2_120, w_iz_2_121, w_iz_2_122, w_iz_2_123, w_iz_2_124, w_iz_2_125, w_iz_2_126, w_iz_2_127, w_iz_2_128, w_iz_2_129, w_iz_2_130, w_iz_2_131, w_iz_2_132, w_iz_2_133, w_iz_2_134, w_iz_2_135, w_iz_2_136, w_iz_2_137, w_iz_2_138, w_iz_2_139, w_iz_2_140, w_iz_2_141, w_iz_2_142, w_iz_2_143, w_iz_2_144, w_iz_2_145, w_iz_2_146, w_iz_2_147, w_iz_2_148, w_iz_2_149, w_iz_2_150, w_iz_2_151, w_iz_2_152, w_iz_2_153, w_iz_2_154, w_iz_2_155, w_iz_2_156, w_iz_2_157, w_iz_2_158, w_iz_2_159, w_iz_2_160, w_iz_2_161, w_iz_2_162, w_iz_2_163, w_iz_2_164, w_iz_2_165, w_iz_2_166, w_iz_2_167, w_iz_2_168, w_iz_2_169, w_iz_2_170, w_iz_2_171, w_iz_2_172, w_iz_2_173, w_iz_2_174, w_iz_2_175, w_iz_2_176, w_iz_2_177, w_iz_2_178, w_iz_2_179, w_iz_2_180, w_iz_2_181, w_iz_2_182, w_iz_2_183, w_iz_2_184, w_iz_2_185, w_iz_2_186, w_iz_2_187, w_iz_2_188, w_iz_2_189, w_iz_2_190, w_iz_2_191, w_iz_2_192, w_iz_2_193, w_iz_2_194, w_iz_2_195, w_iz_2_196, w_iz_2_197, w_iz_2_198, w_iz_2_199, w_iz_2_200, w_iz_2_201, w_iz_2_202, w_iz_2_203, w_iz_2_204, w_iz_2_205, w_iz_2_206, w_iz_2_207, w_iz_2_208, w_iz_2_209, w_iz_2_210, w_iz_2_211, w_iz_2_212, w_iz_2_213, w_iz_2_214, w_iz_2_215, w_iz_2_216, w_iz_2_217, w_iz_2_218, w_iz_2_219, w_iz_2_220, w_iz_2_221, w_iz_2_222, w_iz_2_223, w_iz_2_224, w_iz_2_225, w_iz_2_226, w_iz_2_227, w_iz_2_228, w_iz_2_229, w_iz_2_230, w_iz_2_231, w_iz_2_232, w_iz_2_233, w_iz_2_234, w_iz_2_235, w_iz_2_236, w_iz_2_237, w_iz_2_238, w_iz_2_239, w_iz_2_240, w_iz_2_241, w_iz_2_242, w_iz_2_243, w_iz_2_244, w_iz_2_245, w_iz_2_246, w_iz_2_247, w_iz_2_248, w_iz_2_249, w_iz_2_250, w_iz_2_251, w_iz_2_252, w_iz_2_253, w_iz_2_254, w_iz_2_255, w_iz_3_0, w_iz_3_1, w_iz_3_2, w_iz_3_3, w_iz_3_4, w_iz_3_5, w_iz_3_6, w_iz_3_7, w_iz_3_8, w_iz_3_9, w_iz_3_10, w_iz_3_11, w_iz_3_12, w_iz_3_13, w_iz_3_14, w_iz_3_15, w_iz_3_16, w_iz_3_17, w_iz_3_18, w_iz_3_19, w_iz_3_20, w_iz_3_21, w_iz_3_22, w_iz_3_23, w_iz_3_24, w_iz_3_25, w_iz_3_26, w_iz_3_27, w_iz_3_28, w_iz_3_29, w_iz_3_30, w_iz_3_31, w_iz_3_32, w_iz_3_33, w_iz_3_34, w_iz_3_35, w_iz_3_36, w_iz_3_37, w_iz_3_38, w_iz_3_39, w_iz_3_40, w_iz_3_41, w_iz_3_42, w_iz_3_43, w_iz_3_44, w_iz_3_45, w_iz_3_46, w_iz_3_47, w_iz_3_48, w_iz_3_49, w_iz_3_50, w_iz_3_51, w_iz_3_52, w_iz_3_53, w_iz_3_54, w_iz_3_55, w_iz_3_56, w_iz_3_57, w_iz_3_58, w_iz_3_59, w_iz_3_60, w_iz_3_61, w_iz_3_62, w_iz_3_63, w_iz_3_64, w_iz_3_65, w_iz_3_66, w_iz_3_67, w_iz_3_68, w_iz_3_69, w_iz_3_70, w_iz_3_71, w_iz_3_72, w_iz_3_73, w_iz_3_74, w_iz_3_75, w_iz_3_76, w_iz_3_77, w_iz_3_78, w_iz_3_79, w_iz_3_80, w_iz_3_81, w_iz_3_82, w_iz_3_83, w_iz_3_84, w_iz_3_85, w_iz_3_86, w_iz_3_87, w_iz_3_88, w_iz_3_89, w_iz_3_90, w_iz_3_91, w_iz_3_92, w_iz_3_93, w_iz_3_94, w_iz_3_95, w_iz_3_96, w_iz_3_97, w_iz_3_98, w_iz_3_99, w_iz_3_100, w_iz_3_101, w_iz_3_102, w_iz_3_103, w_iz_3_104, w_iz_3_105, w_iz_3_106, w_iz_3_107, w_iz_3_108, w_iz_3_109, w_iz_3_110, w_iz_3_111, w_iz_3_112, w_iz_3_113, w_iz_3_114, w_iz_3_115, w_iz_3_116, w_iz_3_117, w_iz_3_118, w_iz_3_119, w_iz_3_120, w_iz_3_121, w_iz_3_122, w_iz_3_123, w_iz_3_124, w_iz_3_125, w_iz_3_126, w_iz_3_127, w_iz_3_128, w_iz_3_129, w_iz_3_130, w_iz_3_131, w_iz_3_132, w_iz_3_133, w_iz_3_134, w_iz_3_135, w_iz_3_136, w_iz_3_137, w_iz_3_138, w_iz_3_139, w_iz_3_140, w_iz_3_141, w_iz_3_142, w_iz_3_143, w_iz_3_144, w_iz_3_145, w_iz_3_146, w_iz_3_147, w_iz_3_148, w_iz_3_149, w_iz_3_150, w_iz_3_151, w_iz_3_152, w_iz_3_153, w_iz_3_154, w_iz_3_155, w_iz_3_156, w_iz_3_157, w_iz_3_158, w_iz_3_159, w_iz_3_160, w_iz_3_161, w_iz_3_162, w_iz_3_163, w_iz_3_164, w_iz_3_165, w_iz_3_166, w_iz_3_167, w_iz_3_168, w_iz_3_169, w_iz_3_170, w_iz_3_171, w_iz_3_172, w_iz_3_173, w_iz_3_174, w_iz_3_175, w_iz_3_176, w_iz_3_177, w_iz_3_178, w_iz_3_179, w_iz_3_180, w_iz_3_181, w_iz_3_182, w_iz_3_183, w_iz_3_184, w_iz_3_185, w_iz_3_186, w_iz_3_187, w_iz_3_188, w_iz_3_189, w_iz_3_190, w_iz_3_191, w_iz_3_192, w_iz_3_193, w_iz_3_194, w_iz_3_195, w_iz_3_196, w_iz_3_197, w_iz_3_198, w_iz_3_199, w_iz_3_200, w_iz_3_201, w_iz_3_202, w_iz_3_203, w_iz_3_204, w_iz_3_205, w_iz_3_206, w_iz_3_207, w_iz_3_208, w_iz_3_209, w_iz_3_210, w_iz_3_211, w_iz_3_212, w_iz_3_213, w_iz_3_214, w_iz_3_215, w_iz_3_216, w_iz_3_217, w_iz_3_218, w_iz_3_219, w_iz_3_220, w_iz_3_221, w_iz_3_222, w_iz_3_223, w_iz_3_224, w_iz_3_225, w_iz_3_226, w_iz_3_227, w_iz_3_228, w_iz_3_229, w_iz_3_230, w_iz_3_231, w_iz_3_232, w_iz_3_233, w_iz_3_234, w_iz_3_235, w_iz_3_236, w_iz_3_237, w_iz_3_238, w_iz_3_239, w_iz_3_240, w_iz_3_241, w_iz_3_242, w_iz_3_243, w_iz_3_244, w_iz_3_245, w_iz_3_246, w_iz_3_247, w_iz_3_248, w_iz_3_249, w_iz_3_250, w_iz_3_251, w_iz_3_252, w_iz_3_253, w_iz_3_254, w_iz_3_255, w_iz_4_0, w_iz_4_1, w_iz_4_2, w_iz_4_3, w_iz_4_4, w_iz_4_5, w_iz_4_6, w_iz_4_7, w_iz_4_8, w_iz_4_9, w_iz_4_10, w_iz_4_11, w_iz_4_12, w_iz_4_13, w_iz_4_14, w_iz_4_15, w_iz_4_16, w_iz_4_17, w_iz_4_18, w_iz_4_19, w_iz_4_20, w_iz_4_21, w_iz_4_22, w_iz_4_23, w_iz_4_24, w_iz_4_25, w_iz_4_26, w_iz_4_27, w_iz_4_28, w_iz_4_29, w_iz_4_30, w_iz_4_31, w_iz_4_32, w_iz_4_33, w_iz_4_34, w_iz_4_35, w_iz_4_36, w_iz_4_37, w_iz_4_38, w_iz_4_39, w_iz_4_40, w_iz_4_41, w_iz_4_42, w_iz_4_43, w_iz_4_44, w_iz_4_45, w_iz_4_46, w_iz_4_47, w_iz_4_48, w_iz_4_49, w_iz_4_50, w_iz_4_51, w_iz_4_52, w_iz_4_53, w_iz_4_54, w_iz_4_55, w_iz_4_56, w_iz_4_57, w_iz_4_58, w_iz_4_59, w_iz_4_60, w_iz_4_61, w_iz_4_62, w_iz_4_63, w_iz_4_64, w_iz_4_65, w_iz_4_66, w_iz_4_67, w_iz_4_68, w_iz_4_69, w_iz_4_70, w_iz_4_71, w_iz_4_72, w_iz_4_73, w_iz_4_74, w_iz_4_75, w_iz_4_76, w_iz_4_77, w_iz_4_78, w_iz_4_79, w_iz_4_80, w_iz_4_81, w_iz_4_82, w_iz_4_83, w_iz_4_84, w_iz_4_85, w_iz_4_86, w_iz_4_87, w_iz_4_88, w_iz_4_89, w_iz_4_90, w_iz_4_91, w_iz_4_92, w_iz_4_93, w_iz_4_94, w_iz_4_95, w_iz_4_96, w_iz_4_97, w_iz_4_98, w_iz_4_99, w_iz_4_100, w_iz_4_101, w_iz_4_102, w_iz_4_103, w_iz_4_104, w_iz_4_105, w_iz_4_106, w_iz_4_107, w_iz_4_108, w_iz_4_109, w_iz_4_110, w_iz_4_111, w_iz_4_112, w_iz_4_113, w_iz_4_114, w_iz_4_115, w_iz_4_116, w_iz_4_117, w_iz_4_118, w_iz_4_119, w_iz_4_120, w_iz_4_121, w_iz_4_122, w_iz_4_123, w_iz_4_124, w_iz_4_125, w_iz_4_126, w_iz_4_127, w_iz_4_128, w_iz_4_129, w_iz_4_130, w_iz_4_131, w_iz_4_132, w_iz_4_133, w_iz_4_134, w_iz_4_135, w_iz_4_136, w_iz_4_137, w_iz_4_138, w_iz_4_139, w_iz_4_140, w_iz_4_141, w_iz_4_142, w_iz_4_143, w_iz_4_144, w_iz_4_145, w_iz_4_146, w_iz_4_147, w_iz_4_148, w_iz_4_149, w_iz_4_150, w_iz_4_151, w_iz_4_152, w_iz_4_153, w_iz_4_154, w_iz_4_155, w_iz_4_156, w_iz_4_157, w_iz_4_158, w_iz_4_159, w_iz_4_160, w_iz_4_161, w_iz_4_162, w_iz_4_163, w_iz_4_164, w_iz_4_165, w_iz_4_166, w_iz_4_167, w_iz_4_168, w_iz_4_169, w_iz_4_170, w_iz_4_171, w_iz_4_172, w_iz_4_173, w_iz_4_174, w_iz_4_175, w_iz_4_176, w_iz_4_177, w_iz_4_178, w_iz_4_179, w_iz_4_180, w_iz_4_181, w_iz_4_182, w_iz_4_183, w_iz_4_184, w_iz_4_185, w_iz_4_186, w_iz_4_187, w_iz_4_188, w_iz_4_189, w_iz_4_190, w_iz_4_191, w_iz_4_192, w_iz_4_193, w_iz_4_194, w_iz_4_195, w_iz_4_196, w_iz_4_197, w_iz_4_198, w_iz_4_199, w_iz_4_200, w_iz_4_201, w_iz_4_202, w_iz_4_203, w_iz_4_204, w_iz_4_205, w_iz_4_206, w_iz_4_207, w_iz_4_208, w_iz_4_209, w_iz_4_210, w_iz_4_211, w_iz_4_212, w_iz_4_213, w_iz_4_214, w_iz_4_215, w_iz_4_216, w_iz_4_217, w_iz_4_218, w_iz_4_219, w_iz_4_220, w_iz_4_221, w_iz_4_222, w_iz_4_223, w_iz_4_224, w_iz_4_225, w_iz_4_226, w_iz_4_227, w_iz_4_228, w_iz_4_229, w_iz_4_230, w_iz_4_231, w_iz_4_232, w_iz_4_233, w_iz_4_234, w_iz_4_235, w_iz_4_236, w_iz_4_237, w_iz_4_238, w_iz_4_239, w_iz_4_240, w_iz_4_241, w_iz_4_242, w_iz_4_243, w_iz_4_244, w_iz_4_245, w_iz_4_246, w_iz_4_247, w_iz_4_248, w_iz_4_249, w_iz_4_250, w_iz_4_251, w_iz_4_252, w_iz_4_253, w_iz_4_254, w_iz_4_255, w_iz_5_0, w_iz_5_1, w_iz_5_2, w_iz_5_3, w_iz_5_4, w_iz_5_5, w_iz_5_6, w_iz_5_7, w_iz_5_8, w_iz_5_9, w_iz_5_10, w_iz_5_11, w_iz_5_12, w_iz_5_13, w_iz_5_14, w_iz_5_15, w_iz_5_16, w_iz_5_17, w_iz_5_18, w_iz_5_19, w_iz_5_20, w_iz_5_21, w_iz_5_22, w_iz_5_23, w_iz_5_24, w_iz_5_25, w_iz_5_26, w_iz_5_27, w_iz_5_28, w_iz_5_29, w_iz_5_30, w_iz_5_31, w_iz_5_32, w_iz_5_33, w_iz_5_34, w_iz_5_35, w_iz_5_36, w_iz_5_37, w_iz_5_38, w_iz_5_39, w_iz_5_40, w_iz_5_41, w_iz_5_42, w_iz_5_43, w_iz_5_44, w_iz_5_45, w_iz_5_46, w_iz_5_47, w_iz_5_48, w_iz_5_49, w_iz_5_50, w_iz_5_51, w_iz_5_52, w_iz_5_53, w_iz_5_54, w_iz_5_55, w_iz_5_56, w_iz_5_57, w_iz_5_58, w_iz_5_59, w_iz_5_60, w_iz_5_61, w_iz_5_62, w_iz_5_63, w_iz_5_64, w_iz_5_65, w_iz_5_66, w_iz_5_67, w_iz_5_68, w_iz_5_69, w_iz_5_70, w_iz_5_71, w_iz_5_72, w_iz_5_73, w_iz_5_74, w_iz_5_75, w_iz_5_76, w_iz_5_77, w_iz_5_78, w_iz_5_79, w_iz_5_80, w_iz_5_81, w_iz_5_82, w_iz_5_83, w_iz_5_84, w_iz_5_85, w_iz_5_86, w_iz_5_87, w_iz_5_88, w_iz_5_89, w_iz_5_90, w_iz_5_91, w_iz_5_92, w_iz_5_93, w_iz_5_94, w_iz_5_95, w_iz_5_96, w_iz_5_97, w_iz_5_98, w_iz_5_99, w_iz_5_100, w_iz_5_101, w_iz_5_102, w_iz_5_103, w_iz_5_104, w_iz_5_105, w_iz_5_106, w_iz_5_107, w_iz_5_108, w_iz_5_109, w_iz_5_110, w_iz_5_111, w_iz_5_112, w_iz_5_113, w_iz_5_114, w_iz_5_115, w_iz_5_116, w_iz_5_117, w_iz_5_118, w_iz_5_119, w_iz_5_120, w_iz_5_121, w_iz_5_122, w_iz_5_123, w_iz_5_124, w_iz_5_125, w_iz_5_126, w_iz_5_127, w_iz_5_128, w_iz_5_129, w_iz_5_130, w_iz_5_131, w_iz_5_132, w_iz_5_133, w_iz_5_134, w_iz_5_135, w_iz_5_136, w_iz_5_137, w_iz_5_138, w_iz_5_139, w_iz_5_140, w_iz_5_141, w_iz_5_142, w_iz_5_143, w_iz_5_144, w_iz_5_145, w_iz_5_146, w_iz_5_147, w_iz_5_148, w_iz_5_149, w_iz_5_150, w_iz_5_151, w_iz_5_152, w_iz_5_153, w_iz_5_154, w_iz_5_155, w_iz_5_156, w_iz_5_157, w_iz_5_158, w_iz_5_159, w_iz_5_160, w_iz_5_161, w_iz_5_162, w_iz_5_163, w_iz_5_164, w_iz_5_165, w_iz_5_166, w_iz_5_167, w_iz_5_168, w_iz_5_169, w_iz_5_170, w_iz_5_171, w_iz_5_172, w_iz_5_173, w_iz_5_174, w_iz_5_175, w_iz_5_176, w_iz_5_177, w_iz_5_178, w_iz_5_179, w_iz_5_180, w_iz_5_181, w_iz_5_182, w_iz_5_183, w_iz_5_184, w_iz_5_185, w_iz_5_186, w_iz_5_187, w_iz_5_188, w_iz_5_189, w_iz_5_190, w_iz_5_191, w_iz_5_192, w_iz_5_193, w_iz_5_194, w_iz_5_195, w_iz_5_196, w_iz_5_197, w_iz_5_198, w_iz_5_199, w_iz_5_200, w_iz_5_201, w_iz_5_202, w_iz_5_203, w_iz_5_204, w_iz_5_205, w_iz_5_206, w_iz_5_207, w_iz_5_208, w_iz_5_209, w_iz_5_210, w_iz_5_211, w_iz_5_212, w_iz_5_213, w_iz_5_214, w_iz_5_215, w_iz_5_216, w_iz_5_217, w_iz_5_218, w_iz_5_219, w_iz_5_220, w_iz_5_221, w_iz_5_222, w_iz_5_223, w_iz_5_224, w_iz_5_225, w_iz_5_226, w_iz_5_227, w_iz_5_228, w_iz_5_229, w_iz_5_230, w_iz_5_231, w_iz_5_232, w_iz_5_233, w_iz_5_234, w_iz_5_235, w_iz_5_236, w_iz_5_237, w_iz_5_238, w_iz_5_239, w_iz_5_240, w_iz_5_241, w_iz_5_242, w_iz_5_243, w_iz_5_244, w_iz_5_245, w_iz_5_246, w_iz_5_247, w_iz_5_248, w_iz_5_249, w_iz_5_250, w_iz_5_251, w_iz_5_252, w_iz_5_253, w_iz_5_254, w_iz_5_255, w_iz_6_0, w_iz_6_1, w_iz_6_2, w_iz_6_3, w_iz_6_4, w_iz_6_5, w_iz_6_6, w_iz_6_7, w_iz_6_8, w_iz_6_9, w_iz_6_10, w_iz_6_11, w_iz_6_12, w_iz_6_13, w_iz_6_14, w_iz_6_15, w_iz_6_16, w_iz_6_17, w_iz_6_18, w_iz_6_19, w_iz_6_20, w_iz_6_21, w_iz_6_22, w_iz_6_23, w_iz_6_24, w_iz_6_25, w_iz_6_26, w_iz_6_27, w_iz_6_28, w_iz_6_29, w_iz_6_30, w_iz_6_31, w_iz_6_32, w_iz_6_33, w_iz_6_34, w_iz_6_35, w_iz_6_36, w_iz_6_37, w_iz_6_38, w_iz_6_39, w_iz_6_40, w_iz_6_41, w_iz_6_42, w_iz_6_43, w_iz_6_44, w_iz_6_45, w_iz_6_46, w_iz_6_47, w_iz_6_48, w_iz_6_49, w_iz_6_50, w_iz_6_51, w_iz_6_52, w_iz_6_53, w_iz_6_54, w_iz_6_55, w_iz_6_56, w_iz_6_57, w_iz_6_58, w_iz_6_59, w_iz_6_60, w_iz_6_61, w_iz_6_62, w_iz_6_63, w_iz_6_64, w_iz_6_65, w_iz_6_66, w_iz_6_67, w_iz_6_68, w_iz_6_69, w_iz_6_70, w_iz_6_71, w_iz_6_72, w_iz_6_73, w_iz_6_74, w_iz_6_75, w_iz_6_76, w_iz_6_77, w_iz_6_78, w_iz_6_79, w_iz_6_80, w_iz_6_81, w_iz_6_82, w_iz_6_83, w_iz_6_84, w_iz_6_85, w_iz_6_86, w_iz_6_87, w_iz_6_88, w_iz_6_89, w_iz_6_90, w_iz_6_91, w_iz_6_92, w_iz_6_93, w_iz_6_94, w_iz_6_95, w_iz_6_96, w_iz_6_97, w_iz_6_98, w_iz_6_99, w_iz_6_100, w_iz_6_101, w_iz_6_102, w_iz_6_103, w_iz_6_104, w_iz_6_105, w_iz_6_106, w_iz_6_107, w_iz_6_108, w_iz_6_109, w_iz_6_110, w_iz_6_111, w_iz_6_112, w_iz_6_113, w_iz_6_114, w_iz_6_115, w_iz_6_116, w_iz_6_117, w_iz_6_118, w_iz_6_119, w_iz_6_120, w_iz_6_121, w_iz_6_122, w_iz_6_123, w_iz_6_124, w_iz_6_125, w_iz_6_126, w_iz_6_127, w_iz_6_128, w_iz_6_129, w_iz_6_130, w_iz_6_131, w_iz_6_132, w_iz_6_133, w_iz_6_134, w_iz_6_135, w_iz_6_136, w_iz_6_137, w_iz_6_138, w_iz_6_139, w_iz_6_140, w_iz_6_141, w_iz_6_142, w_iz_6_143, w_iz_6_144, w_iz_6_145, w_iz_6_146, w_iz_6_147, w_iz_6_148, w_iz_6_149, w_iz_6_150, w_iz_6_151, w_iz_6_152, w_iz_6_153, w_iz_6_154, w_iz_6_155, w_iz_6_156, w_iz_6_157, w_iz_6_158, w_iz_6_159, w_iz_6_160, w_iz_6_161, w_iz_6_162, w_iz_6_163, w_iz_6_164, w_iz_6_165, w_iz_6_166, w_iz_6_167, w_iz_6_168, w_iz_6_169, w_iz_6_170, w_iz_6_171, w_iz_6_172, w_iz_6_173, w_iz_6_174, w_iz_6_175, w_iz_6_176, w_iz_6_177, w_iz_6_178, w_iz_6_179, w_iz_6_180, w_iz_6_181, w_iz_6_182, w_iz_6_183, w_iz_6_184, w_iz_6_185, w_iz_6_186, w_iz_6_187, w_iz_6_188, w_iz_6_189, w_iz_6_190, w_iz_6_191, w_iz_6_192, w_iz_6_193, w_iz_6_194, w_iz_6_195, w_iz_6_196, w_iz_6_197, w_iz_6_198, w_iz_6_199, w_iz_6_200, w_iz_6_201, w_iz_6_202, w_iz_6_203, w_iz_6_204, w_iz_6_205, w_iz_6_206, w_iz_6_207, w_iz_6_208, w_iz_6_209, w_iz_6_210, w_iz_6_211, w_iz_6_212, w_iz_6_213, w_iz_6_214, w_iz_6_215, w_iz_6_216, w_iz_6_217, w_iz_6_218, w_iz_6_219, w_iz_6_220, w_iz_6_221, w_iz_6_222, w_iz_6_223, w_iz_6_224, w_iz_6_225, w_iz_6_226, w_iz_6_227, w_iz_6_228, w_iz_6_229, w_iz_6_230, w_iz_6_231, w_iz_6_232, w_iz_6_233, w_iz_6_234, w_iz_6_235, w_iz_6_236, w_iz_6_237, w_iz_6_238, w_iz_6_239, w_iz_6_240, w_iz_6_241, w_iz_6_242, w_iz_6_243, w_iz_6_244, w_iz_6_245, w_iz_6_246, w_iz_6_247, w_iz_6_248, w_iz_6_249, w_iz_6_250, w_iz_6_251, w_iz_6_252, w_iz_6_253, w_iz_6_254, w_iz_6_255, w_iz_7_0, w_iz_7_1, w_iz_7_2, w_iz_7_3, w_iz_7_4, w_iz_7_5, w_iz_7_6, w_iz_7_7, w_iz_7_8, w_iz_7_9, w_iz_7_10, w_iz_7_11, w_iz_7_12, w_iz_7_13, w_iz_7_14, w_iz_7_15, w_iz_7_16, w_iz_7_17, w_iz_7_18, w_iz_7_19, w_iz_7_20, w_iz_7_21, w_iz_7_22, w_iz_7_23, w_iz_7_24, w_iz_7_25, w_iz_7_26, w_iz_7_27, w_iz_7_28, w_iz_7_29, w_iz_7_30, w_iz_7_31, w_iz_7_32, w_iz_7_33, w_iz_7_34, w_iz_7_35, w_iz_7_36, w_iz_7_37, w_iz_7_38, w_iz_7_39, w_iz_7_40, w_iz_7_41, w_iz_7_42, w_iz_7_43, w_iz_7_44, w_iz_7_45, w_iz_7_46, w_iz_7_47, w_iz_7_48, w_iz_7_49, w_iz_7_50, w_iz_7_51, w_iz_7_52, w_iz_7_53, w_iz_7_54, w_iz_7_55, w_iz_7_56, w_iz_7_57, w_iz_7_58, w_iz_7_59, w_iz_7_60, w_iz_7_61, w_iz_7_62, w_iz_7_63, w_iz_7_64, w_iz_7_65, w_iz_7_66, w_iz_7_67, w_iz_7_68, w_iz_7_69, w_iz_7_70, w_iz_7_71, w_iz_7_72, w_iz_7_73, w_iz_7_74, w_iz_7_75, w_iz_7_76, w_iz_7_77, w_iz_7_78, w_iz_7_79, w_iz_7_80, w_iz_7_81, w_iz_7_82, w_iz_7_83, w_iz_7_84, w_iz_7_85, w_iz_7_86, w_iz_7_87, w_iz_7_88, w_iz_7_89, w_iz_7_90, w_iz_7_91, w_iz_7_92, w_iz_7_93, w_iz_7_94, w_iz_7_95, w_iz_7_96, w_iz_7_97, w_iz_7_98, w_iz_7_99, w_iz_7_100, w_iz_7_101, w_iz_7_102, w_iz_7_103, w_iz_7_104, w_iz_7_105, w_iz_7_106, w_iz_7_107, w_iz_7_108, w_iz_7_109, w_iz_7_110, w_iz_7_111, w_iz_7_112, w_iz_7_113, w_iz_7_114, w_iz_7_115, w_iz_7_116, w_iz_7_117, w_iz_7_118, w_iz_7_119, w_iz_7_120, w_iz_7_121, w_iz_7_122, w_iz_7_123, w_iz_7_124, w_iz_7_125, w_iz_7_126, w_iz_7_127, w_iz_7_128, w_iz_7_129, w_iz_7_130, w_iz_7_131, w_iz_7_132, w_iz_7_133, w_iz_7_134, w_iz_7_135, w_iz_7_136, w_iz_7_137, w_iz_7_138, w_iz_7_139, w_iz_7_140, w_iz_7_141, w_iz_7_142, w_iz_7_143, w_iz_7_144, w_iz_7_145, w_iz_7_146, w_iz_7_147, w_iz_7_148, w_iz_7_149, w_iz_7_150, w_iz_7_151, w_iz_7_152, w_iz_7_153, w_iz_7_154, w_iz_7_155, w_iz_7_156, w_iz_7_157, w_iz_7_158, w_iz_7_159, w_iz_7_160, w_iz_7_161, w_iz_7_162, w_iz_7_163, w_iz_7_164, w_iz_7_165, w_iz_7_166, w_iz_7_167, w_iz_7_168, w_iz_7_169, w_iz_7_170, w_iz_7_171, w_iz_7_172, w_iz_7_173, w_iz_7_174, w_iz_7_175, w_iz_7_176, w_iz_7_177, w_iz_7_178, w_iz_7_179, w_iz_7_180, w_iz_7_181, w_iz_7_182, w_iz_7_183, w_iz_7_184, w_iz_7_185, w_iz_7_186, w_iz_7_187, w_iz_7_188, w_iz_7_189, w_iz_7_190, w_iz_7_191, w_iz_7_192, w_iz_7_193, w_iz_7_194, w_iz_7_195, w_iz_7_196, w_iz_7_197, w_iz_7_198, w_iz_7_199, w_iz_7_200, w_iz_7_201, w_iz_7_202, w_iz_7_203, w_iz_7_204, w_iz_7_205, w_iz_7_206, w_iz_7_207, w_iz_7_208, w_iz_7_209, w_iz_7_210, w_iz_7_211, w_iz_7_212, w_iz_7_213, w_iz_7_214, w_iz_7_215, w_iz_7_216, w_iz_7_217, w_iz_7_218, w_iz_7_219, w_iz_7_220, w_iz_7_221, w_iz_7_222, w_iz_7_223, w_iz_7_224, w_iz_7_225, w_iz_7_226, w_iz_7_227, w_iz_7_228, w_iz_7_229, w_iz_7_230, w_iz_7_231, w_iz_7_232, w_iz_7_233, w_iz_7_234, w_iz_7_235, w_iz_7_236, w_iz_7_237, w_iz_7_238, w_iz_7_239, w_iz_7_240, w_iz_7_241, w_iz_7_242, w_iz_7_243, w_iz_7_244, w_iz_7_245, w_iz_7_246, w_iz_7_247, w_iz_7_248, w_iz_7_249, w_iz_7_250, w_iz_7_251, w_iz_7_252, w_iz_7_253, w_iz_7_254, w_iz_7_255,
    input  logic signed [WIDTH-1:0]  w_in_0_0, w_in_0_1, w_in_0_2, w_in_0_3, w_in_0_4, w_in_0_5, w_in_0_6, w_in_0_7, w_in_0_8, w_in_0_9, w_in_0_10, w_in_0_11, w_in_0_12, w_in_0_13, w_in_0_14, w_in_0_15, w_in_0_16, w_in_0_17, w_in_0_18, w_in_0_19, w_in_0_20, w_in_0_21, w_in_0_22, w_in_0_23, w_in_0_24, w_in_0_25, w_in_0_26, w_in_0_27, w_in_0_28, w_in_0_29, w_in_0_30, w_in_0_31, w_in_0_32, w_in_0_33, w_in_0_34, w_in_0_35, w_in_0_36, w_in_0_37, w_in_0_38, w_in_0_39, w_in_0_40, w_in_0_41, w_in_0_42, w_in_0_43, w_in_0_44, w_in_0_45, w_in_0_46, w_in_0_47, w_in_0_48, w_in_0_49, w_in_0_50, w_in_0_51, w_in_0_52, w_in_0_53, w_in_0_54, w_in_0_55, w_in_0_56, w_in_0_57, w_in_0_58, w_in_0_59, w_in_0_60, w_in_0_61, w_in_0_62, w_in_0_63, w_in_0_64, w_in_0_65, w_in_0_66, w_in_0_67, w_in_0_68, w_in_0_69, w_in_0_70, w_in_0_71, w_in_0_72, w_in_0_73, w_in_0_74, w_in_0_75, w_in_0_76, w_in_0_77, w_in_0_78, w_in_0_79, w_in_0_80, w_in_0_81, w_in_0_82, w_in_0_83, w_in_0_84, w_in_0_85, w_in_0_86, w_in_0_87, w_in_0_88, w_in_0_89, w_in_0_90, w_in_0_91, w_in_0_92, w_in_0_93, w_in_0_94, w_in_0_95, w_in_0_96, w_in_0_97, w_in_0_98, w_in_0_99, w_in_0_100, w_in_0_101, w_in_0_102, w_in_0_103, w_in_0_104, w_in_0_105, w_in_0_106, w_in_0_107, w_in_0_108, w_in_0_109, w_in_0_110, w_in_0_111, w_in_0_112, w_in_0_113, w_in_0_114, w_in_0_115, w_in_0_116, w_in_0_117, w_in_0_118, w_in_0_119, w_in_0_120, w_in_0_121, w_in_0_122, w_in_0_123, w_in_0_124, w_in_0_125, w_in_0_126, w_in_0_127, w_in_0_128, w_in_0_129, w_in_0_130, w_in_0_131, w_in_0_132, w_in_0_133, w_in_0_134, w_in_0_135, w_in_0_136, w_in_0_137, w_in_0_138, w_in_0_139, w_in_0_140, w_in_0_141, w_in_0_142, w_in_0_143, w_in_0_144, w_in_0_145, w_in_0_146, w_in_0_147, w_in_0_148, w_in_0_149, w_in_0_150, w_in_0_151, w_in_0_152, w_in_0_153, w_in_0_154, w_in_0_155, w_in_0_156, w_in_0_157, w_in_0_158, w_in_0_159, w_in_0_160, w_in_0_161, w_in_0_162, w_in_0_163, w_in_0_164, w_in_0_165, w_in_0_166, w_in_0_167, w_in_0_168, w_in_0_169, w_in_0_170, w_in_0_171, w_in_0_172, w_in_0_173, w_in_0_174, w_in_0_175, w_in_0_176, w_in_0_177, w_in_0_178, w_in_0_179, w_in_0_180, w_in_0_181, w_in_0_182, w_in_0_183, w_in_0_184, w_in_0_185, w_in_0_186, w_in_0_187, w_in_0_188, w_in_0_189, w_in_0_190, w_in_0_191, w_in_0_192, w_in_0_193, w_in_0_194, w_in_0_195, w_in_0_196, w_in_0_197, w_in_0_198, w_in_0_199, w_in_0_200, w_in_0_201, w_in_0_202, w_in_0_203, w_in_0_204, w_in_0_205, w_in_0_206, w_in_0_207, w_in_0_208, w_in_0_209, w_in_0_210, w_in_0_211, w_in_0_212, w_in_0_213, w_in_0_214, w_in_0_215, w_in_0_216, w_in_0_217, w_in_0_218, w_in_0_219, w_in_0_220, w_in_0_221, w_in_0_222, w_in_0_223, w_in_0_224, w_in_0_225, w_in_0_226, w_in_0_227, w_in_0_228, w_in_0_229, w_in_0_230, w_in_0_231, w_in_0_232, w_in_0_233, w_in_0_234, w_in_0_235, w_in_0_236, w_in_0_237, w_in_0_238, w_in_0_239, w_in_0_240, w_in_0_241, w_in_0_242, w_in_0_243, w_in_0_244, w_in_0_245, w_in_0_246, w_in_0_247, w_in_0_248, w_in_0_249, w_in_0_250, w_in_0_251, w_in_0_252, w_in_0_253, w_in_0_254, w_in_0_255, w_in_1_0, w_in_1_1, w_in_1_2, w_in_1_3, w_in_1_4, w_in_1_5, w_in_1_6, w_in_1_7, w_in_1_8, w_in_1_9, w_in_1_10, w_in_1_11, w_in_1_12, w_in_1_13, w_in_1_14, w_in_1_15, w_in_1_16, w_in_1_17, w_in_1_18, w_in_1_19, w_in_1_20, w_in_1_21, w_in_1_22, w_in_1_23, w_in_1_24, w_in_1_25, w_in_1_26, w_in_1_27, w_in_1_28, w_in_1_29, w_in_1_30, w_in_1_31, w_in_1_32, w_in_1_33, w_in_1_34, w_in_1_35, w_in_1_36, w_in_1_37, w_in_1_38, w_in_1_39, w_in_1_40, w_in_1_41, w_in_1_42, w_in_1_43, w_in_1_44, w_in_1_45, w_in_1_46, w_in_1_47, w_in_1_48, w_in_1_49, w_in_1_50, w_in_1_51, w_in_1_52, w_in_1_53, w_in_1_54, w_in_1_55, w_in_1_56, w_in_1_57, w_in_1_58, w_in_1_59, w_in_1_60, w_in_1_61, w_in_1_62, w_in_1_63, w_in_1_64, w_in_1_65, w_in_1_66, w_in_1_67, w_in_1_68, w_in_1_69, w_in_1_70, w_in_1_71, w_in_1_72, w_in_1_73, w_in_1_74, w_in_1_75, w_in_1_76, w_in_1_77, w_in_1_78, w_in_1_79, w_in_1_80, w_in_1_81, w_in_1_82, w_in_1_83, w_in_1_84, w_in_1_85, w_in_1_86, w_in_1_87, w_in_1_88, w_in_1_89, w_in_1_90, w_in_1_91, w_in_1_92, w_in_1_93, w_in_1_94, w_in_1_95, w_in_1_96, w_in_1_97, w_in_1_98, w_in_1_99, w_in_1_100, w_in_1_101, w_in_1_102, w_in_1_103, w_in_1_104, w_in_1_105, w_in_1_106, w_in_1_107, w_in_1_108, w_in_1_109, w_in_1_110, w_in_1_111, w_in_1_112, w_in_1_113, w_in_1_114, w_in_1_115, w_in_1_116, w_in_1_117, w_in_1_118, w_in_1_119, w_in_1_120, w_in_1_121, w_in_1_122, w_in_1_123, w_in_1_124, w_in_1_125, w_in_1_126, w_in_1_127, w_in_1_128, w_in_1_129, w_in_1_130, w_in_1_131, w_in_1_132, w_in_1_133, w_in_1_134, w_in_1_135, w_in_1_136, w_in_1_137, w_in_1_138, w_in_1_139, w_in_1_140, w_in_1_141, w_in_1_142, w_in_1_143, w_in_1_144, w_in_1_145, w_in_1_146, w_in_1_147, w_in_1_148, w_in_1_149, w_in_1_150, w_in_1_151, w_in_1_152, w_in_1_153, w_in_1_154, w_in_1_155, w_in_1_156, w_in_1_157, w_in_1_158, w_in_1_159, w_in_1_160, w_in_1_161, w_in_1_162, w_in_1_163, w_in_1_164, w_in_1_165, w_in_1_166, w_in_1_167, w_in_1_168, w_in_1_169, w_in_1_170, w_in_1_171, w_in_1_172, w_in_1_173, w_in_1_174, w_in_1_175, w_in_1_176, w_in_1_177, w_in_1_178, w_in_1_179, w_in_1_180, w_in_1_181, w_in_1_182, w_in_1_183, w_in_1_184, w_in_1_185, w_in_1_186, w_in_1_187, w_in_1_188, w_in_1_189, w_in_1_190, w_in_1_191, w_in_1_192, w_in_1_193, w_in_1_194, w_in_1_195, w_in_1_196, w_in_1_197, w_in_1_198, w_in_1_199, w_in_1_200, w_in_1_201, w_in_1_202, w_in_1_203, w_in_1_204, w_in_1_205, w_in_1_206, w_in_1_207, w_in_1_208, w_in_1_209, w_in_1_210, w_in_1_211, w_in_1_212, w_in_1_213, w_in_1_214, w_in_1_215, w_in_1_216, w_in_1_217, w_in_1_218, w_in_1_219, w_in_1_220, w_in_1_221, w_in_1_222, w_in_1_223, w_in_1_224, w_in_1_225, w_in_1_226, w_in_1_227, w_in_1_228, w_in_1_229, w_in_1_230, w_in_1_231, w_in_1_232, w_in_1_233, w_in_1_234, w_in_1_235, w_in_1_236, w_in_1_237, w_in_1_238, w_in_1_239, w_in_1_240, w_in_1_241, w_in_1_242, w_in_1_243, w_in_1_244, w_in_1_245, w_in_1_246, w_in_1_247, w_in_1_248, w_in_1_249, w_in_1_250, w_in_1_251, w_in_1_252, w_in_1_253, w_in_1_254, w_in_1_255, w_in_2_0, w_in_2_1, w_in_2_2, w_in_2_3, w_in_2_4, w_in_2_5, w_in_2_6, w_in_2_7, w_in_2_8, w_in_2_9, w_in_2_10, w_in_2_11, w_in_2_12, w_in_2_13, w_in_2_14, w_in_2_15, w_in_2_16, w_in_2_17, w_in_2_18, w_in_2_19, w_in_2_20, w_in_2_21, w_in_2_22, w_in_2_23, w_in_2_24, w_in_2_25, w_in_2_26, w_in_2_27, w_in_2_28, w_in_2_29, w_in_2_30, w_in_2_31, w_in_2_32, w_in_2_33, w_in_2_34, w_in_2_35, w_in_2_36, w_in_2_37, w_in_2_38, w_in_2_39, w_in_2_40, w_in_2_41, w_in_2_42, w_in_2_43, w_in_2_44, w_in_2_45, w_in_2_46, w_in_2_47, w_in_2_48, w_in_2_49, w_in_2_50, w_in_2_51, w_in_2_52, w_in_2_53, w_in_2_54, w_in_2_55, w_in_2_56, w_in_2_57, w_in_2_58, w_in_2_59, w_in_2_60, w_in_2_61, w_in_2_62, w_in_2_63, w_in_2_64, w_in_2_65, w_in_2_66, w_in_2_67, w_in_2_68, w_in_2_69, w_in_2_70, w_in_2_71, w_in_2_72, w_in_2_73, w_in_2_74, w_in_2_75, w_in_2_76, w_in_2_77, w_in_2_78, w_in_2_79, w_in_2_80, w_in_2_81, w_in_2_82, w_in_2_83, w_in_2_84, w_in_2_85, w_in_2_86, w_in_2_87, w_in_2_88, w_in_2_89, w_in_2_90, w_in_2_91, w_in_2_92, w_in_2_93, w_in_2_94, w_in_2_95, w_in_2_96, w_in_2_97, w_in_2_98, w_in_2_99, w_in_2_100, w_in_2_101, w_in_2_102, w_in_2_103, w_in_2_104, w_in_2_105, w_in_2_106, w_in_2_107, w_in_2_108, w_in_2_109, w_in_2_110, w_in_2_111, w_in_2_112, w_in_2_113, w_in_2_114, w_in_2_115, w_in_2_116, w_in_2_117, w_in_2_118, w_in_2_119, w_in_2_120, w_in_2_121, w_in_2_122, w_in_2_123, w_in_2_124, w_in_2_125, w_in_2_126, w_in_2_127, w_in_2_128, w_in_2_129, w_in_2_130, w_in_2_131, w_in_2_132, w_in_2_133, w_in_2_134, w_in_2_135, w_in_2_136, w_in_2_137, w_in_2_138, w_in_2_139, w_in_2_140, w_in_2_141, w_in_2_142, w_in_2_143, w_in_2_144, w_in_2_145, w_in_2_146, w_in_2_147, w_in_2_148, w_in_2_149, w_in_2_150, w_in_2_151, w_in_2_152, w_in_2_153, w_in_2_154, w_in_2_155, w_in_2_156, w_in_2_157, w_in_2_158, w_in_2_159, w_in_2_160, w_in_2_161, w_in_2_162, w_in_2_163, w_in_2_164, w_in_2_165, w_in_2_166, w_in_2_167, w_in_2_168, w_in_2_169, w_in_2_170, w_in_2_171, w_in_2_172, w_in_2_173, w_in_2_174, w_in_2_175, w_in_2_176, w_in_2_177, w_in_2_178, w_in_2_179, w_in_2_180, w_in_2_181, w_in_2_182, w_in_2_183, w_in_2_184, w_in_2_185, w_in_2_186, w_in_2_187, w_in_2_188, w_in_2_189, w_in_2_190, w_in_2_191, w_in_2_192, w_in_2_193, w_in_2_194, w_in_2_195, w_in_2_196, w_in_2_197, w_in_2_198, w_in_2_199, w_in_2_200, w_in_2_201, w_in_2_202, w_in_2_203, w_in_2_204, w_in_2_205, w_in_2_206, w_in_2_207, w_in_2_208, w_in_2_209, w_in_2_210, w_in_2_211, w_in_2_212, w_in_2_213, w_in_2_214, w_in_2_215, w_in_2_216, w_in_2_217, w_in_2_218, w_in_2_219, w_in_2_220, w_in_2_221, w_in_2_222, w_in_2_223, w_in_2_224, w_in_2_225, w_in_2_226, w_in_2_227, w_in_2_228, w_in_2_229, w_in_2_230, w_in_2_231, w_in_2_232, w_in_2_233, w_in_2_234, w_in_2_235, w_in_2_236, w_in_2_237, w_in_2_238, w_in_2_239, w_in_2_240, w_in_2_241, w_in_2_242, w_in_2_243, w_in_2_244, w_in_2_245, w_in_2_246, w_in_2_247, w_in_2_248, w_in_2_249, w_in_2_250, w_in_2_251, w_in_2_252, w_in_2_253, w_in_2_254, w_in_2_255, w_in_3_0, w_in_3_1, w_in_3_2, w_in_3_3, w_in_3_4, w_in_3_5, w_in_3_6, w_in_3_7, w_in_3_8, w_in_3_9, w_in_3_10, w_in_3_11, w_in_3_12, w_in_3_13, w_in_3_14, w_in_3_15, w_in_3_16, w_in_3_17, w_in_3_18, w_in_3_19, w_in_3_20, w_in_3_21, w_in_3_22, w_in_3_23, w_in_3_24, w_in_3_25, w_in_3_26, w_in_3_27, w_in_3_28, w_in_3_29, w_in_3_30, w_in_3_31, w_in_3_32, w_in_3_33, w_in_3_34, w_in_3_35, w_in_3_36, w_in_3_37, w_in_3_38, w_in_3_39, w_in_3_40, w_in_3_41, w_in_3_42, w_in_3_43, w_in_3_44, w_in_3_45, w_in_3_46, w_in_3_47, w_in_3_48, w_in_3_49, w_in_3_50, w_in_3_51, w_in_3_52, w_in_3_53, w_in_3_54, w_in_3_55, w_in_3_56, w_in_3_57, w_in_3_58, w_in_3_59, w_in_3_60, w_in_3_61, w_in_3_62, w_in_3_63, w_in_3_64, w_in_3_65, w_in_3_66, w_in_3_67, w_in_3_68, w_in_3_69, w_in_3_70, w_in_3_71, w_in_3_72, w_in_3_73, w_in_3_74, w_in_3_75, w_in_3_76, w_in_3_77, w_in_3_78, w_in_3_79, w_in_3_80, w_in_3_81, w_in_3_82, w_in_3_83, w_in_3_84, w_in_3_85, w_in_3_86, w_in_3_87, w_in_3_88, w_in_3_89, w_in_3_90, w_in_3_91, w_in_3_92, w_in_3_93, w_in_3_94, w_in_3_95, w_in_3_96, w_in_3_97, w_in_3_98, w_in_3_99, w_in_3_100, w_in_3_101, w_in_3_102, w_in_3_103, w_in_3_104, w_in_3_105, w_in_3_106, w_in_3_107, w_in_3_108, w_in_3_109, w_in_3_110, w_in_3_111, w_in_3_112, w_in_3_113, w_in_3_114, w_in_3_115, w_in_3_116, w_in_3_117, w_in_3_118, w_in_3_119, w_in_3_120, w_in_3_121, w_in_3_122, w_in_3_123, w_in_3_124, w_in_3_125, w_in_3_126, w_in_3_127, w_in_3_128, w_in_3_129, w_in_3_130, w_in_3_131, w_in_3_132, w_in_3_133, w_in_3_134, w_in_3_135, w_in_3_136, w_in_3_137, w_in_3_138, w_in_3_139, w_in_3_140, w_in_3_141, w_in_3_142, w_in_3_143, w_in_3_144, w_in_3_145, w_in_3_146, w_in_3_147, w_in_3_148, w_in_3_149, w_in_3_150, w_in_3_151, w_in_3_152, w_in_3_153, w_in_3_154, w_in_3_155, w_in_3_156, w_in_3_157, w_in_3_158, w_in_3_159, w_in_3_160, w_in_3_161, w_in_3_162, w_in_3_163, w_in_3_164, w_in_3_165, w_in_3_166, w_in_3_167, w_in_3_168, w_in_3_169, w_in_3_170, w_in_3_171, w_in_3_172, w_in_3_173, w_in_3_174, w_in_3_175, w_in_3_176, w_in_3_177, w_in_3_178, w_in_3_179, w_in_3_180, w_in_3_181, w_in_3_182, w_in_3_183, w_in_3_184, w_in_3_185, w_in_3_186, w_in_3_187, w_in_3_188, w_in_3_189, w_in_3_190, w_in_3_191, w_in_3_192, w_in_3_193, w_in_3_194, w_in_3_195, w_in_3_196, w_in_3_197, w_in_3_198, w_in_3_199, w_in_3_200, w_in_3_201, w_in_3_202, w_in_3_203, w_in_3_204, w_in_3_205, w_in_3_206, w_in_3_207, w_in_3_208, w_in_3_209, w_in_3_210, w_in_3_211, w_in_3_212, w_in_3_213, w_in_3_214, w_in_3_215, w_in_3_216, w_in_3_217, w_in_3_218, w_in_3_219, w_in_3_220, w_in_3_221, w_in_3_222, w_in_3_223, w_in_3_224, w_in_3_225, w_in_3_226, w_in_3_227, w_in_3_228, w_in_3_229, w_in_3_230, w_in_3_231, w_in_3_232, w_in_3_233, w_in_3_234, w_in_3_235, w_in_3_236, w_in_3_237, w_in_3_238, w_in_3_239, w_in_3_240, w_in_3_241, w_in_3_242, w_in_3_243, w_in_3_244, w_in_3_245, w_in_3_246, w_in_3_247, w_in_3_248, w_in_3_249, w_in_3_250, w_in_3_251, w_in_3_252, w_in_3_253, w_in_3_254, w_in_3_255, w_in_4_0, w_in_4_1, w_in_4_2, w_in_4_3, w_in_4_4, w_in_4_5, w_in_4_6, w_in_4_7, w_in_4_8, w_in_4_9, w_in_4_10, w_in_4_11, w_in_4_12, w_in_4_13, w_in_4_14, w_in_4_15, w_in_4_16, w_in_4_17, w_in_4_18, w_in_4_19, w_in_4_20, w_in_4_21, w_in_4_22, w_in_4_23, w_in_4_24, w_in_4_25, w_in_4_26, w_in_4_27, w_in_4_28, w_in_4_29, w_in_4_30, w_in_4_31, w_in_4_32, w_in_4_33, w_in_4_34, w_in_4_35, w_in_4_36, w_in_4_37, w_in_4_38, w_in_4_39, w_in_4_40, w_in_4_41, w_in_4_42, w_in_4_43, w_in_4_44, w_in_4_45, w_in_4_46, w_in_4_47, w_in_4_48, w_in_4_49, w_in_4_50, w_in_4_51, w_in_4_52, w_in_4_53, w_in_4_54, w_in_4_55, w_in_4_56, w_in_4_57, w_in_4_58, w_in_4_59, w_in_4_60, w_in_4_61, w_in_4_62, w_in_4_63, w_in_4_64, w_in_4_65, w_in_4_66, w_in_4_67, w_in_4_68, w_in_4_69, w_in_4_70, w_in_4_71, w_in_4_72, w_in_4_73, w_in_4_74, w_in_4_75, w_in_4_76, w_in_4_77, w_in_4_78, w_in_4_79, w_in_4_80, w_in_4_81, w_in_4_82, w_in_4_83, w_in_4_84, w_in_4_85, w_in_4_86, w_in_4_87, w_in_4_88, w_in_4_89, w_in_4_90, w_in_4_91, w_in_4_92, w_in_4_93, w_in_4_94, w_in_4_95, w_in_4_96, w_in_4_97, w_in_4_98, w_in_4_99, w_in_4_100, w_in_4_101, w_in_4_102, w_in_4_103, w_in_4_104, w_in_4_105, w_in_4_106, w_in_4_107, w_in_4_108, w_in_4_109, w_in_4_110, w_in_4_111, w_in_4_112, w_in_4_113, w_in_4_114, w_in_4_115, w_in_4_116, w_in_4_117, w_in_4_118, w_in_4_119, w_in_4_120, w_in_4_121, w_in_4_122, w_in_4_123, w_in_4_124, w_in_4_125, w_in_4_126, w_in_4_127, w_in_4_128, w_in_4_129, w_in_4_130, w_in_4_131, w_in_4_132, w_in_4_133, w_in_4_134, w_in_4_135, w_in_4_136, w_in_4_137, w_in_4_138, w_in_4_139, w_in_4_140, w_in_4_141, w_in_4_142, w_in_4_143, w_in_4_144, w_in_4_145, w_in_4_146, w_in_4_147, w_in_4_148, w_in_4_149, w_in_4_150, w_in_4_151, w_in_4_152, w_in_4_153, w_in_4_154, w_in_4_155, w_in_4_156, w_in_4_157, w_in_4_158, w_in_4_159, w_in_4_160, w_in_4_161, w_in_4_162, w_in_4_163, w_in_4_164, w_in_4_165, w_in_4_166, w_in_4_167, w_in_4_168, w_in_4_169, w_in_4_170, w_in_4_171, w_in_4_172, w_in_4_173, w_in_4_174, w_in_4_175, w_in_4_176, w_in_4_177, w_in_4_178, w_in_4_179, w_in_4_180, w_in_4_181, w_in_4_182, w_in_4_183, w_in_4_184, w_in_4_185, w_in_4_186, w_in_4_187, w_in_4_188, w_in_4_189, w_in_4_190, w_in_4_191, w_in_4_192, w_in_4_193, w_in_4_194, w_in_4_195, w_in_4_196, w_in_4_197, w_in_4_198, w_in_4_199, w_in_4_200, w_in_4_201, w_in_4_202, w_in_4_203, w_in_4_204, w_in_4_205, w_in_4_206, w_in_4_207, w_in_4_208, w_in_4_209, w_in_4_210, w_in_4_211, w_in_4_212, w_in_4_213, w_in_4_214, w_in_4_215, w_in_4_216, w_in_4_217, w_in_4_218, w_in_4_219, w_in_4_220, w_in_4_221, w_in_4_222, w_in_4_223, w_in_4_224, w_in_4_225, w_in_4_226, w_in_4_227, w_in_4_228, w_in_4_229, w_in_4_230, w_in_4_231, w_in_4_232, w_in_4_233, w_in_4_234, w_in_4_235, w_in_4_236, w_in_4_237, w_in_4_238, w_in_4_239, w_in_4_240, w_in_4_241, w_in_4_242, w_in_4_243, w_in_4_244, w_in_4_245, w_in_4_246, w_in_4_247, w_in_4_248, w_in_4_249, w_in_4_250, w_in_4_251, w_in_4_252, w_in_4_253, w_in_4_254, w_in_4_255, w_in_5_0, w_in_5_1, w_in_5_2, w_in_5_3, w_in_5_4, w_in_5_5, w_in_5_6, w_in_5_7, w_in_5_8, w_in_5_9, w_in_5_10, w_in_5_11, w_in_5_12, w_in_5_13, w_in_5_14, w_in_5_15, w_in_5_16, w_in_5_17, w_in_5_18, w_in_5_19, w_in_5_20, w_in_5_21, w_in_5_22, w_in_5_23, w_in_5_24, w_in_5_25, w_in_5_26, w_in_5_27, w_in_5_28, w_in_5_29, w_in_5_30, w_in_5_31, w_in_5_32, w_in_5_33, w_in_5_34, w_in_5_35, w_in_5_36, w_in_5_37, w_in_5_38, w_in_5_39, w_in_5_40, w_in_5_41, w_in_5_42, w_in_5_43, w_in_5_44, w_in_5_45, w_in_5_46, w_in_5_47, w_in_5_48, w_in_5_49, w_in_5_50, w_in_5_51, w_in_5_52, w_in_5_53, w_in_5_54, w_in_5_55, w_in_5_56, w_in_5_57, w_in_5_58, w_in_5_59, w_in_5_60, w_in_5_61, w_in_5_62, w_in_5_63, w_in_5_64, w_in_5_65, w_in_5_66, w_in_5_67, w_in_5_68, w_in_5_69, w_in_5_70, w_in_5_71, w_in_5_72, w_in_5_73, w_in_5_74, w_in_5_75, w_in_5_76, w_in_5_77, w_in_5_78, w_in_5_79, w_in_5_80, w_in_5_81, w_in_5_82, w_in_5_83, w_in_5_84, w_in_5_85, w_in_5_86, w_in_5_87, w_in_5_88, w_in_5_89, w_in_5_90, w_in_5_91, w_in_5_92, w_in_5_93, w_in_5_94, w_in_5_95, w_in_5_96, w_in_5_97, w_in_5_98, w_in_5_99, w_in_5_100, w_in_5_101, w_in_5_102, w_in_5_103, w_in_5_104, w_in_5_105, w_in_5_106, w_in_5_107, w_in_5_108, w_in_5_109, w_in_5_110, w_in_5_111, w_in_5_112, w_in_5_113, w_in_5_114, w_in_5_115, w_in_5_116, w_in_5_117, w_in_5_118, w_in_5_119, w_in_5_120, w_in_5_121, w_in_5_122, w_in_5_123, w_in_5_124, w_in_5_125, w_in_5_126, w_in_5_127, w_in_5_128, w_in_5_129, w_in_5_130, w_in_5_131, w_in_5_132, w_in_5_133, w_in_5_134, w_in_5_135, w_in_5_136, w_in_5_137, w_in_5_138, w_in_5_139, w_in_5_140, w_in_5_141, w_in_5_142, w_in_5_143, w_in_5_144, w_in_5_145, w_in_5_146, w_in_5_147, w_in_5_148, w_in_5_149, w_in_5_150, w_in_5_151, w_in_5_152, w_in_5_153, w_in_5_154, w_in_5_155, w_in_5_156, w_in_5_157, w_in_5_158, w_in_5_159, w_in_5_160, w_in_5_161, w_in_5_162, w_in_5_163, w_in_5_164, w_in_5_165, w_in_5_166, w_in_5_167, w_in_5_168, w_in_5_169, w_in_5_170, w_in_5_171, w_in_5_172, w_in_5_173, w_in_5_174, w_in_5_175, w_in_5_176, w_in_5_177, w_in_5_178, w_in_5_179, w_in_5_180, w_in_5_181, w_in_5_182, w_in_5_183, w_in_5_184, w_in_5_185, w_in_5_186, w_in_5_187, w_in_5_188, w_in_5_189, w_in_5_190, w_in_5_191, w_in_5_192, w_in_5_193, w_in_5_194, w_in_5_195, w_in_5_196, w_in_5_197, w_in_5_198, w_in_5_199, w_in_5_200, w_in_5_201, w_in_5_202, w_in_5_203, w_in_5_204, w_in_5_205, w_in_5_206, w_in_5_207, w_in_5_208, w_in_5_209, w_in_5_210, w_in_5_211, w_in_5_212, w_in_5_213, w_in_5_214, w_in_5_215, w_in_5_216, w_in_5_217, w_in_5_218, w_in_5_219, w_in_5_220, w_in_5_221, w_in_5_222, w_in_5_223, w_in_5_224, w_in_5_225, w_in_5_226, w_in_5_227, w_in_5_228, w_in_5_229, w_in_5_230, w_in_5_231, w_in_5_232, w_in_5_233, w_in_5_234, w_in_5_235, w_in_5_236, w_in_5_237, w_in_5_238, w_in_5_239, w_in_5_240, w_in_5_241, w_in_5_242, w_in_5_243, w_in_5_244, w_in_5_245, w_in_5_246, w_in_5_247, w_in_5_248, w_in_5_249, w_in_5_250, w_in_5_251, w_in_5_252, w_in_5_253, w_in_5_254, w_in_5_255, w_in_6_0, w_in_6_1, w_in_6_2, w_in_6_3, w_in_6_4, w_in_6_5, w_in_6_6, w_in_6_7, w_in_6_8, w_in_6_9, w_in_6_10, w_in_6_11, w_in_6_12, w_in_6_13, w_in_6_14, w_in_6_15, w_in_6_16, w_in_6_17, w_in_6_18, w_in_6_19, w_in_6_20, w_in_6_21, w_in_6_22, w_in_6_23, w_in_6_24, w_in_6_25, w_in_6_26, w_in_6_27, w_in_6_28, w_in_6_29, w_in_6_30, w_in_6_31, w_in_6_32, w_in_6_33, w_in_6_34, w_in_6_35, w_in_6_36, w_in_6_37, w_in_6_38, w_in_6_39, w_in_6_40, w_in_6_41, w_in_6_42, w_in_6_43, w_in_6_44, w_in_6_45, w_in_6_46, w_in_6_47, w_in_6_48, w_in_6_49, w_in_6_50, w_in_6_51, w_in_6_52, w_in_6_53, w_in_6_54, w_in_6_55, w_in_6_56, w_in_6_57, w_in_6_58, w_in_6_59, w_in_6_60, w_in_6_61, w_in_6_62, w_in_6_63, w_in_6_64, w_in_6_65, w_in_6_66, w_in_6_67, w_in_6_68, w_in_6_69, w_in_6_70, w_in_6_71, w_in_6_72, w_in_6_73, w_in_6_74, w_in_6_75, w_in_6_76, w_in_6_77, w_in_6_78, w_in_6_79, w_in_6_80, w_in_6_81, w_in_6_82, w_in_6_83, w_in_6_84, w_in_6_85, w_in_6_86, w_in_6_87, w_in_6_88, w_in_6_89, w_in_6_90, w_in_6_91, w_in_6_92, w_in_6_93, w_in_6_94, w_in_6_95, w_in_6_96, w_in_6_97, w_in_6_98, w_in_6_99, w_in_6_100, w_in_6_101, w_in_6_102, w_in_6_103, w_in_6_104, w_in_6_105, w_in_6_106, w_in_6_107, w_in_6_108, w_in_6_109, w_in_6_110, w_in_6_111, w_in_6_112, w_in_6_113, w_in_6_114, w_in_6_115, w_in_6_116, w_in_6_117, w_in_6_118, w_in_6_119, w_in_6_120, w_in_6_121, w_in_6_122, w_in_6_123, w_in_6_124, w_in_6_125, w_in_6_126, w_in_6_127, w_in_6_128, w_in_6_129, w_in_6_130, w_in_6_131, w_in_6_132, w_in_6_133, w_in_6_134, w_in_6_135, w_in_6_136, w_in_6_137, w_in_6_138, w_in_6_139, w_in_6_140, w_in_6_141, w_in_6_142, w_in_6_143, w_in_6_144, w_in_6_145, w_in_6_146, w_in_6_147, w_in_6_148, w_in_6_149, w_in_6_150, w_in_6_151, w_in_6_152, w_in_6_153, w_in_6_154, w_in_6_155, w_in_6_156, w_in_6_157, w_in_6_158, w_in_6_159, w_in_6_160, w_in_6_161, w_in_6_162, w_in_6_163, w_in_6_164, w_in_6_165, w_in_6_166, w_in_6_167, w_in_6_168, w_in_6_169, w_in_6_170, w_in_6_171, w_in_6_172, w_in_6_173, w_in_6_174, w_in_6_175, w_in_6_176, w_in_6_177, w_in_6_178, w_in_6_179, w_in_6_180, w_in_6_181, w_in_6_182, w_in_6_183, w_in_6_184, w_in_6_185, w_in_6_186, w_in_6_187, w_in_6_188, w_in_6_189, w_in_6_190, w_in_6_191, w_in_6_192, w_in_6_193, w_in_6_194, w_in_6_195, w_in_6_196, w_in_6_197, w_in_6_198, w_in_6_199, w_in_6_200, w_in_6_201, w_in_6_202, w_in_6_203, w_in_6_204, w_in_6_205, w_in_6_206, w_in_6_207, w_in_6_208, w_in_6_209, w_in_6_210, w_in_6_211, w_in_6_212, w_in_6_213, w_in_6_214, w_in_6_215, w_in_6_216, w_in_6_217, w_in_6_218, w_in_6_219, w_in_6_220, w_in_6_221, w_in_6_222, w_in_6_223, w_in_6_224, w_in_6_225, w_in_6_226, w_in_6_227, w_in_6_228, w_in_6_229, w_in_6_230, w_in_6_231, w_in_6_232, w_in_6_233, w_in_6_234, w_in_6_235, w_in_6_236, w_in_6_237, w_in_6_238, w_in_6_239, w_in_6_240, w_in_6_241, w_in_6_242, w_in_6_243, w_in_6_244, w_in_6_245, w_in_6_246, w_in_6_247, w_in_6_248, w_in_6_249, w_in_6_250, w_in_6_251, w_in_6_252, w_in_6_253, w_in_6_254, w_in_6_255, w_in_7_0, w_in_7_1, w_in_7_2, w_in_7_3, w_in_7_4, w_in_7_5, w_in_7_6, w_in_7_7, w_in_7_8, w_in_7_9, w_in_7_10, w_in_7_11, w_in_7_12, w_in_7_13, w_in_7_14, w_in_7_15, w_in_7_16, w_in_7_17, w_in_7_18, w_in_7_19, w_in_7_20, w_in_7_21, w_in_7_22, w_in_7_23, w_in_7_24, w_in_7_25, w_in_7_26, w_in_7_27, w_in_7_28, w_in_7_29, w_in_7_30, w_in_7_31, w_in_7_32, w_in_7_33, w_in_7_34, w_in_7_35, w_in_7_36, w_in_7_37, w_in_7_38, w_in_7_39, w_in_7_40, w_in_7_41, w_in_7_42, w_in_7_43, w_in_7_44, w_in_7_45, w_in_7_46, w_in_7_47, w_in_7_48, w_in_7_49, w_in_7_50, w_in_7_51, w_in_7_52, w_in_7_53, w_in_7_54, w_in_7_55, w_in_7_56, w_in_7_57, w_in_7_58, w_in_7_59, w_in_7_60, w_in_7_61, w_in_7_62, w_in_7_63, w_in_7_64, w_in_7_65, w_in_7_66, w_in_7_67, w_in_7_68, w_in_7_69, w_in_7_70, w_in_7_71, w_in_7_72, w_in_7_73, w_in_7_74, w_in_7_75, w_in_7_76, w_in_7_77, w_in_7_78, w_in_7_79, w_in_7_80, w_in_7_81, w_in_7_82, w_in_7_83, w_in_7_84, w_in_7_85, w_in_7_86, w_in_7_87, w_in_7_88, w_in_7_89, w_in_7_90, w_in_7_91, w_in_7_92, w_in_7_93, w_in_7_94, w_in_7_95, w_in_7_96, w_in_7_97, w_in_7_98, w_in_7_99, w_in_7_100, w_in_7_101, w_in_7_102, w_in_7_103, w_in_7_104, w_in_7_105, w_in_7_106, w_in_7_107, w_in_7_108, w_in_7_109, w_in_7_110, w_in_7_111, w_in_7_112, w_in_7_113, w_in_7_114, w_in_7_115, w_in_7_116, w_in_7_117, w_in_7_118, w_in_7_119, w_in_7_120, w_in_7_121, w_in_7_122, w_in_7_123, w_in_7_124, w_in_7_125, w_in_7_126, w_in_7_127, w_in_7_128, w_in_7_129, w_in_7_130, w_in_7_131, w_in_7_132, w_in_7_133, w_in_7_134, w_in_7_135, w_in_7_136, w_in_7_137, w_in_7_138, w_in_7_139, w_in_7_140, w_in_7_141, w_in_7_142, w_in_7_143, w_in_7_144, w_in_7_145, w_in_7_146, w_in_7_147, w_in_7_148, w_in_7_149, w_in_7_150, w_in_7_151, w_in_7_152, w_in_7_153, w_in_7_154, w_in_7_155, w_in_7_156, w_in_7_157, w_in_7_158, w_in_7_159, w_in_7_160, w_in_7_161, w_in_7_162, w_in_7_163, w_in_7_164, w_in_7_165, w_in_7_166, w_in_7_167, w_in_7_168, w_in_7_169, w_in_7_170, w_in_7_171, w_in_7_172, w_in_7_173, w_in_7_174, w_in_7_175, w_in_7_176, w_in_7_177, w_in_7_178, w_in_7_179, w_in_7_180, w_in_7_181, w_in_7_182, w_in_7_183, w_in_7_184, w_in_7_185, w_in_7_186, w_in_7_187, w_in_7_188, w_in_7_189, w_in_7_190, w_in_7_191, w_in_7_192, w_in_7_193, w_in_7_194, w_in_7_195, w_in_7_196, w_in_7_197, w_in_7_198, w_in_7_199, w_in_7_200, w_in_7_201, w_in_7_202, w_in_7_203, w_in_7_204, w_in_7_205, w_in_7_206, w_in_7_207, w_in_7_208, w_in_7_209, w_in_7_210, w_in_7_211, w_in_7_212, w_in_7_213, w_in_7_214, w_in_7_215, w_in_7_216, w_in_7_217, w_in_7_218, w_in_7_219, w_in_7_220, w_in_7_221, w_in_7_222, w_in_7_223, w_in_7_224, w_in_7_225, w_in_7_226, w_in_7_227, w_in_7_228, w_in_7_229, w_in_7_230, w_in_7_231, w_in_7_232, w_in_7_233, w_in_7_234, w_in_7_235, w_in_7_236, w_in_7_237, w_in_7_238, w_in_7_239, w_in_7_240, w_in_7_241, w_in_7_242, w_in_7_243, w_in_7_244, w_in_7_245, w_in_7_246, w_in_7_247, w_in_7_248, w_in_7_249, w_in_7_250, w_in_7_251, w_in_7_252, w_in_7_253, w_in_7_254, w_in_7_255,

    // Recurrent weights (h×h for each gate)
    input  logic signed [WIDTH-1:0]  w_hr_0_0, w_hr_0_1, w_hr_0_2, w_hr_0_3, w_hr_0_4, w_hr_0_5, w_hr_0_6, w_hr_0_7, w_hr_1_0, w_hr_1_1, w_hr_1_2, w_hr_1_3, w_hr_1_4, w_hr_1_5, w_hr_1_6, w_hr_1_7, w_hr_2_0, w_hr_2_1, w_hr_2_2, w_hr_2_3, w_hr_2_4, w_hr_2_5, w_hr_2_6, w_hr_2_7, w_hr_3_0, w_hr_3_1, w_hr_3_2, w_hr_3_3, w_hr_3_4, w_hr_3_5, w_hr_3_6, w_hr_3_7, w_hr_4_0, w_hr_4_1, w_hr_4_2, w_hr_4_3, w_hr_4_4, w_hr_4_5, w_hr_4_6, w_hr_4_7, w_hr_5_0, w_hr_5_1, w_hr_5_2, w_hr_5_3, w_hr_5_4, w_hr_5_5, w_hr_5_6, w_hr_5_7, w_hr_6_0, w_hr_6_1, w_hr_6_2, w_hr_6_3, w_hr_6_4, w_hr_6_5, w_hr_6_6, w_hr_6_7, w_hr_7_0, w_hr_7_1, w_hr_7_2, w_hr_7_3, w_hr_7_4, w_hr_7_5, w_hr_7_6, w_hr_7_7,
    input  logic signed [WIDTH-1:0]  w_hz_0_0, w_hz_0_1, w_hz_0_2, w_hz_0_3, w_hz_0_4, w_hz_0_5, w_hz_0_6, w_hz_0_7, w_hz_1_0, w_hz_1_1, w_hz_1_2, w_hz_1_3, w_hz_1_4, w_hz_1_5, w_hz_1_6, w_hz_1_7, w_hz_2_0, w_hz_2_1, w_hz_2_2, w_hz_2_3, w_hz_2_4, w_hz_2_5, w_hz_2_6, w_hz_2_7, w_hz_3_0, w_hz_3_1, w_hz_3_2, w_hz_3_3, w_hz_3_4, w_hz_3_5, w_hz_3_6, w_hz_3_7, w_hz_4_0, w_hz_4_1, w_hz_4_2, w_hz_4_3, w_hz_4_4, w_hz_4_5, w_hz_4_6, w_hz_4_7, w_hz_5_0, w_hz_5_1, w_hz_5_2, w_hz_5_3, w_hz_5_4, w_hz_5_5, w_hz_5_6, w_hz_5_7, w_hz_6_0, w_hz_6_1, w_hz_6_2, w_hz_6_3, w_hz_6_4, w_hz_6_5, w_hz_6_6, w_hz_6_7, w_hz_7_0, w_hz_7_1, w_hz_7_2, w_hz_7_3, w_hz_7_4, w_hz_7_5, w_hz_7_6, w_hz_7_7,
    input  logic signed [WIDTH-1:0]  w_hn_0_0, w_hn_0_1, w_hn_0_2, w_hn_0_3, w_hn_0_4, w_hn_0_5, w_hn_0_6, w_hn_0_7, w_hn_1_0, w_hn_1_1, w_hn_1_2, w_hn_1_3, w_hn_1_4, w_hn_1_5, w_hn_1_6, w_hn_1_7, w_hn_2_0, w_hn_2_1, w_hn_2_2, w_hn_2_3, w_hn_2_4, w_hn_2_5, w_hn_2_6, w_hn_2_7, w_hn_3_0, w_hn_3_1, w_hn_3_2, w_hn_3_3, w_hn_3_4, w_hn_3_5, w_hn_3_6, w_hn_3_7, w_hn_4_0, w_hn_4_1, w_hn_4_2, w_hn_4_3, w_hn_4_4, w_hn_4_5, w_hn_4_6, w_hn_4_7, w_hn_5_0, w_hn_5_1, w_hn_5_2, w_hn_5_3, w_hn_5_4, w_hn_5_5, w_hn_5_6, w_hn_5_7, w_hn_6_0, w_hn_6_1, w_hn_6_2, w_hn_6_3, w_hn_6_4, w_hn_6_5, w_hn_6_6, w_hn_6_7, w_hn_7_0, w_hn_7_1, w_hn_7_2, w_hn_7_3, w_hn_7_4, w_hn_7_5, w_hn_7_6, w_hn_7_7,

    // Biases (h for each gate type)
    input  logic signed [WIDTH-1:0]  b_ir_0, b_ir_1, b_ir_2, b_ir_3, b_ir_4, b_ir_5, b_ir_6, b_ir_7, b_iz_0, b_iz_1, b_iz_2, b_iz_3, b_iz_4, b_iz_5, b_iz_6, b_iz_7, b_in_0, b_in_1, b_in_2, b_in_3, b_in_4, b_in_5, b_in_6, b_in_7, b_hr_0, b_hr_1, b_hr_2, b_hr_3, b_hr_4, b_hr_5, b_hr_6, b_hr_7, b_hz_0, b_hz_1, b_hz_2, b_hz_3, b_hz_4, b_hz_5, b_hz_6, b_hz_7, b_hn_0, b_hn_1, b_hn_2, b_hn_3, b_hn_4, b_hn_5, b_hn_6, b_hn_7,

    // Outputs (h=8)
        output logic signed [WIDTH-1:0]  y_0,
    output logic signed [WIDTH-1:0]  y_1,
    output logic signed [WIDTH-1:0]  y_2,
    output logic signed [WIDTH-1:0]  y_3,
    output logic signed [WIDTH-1:0]  y_4,
    output logic signed [WIDTH-1:0]  y_5,
    output logic signed [WIDTH-1:0]  y_6,
    output logic signed [WIDTH-1:0]  y_7
);

    // Helper functions
    function automatic logic signed [WIDTH-1:0] sat_add(
        input logic signed [WIDTH-1:0] a,
        input logic signed [WIDTH-1:0] b
    );
        logic signed [WIDTH:0] sum_ext;
        sum_ext = {a[WIDTH-1], a} + {b[WIDTH-1], b};

        if (sum_ext[WIDTH] != sum_ext[WIDTH-1]) begin
            sat_add = sum_ext[WIDTH] ? {1'b1, {(WIDTH-1){1'b0}}} : {1'b0, {(WIDTH-1){1'b1}}};
        end else begin
            sat_add = sum_ext[WIDTH-1:0];
        end
    endfunction

    function automatic logic signed [WIDTH-1:0] fx_mult_round(
        input logic signed [WIDTH-1:0] a,
        input logic signed [WIDTH-1:0] b
    );
        logic signed [(2*WIDTH)-1:0] product;
        logic signed [WIDTH:0] rounded;

        product = a * b;
        rounded = (product[(2*WIDTH)-1:FRAC_WIDTH] + product[FRAC_WIDTH-1]);

        if (rounded[WIDTH] != rounded[WIDTH-1]) begin
            fx_mult_round = rounded[WIDTH] ? {1'b1, {(WIDTH-1){1'b0}}} : {1'b0, {(WIDTH-1){1'b1}}};
        end else begin
            fx_mult_round = rounded[WIDTH-1:0];
        end
    endfunction

    localparam logic signed [WIDTH-1:0] ONE = (1 <<< FRAC_WIDTH);

    // Reset gate: r_t = σ(W_ir*x + b_ir + W_hr*h + b_hr)
    // r gate computation
    logic signed [WIDTH-1:0] r_sum[8];
    logic signed [WIDTH-1:0] r_act[8];

    always_comb begin
        // r_sum[0]
        r_sum[0] = b_ir_0;
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_0, x_0));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_1, x_1));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_2, x_2));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_3, x_3));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_4, x_4));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_5, x_5));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_6, x_6));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_7, x_7));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_8, x_8));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_9, x_9));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_10, x_10));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_11, x_11));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_12, x_12));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_13, x_13));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_14, x_14));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_15, x_15));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_16, x_16));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_17, x_17));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_18, x_18));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_19, x_19));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_20, x_20));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_21, x_21));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_22, x_22));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_23, x_23));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_24, x_24));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_25, x_25));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_26, x_26));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_27, x_27));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_28, x_28));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_29, x_29));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_30, x_30));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_31, x_31));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_32, x_32));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_33, x_33));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_34, x_34));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_35, x_35));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_36, x_36));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_37, x_37));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_38, x_38));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_39, x_39));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_40, x_40));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_41, x_41));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_42, x_42));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_43, x_43));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_44, x_44));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_45, x_45));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_46, x_46));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_47, x_47));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_48, x_48));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_49, x_49));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_50, x_50));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_51, x_51));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_52, x_52));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_53, x_53));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_54, x_54));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_55, x_55));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_56, x_56));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_57, x_57));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_58, x_58));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_59, x_59));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_60, x_60));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_61, x_61));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_62, x_62));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_63, x_63));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_64, x_64));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_65, x_65));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_66, x_66));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_67, x_67));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_68, x_68));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_69, x_69));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_70, x_70));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_71, x_71));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_72, x_72));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_73, x_73));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_74, x_74));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_75, x_75));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_76, x_76));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_77, x_77));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_78, x_78));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_79, x_79));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_80, x_80));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_81, x_81));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_82, x_82));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_83, x_83));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_84, x_84));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_85, x_85));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_86, x_86));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_87, x_87));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_88, x_88));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_89, x_89));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_90, x_90));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_91, x_91));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_92, x_92));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_93, x_93));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_94, x_94));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_95, x_95));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_96, x_96));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_97, x_97));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_98, x_98));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_99, x_99));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_100, x_100));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_101, x_101));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_102, x_102));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_103, x_103));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_104, x_104));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_105, x_105));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_106, x_106));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_107, x_107));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_108, x_108));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_109, x_109));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_110, x_110));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_111, x_111));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_112, x_112));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_113, x_113));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_114, x_114));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_115, x_115));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_116, x_116));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_117, x_117));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_118, x_118));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_119, x_119));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_120, x_120));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_121, x_121));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_122, x_122));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_123, x_123));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_124, x_124));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_125, x_125));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_126, x_126));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_127, x_127));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_128, x_128));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_129, x_129));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_130, x_130));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_131, x_131));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_132, x_132));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_133, x_133));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_134, x_134));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_135, x_135));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_136, x_136));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_137, x_137));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_138, x_138));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_139, x_139));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_140, x_140));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_141, x_141));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_142, x_142));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_143, x_143));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_144, x_144));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_145, x_145));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_146, x_146));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_147, x_147));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_148, x_148));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_149, x_149));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_150, x_150));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_151, x_151));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_152, x_152));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_153, x_153));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_154, x_154));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_155, x_155));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_156, x_156));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_157, x_157));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_158, x_158));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_159, x_159));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_160, x_160));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_161, x_161));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_162, x_162));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_163, x_163));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_164, x_164));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_165, x_165));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_166, x_166));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_167, x_167));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_168, x_168));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_169, x_169));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_170, x_170));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_171, x_171));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_172, x_172));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_173, x_173));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_174, x_174));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_175, x_175));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_176, x_176));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_177, x_177));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_178, x_178));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_179, x_179));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_180, x_180));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_181, x_181));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_182, x_182));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_183, x_183));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_184, x_184));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_185, x_185));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_186, x_186));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_187, x_187));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_188, x_188));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_189, x_189));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_190, x_190));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_191, x_191));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_192, x_192));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_193, x_193));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_194, x_194));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_195, x_195));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_196, x_196));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_197, x_197));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_198, x_198));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_199, x_199));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_200, x_200));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_201, x_201));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_202, x_202));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_203, x_203));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_204, x_204));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_205, x_205));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_206, x_206));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_207, x_207));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_208, x_208));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_209, x_209));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_210, x_210));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_211, x_211));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_212, x_212));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_213, x_213));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_214, x_214));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_215, x_215));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_216, x_216));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_217, x_217));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_218, x_218));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_219, x_219));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_220, x_220));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_221, x_221));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_222, x_222));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_223, x_223));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_224, x_224));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_225, x_225));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_226, x_226));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_227, x_227));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_228, x_228));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_229, x_229));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_230, x_230));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_231, x_231));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_232, x_232));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_233, x_233));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_234, x_234));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_235, x_235));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_236, x_236));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_237, x_237));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_238, x_238));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_239, x_239));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_240, x_240));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_241, x_241));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_242, x_242));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_243, x_243));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_244, x_244));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_245, x_245));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_246, x_246));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_247, x_247));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_248, x_248));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_249, x_249));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_250, x_250));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_251, x_251));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_252, x_252));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_253, x_253));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_254, x_254));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_ir_0_255, x_255));
        r_sum[0] = sat_add(r_sum[0], b_hr_0);
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_hr_0_0, h_0));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_hr_0_1, h_1));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_hr_0_2, h_2));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_hr_0_3, h_3));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_hr_0_4, h_4));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_hr_0_5, h_5));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_hr_0_6, h_6));
        r_sum[0] = sat_add(r_sum[0], fx_mult_round(w_hr_0_7, h_7));

        // r_sum[1]
        r_sum[1] = b_ir_1;
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_0, x_0));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_1, x_1));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_2, x_2));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_3, x_3));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_4, x_4));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_5, x_5));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_6, x_6));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_7, x_7));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_8, x_8));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_9, x_9));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_10, x_10));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_11, x_11));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_12, x_12));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_13, x_13));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_14, x_14));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_15, x_15));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_16, x_16));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_17, x_17));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_18, x_18));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_19, x_19));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_20, x_20));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_21, x_21));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_22, x_22));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_23, x_23));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_24, x_24));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_25, x_25));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_26, x_26));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_27, x_27));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_28, x_28));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_29, x_29));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_30, x_30));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_31, x_31));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_32, x_32));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_33, x_33));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_34, x_34));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_35, x_35));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_36, x_36));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_37, x_37));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_38, x_38));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_39, x_39));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_40, x_40));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_41, x_41));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_42, x_42));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_43, x_43));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_44, x_44));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_45, x_45));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_46, x_46));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_47, x_47));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_48, x_48));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_49, x_49));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_50, x_50));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_51, x_51));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_52, x_52));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_53, x_53));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_54, x_54));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_55, x_55));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_56, x_56));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_57, x_57));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_58, x_58));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_59, x_59));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_60, x_60));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_61, x_61));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_62, x_62));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_63, x_63));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_64, x_64));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_65, x_65));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_66, x_66));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_67, x_67));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_68, x_68));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_69, x_69));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_70, x_70));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_71, x_71));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_72, x_72));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_73, x_73));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_74, x_74));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_75, x_75));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_76, x_76));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_77, x_77));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_78, x_78));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_79, x_79));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_80, x_80));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_81, x_81));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_82, x_82));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_83, x_83));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_84, x_84));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_85, x_85));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_86, x_86));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_87, x_87));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_88, x_88));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_89, x_89));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_90, x_90));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_91, x_91));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_92, x_92));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_93, x_93));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_94, x_94));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_95, x_95));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_96, x_96));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_97, x_97));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_98, x_98));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_99, x_99));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_100, x_100));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_101, x_101));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_102, x_102));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_103, x_103));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_104, x_104));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_105, x_105));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_106, x_106));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_107, x_107));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_108, x_108));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_109, x_109));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_110, x_110));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_111, x_111));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_112, x_112));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_113, x_113));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_114, x_114));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_115, x_115));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_116, x_116));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_117, x_117));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_118, x_118));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_119, x_119));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_120, x_120));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_121, x_121));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_122, x_122));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_123, x_123));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_124, x_124));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_125, x_125));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_126, x_126));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_127, x_127));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_128, x_128));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_129, x_129));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_130, x_130));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_131, x_131));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_132, x_132));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_133, x_133));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_134, x_134));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_135, x_135));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_136, x_136));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_137, x_137));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_138, x_138));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_139, x_139));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_140, x_140));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_141, x_141));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_142, x_142));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_143, x_143));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_144, x_144));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_145, x_145));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_146, x_146));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_147, x_147));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_148, x_148));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_149, x_149));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_150, x_150));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_151, x_151));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_152, x_152));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_153, x_153));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_154, x_154));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_155, x_155));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_156, x_156));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_157, x_157));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_158, x_158));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_159, x_159));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_160, x_160));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_161, x_161));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_162, x_162));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_163, x_163));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_164, x_164));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_165, x_165));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_166, x_166));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_167, x_167));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_168, x_168));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_169, x_169));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_170, x_170));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_171, x_171));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_172, x_172));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_173, x_173));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_174, x_174));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_175, x_175));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_176, x_176));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_177, x_177));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_178, x_178));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_179, x_179));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_180, x_180));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_181, x_181));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_182, x_182));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_183, x_183));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_184, x_184));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_185, x_185));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_186, x_186));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_187, x_187));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_188, x_188));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_189, x_189));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_190, x_190));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_191, x_191));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_192, x_192));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_193, x_193));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_194, x_194));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_195, x_195));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_196, x_196));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_197, x_197));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_198, x_198));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_199, x_199));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_200, x_200));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_201, x_201));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_202, x_202));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_203, x_203));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_204, x_204));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_205, x_205));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_206, x_206));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_207, x_207));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_208, x_208));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_209, x_209));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_210, x_210));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_211, x_211));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_212, x_212));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_213, x_213));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_214, x_214));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_215, x_215));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_216, x_216));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_217, x_217));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_218, x_218));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_219, x_219));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_220, x_220));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_221, x_221));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_222, x_222));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_223, x_223));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_224, x_224));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_225, x_225));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_226, x_226));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_227, x_227));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_228, x_228));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_229, x_229));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_230, x_230));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_231, x_231));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_232, x_232));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_233, x_233));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_234, x_234));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_235, x_235));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_236, x_236));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_237, x_237));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_238, x_238));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_239, x_239));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_240, x_240));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_241, x_241));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_242, x_242));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_243, x_243));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_244, x_244));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_245, x_245));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_246, x_246));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_247, x_247));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_248, x_248));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_249, x_249));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_250, x_250));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_251, x_251));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_252, x_252));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_253, x_253));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_254, x_254));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_ir_1_255, x_255));
        r_sum[1] = sat_add(r_sum[1], b_hr_1);
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_hr_1_0, h_0));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_hr_1_1, h_1));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_hr_1_2, h_2));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_hr_1_3, h_3));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_hr_1_4, h_4));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_hr_1_5, h_5));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_hr_1_6, h_6));
        r_sum[1] = sat_add(r_sum[1], fx_mult_round(w_hr_1_7, h_7));

        // r_sum[2]
        r_sum[2] = b_ir_2;
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_0, x_0));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_1, x_1));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_2, x_2));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_3, x_3));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_4, x_4));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_5, x_5));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_6, x_6));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_7, x_7));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_8, x_8));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_9, x_9));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_10, x_10));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_11, x_11));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_12, x_12));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_13, x_13));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_14, x_14));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_15, x_15));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_16, x_16));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_17, x_17));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_18, x_18));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_19, x_19));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_20, x_20));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_21, x_21));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_22, x_22));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_23, x_23));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_24, x_24));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_25, x_25));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_26, x_26));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_27, x_27));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_28, x_28));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_29, x_29));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_30, x_30));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_31, x_31));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_32, x_32));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_33, x_33));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_34, x_34));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_35, x_35));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_36, x_36));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_37, x_37));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_38, x_38));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_39, x_39));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_40, x_40));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_41, x_41));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_42, x_42));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_43, x_43));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_44, x_44));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_45, x_45));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_46, x_46));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_47, x_47));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_48, x_48));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_49, x_49));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_50, x_50));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_51, x_51));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_52, x_52));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_53, x_53));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_54, x_54));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_55, x_55));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_56, x_56));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_57, x_57));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_58, x_58));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_59, x_59));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_60, x_60));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_61, x_61));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_62, x_62));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_63, x_63));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_64, x_64));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_65, x_65));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_66, x_66));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_67, x_67));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_68, x_68));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_69, x_69));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_70, x_70));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_71, x_71));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_72, x_72));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_73, x_73));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_74, x_74));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_75, x_75));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_76, x_76));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_77, x_77));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_78, x_78));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_79, x_79));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_80, x_80));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_81, x_81));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_82, x_82));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_83, x_83));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_84, x_84));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_85, x_85));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_86, x_86));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_87, x_87));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_88, x_88));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_89, x_89));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_90, x_90));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_91, x_91));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_92, x_92));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_93, x_93));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_94, x_94));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_95, x_95));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_96, x_96));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_97, x_97));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_98, x_98));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_99, x_99));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_100, x_100));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_101, x_101));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_102, x_102));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_103, x_103));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_104, x_104));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_105, x_105));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_106, x_106));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_107, x_107));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_108, x_108));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_109, x_109));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_110, x_110));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_111, x_111));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_112, x_112));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_113, x_113));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_114, x_114));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_115, x_115));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_116, x_116));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_117, x_117));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_118, x_118));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_119, x_119));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_120, x_120));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_121, x_121));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_122, x_122));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_123, x_123));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_124, x_124));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_125, x_125));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_126, x_126));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_127, x_127));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_128, x_128));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_129, x_129));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_130, x_130));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_131, x_131));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_132, x_132));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_133, x_133));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_134, x_134));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_135, x_135));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_136, x_136));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_137, x_137));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_138, x_138));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_139, x_139));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_140, x_140));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_141, x_141));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_142, x_142));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_143, x_143));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_144, x_144));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_145, x_145));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_146, x_146));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_147, x_147));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_148, x_148));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_149, x_149));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_150, x_150));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_151, x_151));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_152, x_152));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_153, x_153));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_154, x_154));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_155, x_155));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_156, x_156));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_157, x_157));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_158, x_158));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_159, x_159));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_160, x_160));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_161, x_161));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_162, x_162));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_163, x_163));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_164, x_164));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_165, x_165));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_166, x_166));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_167, x_167));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_168, x_168));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_169, x_169));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_170, x_170));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_171, x_171));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_172, x_172));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_173, x_173));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_174, x_174));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_175, x_175));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_176, x_176));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_177, x_177));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_178, x_178));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_179, x_179));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_180, x_180));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_181, x_181));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_182, x_182));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_183, x_183));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_184, x_184));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_185, x_185));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_186, x_186));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_187, x_187));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_188, x_188));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_189, x_189));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_190, x_190));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_191, x_191));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_192, x_192));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_193, x_193));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_194, x_194));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_195, x_195));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_196, x_196));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_197, x_197));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_198, x_198));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_199, x_199));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_200, x_200));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_201, x_201));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_202, x_202));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_203, x_203));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_204, x_204));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_205, x_205));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_206, x_206));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_207, x_207));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_208, x_208));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_209, x_209));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_210, x_210));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_211, x_211));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_212, x_212));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_213, x_213));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_214, x_214));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_215, x_215));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_216, x_216));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_217, x_217));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_218, x_218));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_219, x_219));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_220, x_220));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_221, x_221));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_222, x_222));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_223, x_223));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_224, x_224));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_225, x_225));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_226, x_226));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_227, x_227));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_228, x_228));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_229, x_229));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_230, x_230));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_231, x_231));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_232, x_232));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_233, x_233));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_234, x_234));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_235, x_235));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_236, x_236));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_237, x_237));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_238, x_238));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_239, x_239));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_240, x_240));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_241, x_241));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_242, x_242));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_243, x_243));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_244, x_244));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_245, x_245));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_246, x_246));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_247, x_247));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_248, x_248));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_249, x_249));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_250, x_250));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_251, x_251));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_252, x_252));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_253, x_253));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_254, x_254));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_ir_2_255, x_255));
        r_sum[2] = sat_add(r_sum[2], b_hr_2);
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_hr_2_0, h_0));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_hr_2_1, h_1));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_hr_2_2, h_2));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_hr_2_3, h_3));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_hr_2_4, h_4));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_hr_2_5, h_5));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_hr_2_6, h_6));
        r_sum[2] = sat_add(r_sum[2], fx_mult_round(w_hr_2_7, h_7));

        // r_sum[3]
        r_sum[3] = b_ir_3;
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_0, x_0));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_1, x_1));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_2, x_2));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_3, x_3));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_4, x_4));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_5, x_5));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_6, x_6));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_7, x_7));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_8, x_8));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_9, x_9));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_10, x_10));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_11, x_11));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_12, x_12));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_13, x_13));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_14, x_14));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_15, x_15));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_16, x_16));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_17, x_17));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_18, x_18));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_19, x_19));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_20, x_20));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_21, x_21));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_22, x_22));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_23, x_23));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_24, x_24));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_25, x_25));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_26, x_26));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_27, x_27));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_28, x_28));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_29, x_29));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_30, x_30));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_31, x_31));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_32, x_32));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_33, x_33));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_34, x_34));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_35, x_35));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_36, x_36));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_37, x_37));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_38, x_38));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_39, x_39));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_40, x_40));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_41, x_41));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_42, x_42));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_43, x_43));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_44, x_44));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_45, x_45));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_46, x_46));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_47, x_47));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_48, x_48));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_49, x_49));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_50, x_50));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_51, x_51));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_52, x_52));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_53, x_53));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_54, x_54));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_55, x_55));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_56, x_56));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_57, x_57));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_58, x_58));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_59, x_59));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_60, x_60));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_61, x_61));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_62, x_62));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_63, x_63));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_64, x_64));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_65, x_65));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_66, x_66));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_67, x_67));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_68, x_68));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_69, x_69));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_70, x_70));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_71, x_71));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_72, x_72));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_73, x_73));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_74, x_74));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_75, x_75));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_76, x_76));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_77, x_77));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_78, x_78));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_79, x_79));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_80, x_80));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_81, x_81));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_82, x_82));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_83, x_83));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_84, x_84));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_85, x_85));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_86, x_86));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_87, x_87));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_88, x_88));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_89, x_89));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_90, x_90));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_91, x_91));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_92, x_92));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_93, x_93));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_94, x_94));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_95, x_95));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_96, x_96));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_97, x_97));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_98, x_98));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_99, x_99));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_100, x_100));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_101, x_101));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_102, x_102));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_103, x_103));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_104, x_104));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_105, x_105));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_106, x_106));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_107, x_107));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_108, x_108));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_109, x_109));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_110, x_110));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_111, x_111));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_112, x_112));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_113, x_113));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_114, x_114));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_115, x_115));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_116, x_116));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_117, x_117));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_118, x_118));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_119, x_119));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_120, x_120));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_121, x_121));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_122, x_122));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_123, x_123));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_124, x_124));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_125, x_125));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_126, x_126));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_127, x_127));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_128, x_128));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_129, x_129));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_130, x_130));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_131, x_131));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_132, x_132));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_133, x_133));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_134, x_134));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_135, x_135));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_136, x_136));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_137, x_137));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_138, x_138));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_139, x_139));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_140, x_140));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_141, x_141));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_142, x_142));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_143, x_143));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_144, x_144));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_145, x_145));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_146, x_146));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_147, x_147));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_148, x_148));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_149, x_149));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_150, x_150));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_151, x_151));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_152, x_152));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_153, x_153));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_154, x_154));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_155, x_155));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_156, x_156));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_157, x_157));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_158, x_158));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_159, x_159));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_160, x_160));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_161, x_161));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_162, x_162));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_163, x_163));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_164, x_164));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_165, x_165));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_166, x_166));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_167, x_167));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_168, x_168));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_169, x_169));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_170, x_170));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_171, x_171));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_172, x_172));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_173, x_173));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_174, x_174));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_175, x_175));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_176, x_176));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_177, x_177));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_178, x_178));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_179, x_179));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_180, x_180));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_181, x_181));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_182, x_182));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_183, x_183));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_184, x_184));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_185, x_185));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_186, x_186));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_187, x_187));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_188, x_188));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_189, x_189));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_190, x_190));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_191, x_191));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_192, x_192));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_193, x_193));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_194, x_194));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_195, x_195));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_196, x_196));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_197, x_197));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_198, x_198));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_199, x_199));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_200, x_200));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_201, x_201));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_202, x_202));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_203, x_203));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_204, x_204));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_205, x_205));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_206, x_206));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_207, x_207));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_208, x_208));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_209, x_209));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_210, x_210));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_211, x_211));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_212, x_212));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_213, x_213));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_214, x_214));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_215, x_215));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_216, x_216));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_217, x_217));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_218, x_218));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_219, x_219));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_220, x_220));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_221, x_221));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_222, x_222));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_223, x_223));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_224, x_224));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_225, x_225));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_226, x_226));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_227, x_227));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_228, x_228));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_229, x_229));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_230, x_230));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_231, x_231));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_232, x_232));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_233, x_233));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_234, x_234));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_235, x_235));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_236, x_236));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_237, x_237));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_238, x_238));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_239, x_239));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_240, x_240));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_241, x_241));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_242, x_242));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_243, x_243));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_244, x_244));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_245, x_245));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_246, x_246));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_247, x_247));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_248, x_248));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_249, x_249));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_250, x_250));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_251, x_251));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_252, x_252));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_253, x_253));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_254, x_254));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_ir_3_255, x_255));
        r_sum[3] = sat_add(r_sum[3], b_hr_3);
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_hr_3_0, h_0));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_hr_3_1, h_1));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_hr_3_2, h_2));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_hr_3_3, h_3));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_hr_3_4, h_4));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_hr_3_5, h_5));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_hr_3_6, h_6));
        r_sum[3] = sat_add(r_sum[3], fx_mult_round(w_hr_3_7, h_7));

        // r_sum[4]
        r_sum[4] = b_ir_4;
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_0, x_0));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_1, x_1));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_2, x_2));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_3, x_3));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_4, x_4));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_5, x_5));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_6, x_6));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_7, x_7));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_8, x_8));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_9, x_9));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_10, x_10));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_11, x_11));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_12, x_12));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_13, x_13));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_14, x_14));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_15, x_15));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_16, x_16));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_17, x_17));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_18, x_18));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_19, x_19));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_20, x_20));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_21, x_21));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_22, x_22));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_23, x_23));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_24, x_24));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_25, x_25));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_26, x_26));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_27, x_27));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_28, x_28));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_29, x_29));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_30, x_30));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_31, x_31));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_32, x_32));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_33, x_33));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_34, x_34));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_35, x_35));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_36, x_36));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_37, x_37));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_38, x_38));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_39, x_39));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_40, x_40));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_41, x_41));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_42, x_42));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_43, x_43));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_44, x_44));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_45, x_45));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_46, x_46));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_47, x_47));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_48, x_48));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_49, x_49));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_50, x_50));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_51, x_51));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_52, x_52));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_53, x_53));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_54, x_54));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_55, x_55));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_56, x_56));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_57, x_57));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_58, x_58));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_59, x_59));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_60, x_60));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_61, x_61));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_62, x_62));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_63, x_63));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_64, x_64));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_65, x_65));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_66, x_66));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_67, x_67));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_68, x_68));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_69, x_69));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_70, x_70));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_71, x_71));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_72, x_72));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_73, x_73));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_74, x_74));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_75, x_75));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_76, x_76));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_77, x_77));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_78, x_78));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_79, x_79));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_80, x_80));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_81, x_81));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_82, x_82));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_83, x_83));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_84, x_84));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_85, x_85));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_86, x_86));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_87, x_87));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_88, x_88));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_89, x_89));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_90, x_90));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_91, x_91));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_92, x_92));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_93, x_93));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_94, x_94));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_95, x_95));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_96, x_96));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_97, x_97));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_98, x_98));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_99, x_99));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_100, x_100));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_101, x_101));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_102, x_102));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_103, x_103));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_104, x_104));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_105, x_105));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_106, x_106));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_107, x_107));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_108, x_108));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_109, x_109));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_110, x_110));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_111, x_111));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_112, x_112));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_113, x_113));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_114, x_114));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_115, x_115));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_116, x_116));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_117, x_117));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_118, x_118));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_119, x_119));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_120, x_120));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_121, x_121));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_122, x_122));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_123, x_123));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_124, x_124));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_125, x_125));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_126, x_126));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_127, x_127));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_128, x_128));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_129, x_129));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_130, x_130));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_131, x_131));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_132, x_132));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_133, x_133));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_134, x_134));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_135, x_135));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_136, x_136));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_137, x_137));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_138, x_138));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_139, x_139));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_140, x_140));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_141, x_141));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_142, x_142));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_143, x_143));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_144, x_144));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_145, x_145));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_146, x_146));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_147, x_147));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_148, x_148));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_149, x_149));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_150, x_150));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_151, x_151));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_152, x_152));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_153, x_153));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_154, x_154));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_155, x_155));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_156, x_156));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_157, x_157));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_158, x_158));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_159, x_159));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_160, x_160));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_161, x_161));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_162, x_162));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_163, x_163));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_164, x_164));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_165, x_165));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_166, x_166));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_167, x_167));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_168, x_168));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_169, x_169));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_170, x_170));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_171, x_171));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_172, x_172));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_173, x_173));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_174, x_174));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_175, x_175));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_176, x_176));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_177, x_177));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_178, x_178));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_179, x_179));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_180, x_180));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_181, x_181));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_182, x_182));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_183, x_183));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_184, x_184));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_185, x_185));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_186, x_186));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_187, x_187));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_188, x_188));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_189, x_189));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_190, x_190));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_191, x_191));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_192, x_192));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_193, x_193));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_194, x_194));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_195, x_195));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_196, x_196));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_197, x_197));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_198, x_198));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_199, x_199));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_200, x_200));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_201, x_201));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_202, x_202));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_203, x_203));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_204, x_204));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_205, x_205));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_206, x_206));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_207, x_207));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_208, x_208));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_209, x_209));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_210, x_210));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_211, x_211));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_212, x_212));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_213, x_213));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_214, x_214));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_215, x_215));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_216, x_216));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_217, x_217));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_218, x_218));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_219, x_219));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_220, x_220));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_221, x_221));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_222, x_222));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_223, x_223));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_224, x_224));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_225, x_225));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_226, x_226));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_227, x_227));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_228, x_228));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_229, x_229));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_230, x_230));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_231, x_231));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_232, x_232));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_233, x_233));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_234, x_234));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_235, x_235));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_236, x_236));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_237, x_237));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_238, x_238));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_239, x_239));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_240, x_240));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_241, x_241));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_242, x_242));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_243, x_243));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_244, x_244));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_245, x_245));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_246, x_246));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_247, x_247));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_248, x_248));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_249, x_249));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_250, x_250));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_251, x_251));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_252, x_252));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_253, x_253));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_254, x_254));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_ir_4_255, x_255));
        r_sum[4] = sat_add(r_sum[4], b_hr_4);
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_hr_4_0, h_0));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_hr_4_1, h_1));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_hr_4_2, h_2));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_hr_4_3, h_3));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_hr_4_4, h_4));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_hr_4_5, h_5));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_hr_4_6, h_6));
        r_sum[4] = sat_add(r_sum[4], fx_mult_round(w_hr_4_7, h_7));

        // r_sum[5]
        r_sum[5] = b_ir_5;
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_0, x_0));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_1, x_1));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_2, x_2));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_3, x_3));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_4, x_4));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_5, x_5));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_6, x_6));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_7, x_7));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_8, x_8));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_9, x_9));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_10, x_10));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_11, x_11));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_12, x_12));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_13, x_13));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_14, x_14));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_15, x_15));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_16, x_16));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_17, x_17));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_18, x_18));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_19, x_19));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_20, x_20));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_21, x_21));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_22, x_22));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_23, x_23));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_24, x_24));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_25, x_25));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_26, x_26));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_27, x_27));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_28, x_28));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_29, x_29));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_30, x_30));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_31, x_31));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_32, x_32));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_33, x_33));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_34, x_34));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_35, x_35));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_36, x_36));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_37, x_37));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_38, x_38));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_39, x_39));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_40, x_40));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_41, x_41));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_42, x_42));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_43, x_43));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_44, x_44));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_45, x_45));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_46, x_46));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_47, x_47));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_48, x_48));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_49, x_49));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_50, x_50));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_51, x_51));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_52, x_52));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_53, x_53));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_54, x_54));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_55, x_55));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_56, x_56));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_57, x_57));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_58, x_58));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_59, x_59));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_60, x_60));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_61, x_61));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_62, x_62));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_63, x_63));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_64, x_64));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_65, x_65));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_66, x_66));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_67, x_67));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_68, x_68));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_69, x_69));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_70, x_70));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_71, x_71));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_72, x_72));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_73, x_73));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_74, x_74));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_75, x_75));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_76, x_76));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_77, x_77));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_78, x_78));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_79, x_79));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_80, x_80));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_81, x_81));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_82, x_82));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_83, x_83));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_84, x_84));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_85, x_85));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_86, x_86));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_87, x_87));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_88, x_88));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_89, x_89));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_90, x_90));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_91, x_91));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_92, x_92));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_93, x_93));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_94, x_94));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_95, x_95));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_96, x_96));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_97, x_97));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_98, x_98));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_99, x_99));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_100, x_100));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_101, x_101));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_102, x_102));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_103, x_103));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_104, x_104));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_105, x_105));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_106, x_106));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_107, x_107));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_108, x_108));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_109, x_109));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_110, x_110));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_111, x_111));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_112, x_112));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_113, x_113));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_114, x_114));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_115, x_115));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_116, x_116));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_117, x_117));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_118, x_118));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_119, x_119));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_120, x_120));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_121, x_121));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_122, x_122));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_123, x_123));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_124, x_124));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_125, x_125));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_126, x_126));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_127, x_127));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_128, x_128));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_129, x_129));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_130, x_130));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_131, x_131));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_132, x_132));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_133, x_133));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_134, x_134));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_135, x_135));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_136, x_136));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_137, x_137));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_138, x_138));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_139, x_139));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_140, x_140));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_141, x_141));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_142, x_142));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_143, x_143));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_144, x_144));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_145, x_145));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_146, x_146));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_147, x_147));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_148, x_148));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_149, x_149));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_150, x_150));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_151, x_151));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_152, x_152));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_153, x_153));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_154, x_154));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_155, x_155));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_156, x_156));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_157, x_157));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_158, x_158));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_159, x_159));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_160, x_160));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_161, x_161));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_162, x_162));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_163, x_163));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_164, x_164));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_165, x_165));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_166, x_166));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_167, x_167));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_168, x_168));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_169, x_169));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_170, x_170));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_171, x_171));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_172, x_172));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_173, x_173));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_174, x_174));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_175, x_175));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_176, x_176));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_177, x_177));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_178, x_178));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_179, x_179));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_180, x_180));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_181, x_181));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_182, x_182));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_183, x_183));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_184, x_184));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_185, x_185));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_186, x_186));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_187, x_187));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_188, x_188));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_189, x_189));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_190, x_190));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_191, x_191));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_192, x_192));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_193, x_193));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_194, x_194));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_195, x_195));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_196, x_196));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_197, x_197));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_198, x_198));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_199, x_199));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_200, x_200));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_201, x_201));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_202, x_202));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_203, x_203));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_204, x_204));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_205, x_205));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_206, x_206));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_207, x_207));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_208, x_208));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_209, x_209));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_210, x_210));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_211, x_211));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_212, x_212));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_213, x_213));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_214, x_214));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_215, x_215));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_216, x_216));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_217, x_217));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_218, x_218));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_219, x_219));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_220, x_220));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_221, x_221));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_222, x_222));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_223, x_223));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_224, x_224));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_225, x_225));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_226, x_226));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_227, x_227));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_228, x_228));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_229, x_229));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_230, x_230));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_231, x_231));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_232, x_232));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_233, x_233));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_234, x_234));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_235, x_235));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_236, x_236));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_237, x_237));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_238, x_238));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_239, x_239));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_240, x_240));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_241, x_241));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_242, x_242));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_243, x_243));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_244, x_244));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_245, x_245));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_246, x_246));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_247, x_247));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_248, x_248));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_249, x_249));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_250, x_250));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_251, x_251));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_252, x_252));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_253, x_253));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_254, x_254));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_ir_5_255, x_255));
        r_sum[5] = sat_add(r_sum[5], b_hr_5);
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_hr_5_0, h_0));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_hr_5_1, h_1));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_hr_5_2, h_2));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_hr_5_3, h_3));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_hr_5_4, h_4));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_hr_5_5, h_5));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_hr_5_6, h_6));
        r_sum[5] = sat_add(r_sum[5], fx_mult_round(w_hr_5_7, h_7));

        // r_sum[6]
        r_sum[6] = b_ir_6;
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_0, x_0));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_1, x_1));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_2, x_2));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_3, x_3));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_4, x_4));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_5, x_5));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_6, x_6));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_7, x_7));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_8, x_8));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_9, x_9));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_10, x_10));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_11, x_11));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_12, x_12));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_13, x_13));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_14, x_14));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_15, x_15));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_16, x_16));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_17, x_17));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_18, x_18));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_19, x_19));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_20, x_20));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_21, x_21));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_22, x_22));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_23, x_23));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_24, x_24));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_25, x_25));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_26, x_26));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_27, x_27));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_28, x_28));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_29, x_29));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_30, x_30));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_31, x_31));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_32, x_32));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_33, x_33));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_34, x_34));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_35, x_35));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_36, x_36));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_37, x_37));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_38, x_38));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_39, x_39));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_40, x_40));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_41, x_41));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_42, x_42));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_43, x_43));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_44, x_44));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_45, x_45));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_46, x_46));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_47, x_47));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_48, x_48));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_49, x_49));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_50, x_50));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_51, x_51));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_52, x_52));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_53, x_53));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_54, x_54));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_55, x_55));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_56, x_56));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_57, x_57));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_58, x_58));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_59, x_59));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_60, x_60));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_61, x_61));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_62, x_62));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_63, x_63));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_64, x_64));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_65, x_65));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_66, x_66));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_67, x_67));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_68, x_68));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_69, x_69));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_70, x_70));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_71, x_71));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_72, x_72));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_73, x_73));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_74, x_74));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_75, x_75));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_76, x_76));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_77, x_77));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_78, x_78));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_79, x_79));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_80, x_80));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_81, x_81));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_82, x_82));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_83, x_83));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_84, x_84));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_85, x_85));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_86, x_86));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_87, x_87));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_88, x_88));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_89, x_89));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_90, x_90));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_91, x_91));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_92, x_92));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_93, x_93));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_94, x_94));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_95, x_95));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_96, x_96));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_97, x_97));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_98, x_98));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_99, x_99));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_100, x_100));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_101, x_101));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_102, x_102));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_103, x_103));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_104, x_104));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_105, x_105));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_106, x_106));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_107, x_107));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_108, x_108));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_109, x_109));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_110, x_110));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_111, x_111));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_112, x_112));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_113, x_113));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_114, x_114));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_115, x_115));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_116, x_116));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_117, x_117));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_118, x_118));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_119, x_119));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_120, x_120));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_121, x_121));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_122, x_122));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_123, x_123));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_124, x_124));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_125, x_125));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_126, x_126));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_127, x_127));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_128, x_128));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_129, x_129));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_130, x_130));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_131, x_131));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_132, x_132));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_133, x_133));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_134, x_134));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_135, x_135));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_136, x_136));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_137, x_137));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_138, x_138));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_139, x_139));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_140, x_140));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_141, x_141));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_142, x_142));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_143, x_143));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_144, x_144));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_145, x_145));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_146, x_146));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_147, x_147));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_148, x_148));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_149, x_149));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_150, x_150));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_151, x_151));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_152, x_152));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_153, x_153));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_154, x_154));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_155, x_155));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_156, x_156));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_157, x_157));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_158, x_158));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_159, x_159));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_160, x_160));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_161, x_161));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_162, x_162));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_163, x_163));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_164, x_164));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_165, x_165));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_166, x_166));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_167, x_167));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_168, x_168));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_169, x_169));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_170, x_170));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_171, x_171));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_172, x_172));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_173, x_173));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_174, x_174));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_175, x_175));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_176, x_176));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_177, x_177));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_178, x_178));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_179, x_179));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_180, x_180));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_181, x_181));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_182, x_182));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_183, x_183));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_184, x_184));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_185, x_185));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_186, x_186));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_187, x_187));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_188, x_188));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_189, x_189));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_190, x_190));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_191, x_191));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_192, x_192));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_193, x_193));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_194, x_194));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_195, x_195));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_196, x_196));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_197, x_197));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_198, x_198));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_199, x_199));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_200, x_200));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_201, x_201));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_202, x_202));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_203, x_203));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_204, x_204));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_205, x_205));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_206, x_206));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_207, x_207));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_208, x_208));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_209, x_209));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_210, x_210));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_211, x_211));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_212, x_212));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_213, x_213));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_214, x_214));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_215, x_215));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_216, x_216));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_217, x_217));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_218, x_218));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_219, x_219));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_220, x_220));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_221, x_221));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_222, x_222));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_223, x_223));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_224, x_224));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_225, x_225));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_226, x_226));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_227, x_227));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_228, x_228));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_229, x_229));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_230, x_230));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_231, x_231));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_232, x_232));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_233, x_233));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_234, x_234));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_235, x_235));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_236, x_236));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_237, x_237));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_238, x_238));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_239, x_239));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_240, x_240));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_241, x_241));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_242, x_242));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_243, x_243));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_244, x_244));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_245, x_245));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_246, x_246));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_247, x_247));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_248, x_248));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_249, x_249));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_250, x_250));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_251, x_251));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_252, x_252));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_253, x_253));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_254, x_254));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_ir_6_255, x_255));
        r_sum[6] = sat_add(r_sum[6], b_hr_6);
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_hr_6_0, h_0));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_hr_6_1, h_1));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_hr_6_2, h_2));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_hr_6_3, h_3));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_hr_6_4, h_4));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_hr_6_5, h_5));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_hr_6_6, h_6));
        r_sum[6] = sat_add(r_sum[6], fx_mult_round(w_hr_6_7, h_7));

        // r_sum[7]
        r_sum[7] = b_ir_7;
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_0, x_0));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_1, x_1));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_2, x_2));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_3, x_3));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_4, x_4));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_5, x_5));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_6, x_6));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_7, x_7));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_8, x_8));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_9, x_9));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_10, x_10));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_11, x_11));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_12, x_12));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_13, x_13));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_14, x_14));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_15, x_15));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_16, x_16));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_17, x_17));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_18, x_18));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_19, x_19));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_20, x_20));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_21, x_21));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_22, x_22));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_23, x_23));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_24, x_24));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_25, x_25));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_26, x_26));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_27, x_27));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_28, x_28));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_29, x_29));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_30, x_30));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_31, x_31));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_32, x_32));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_33, x_33));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_34, x_34));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_35, x_35));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_36, x_36));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_37, x_37));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_38, x_38));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_39, x_39));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_40, x_40));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_41, x_41));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_42, x_42));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_43, x_43));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_44, x_44));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_45, x_45));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_46, x_46));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_47, x_47));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_48, x_48));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_49, x_49));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_50, x_50));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_51, x_51));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_52, x_52));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_53, x_53));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_54, x_54));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_55, x_55));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_56, x_56));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_57, x_57));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_58, x_58));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_59, x_59));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_60, x_60));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_61, x_61));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_62, x_62));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_63, x_63));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_64, x_64));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_65, x_65));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_66, x_66));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_67, x_67));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_68, x_68));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_69, x_69));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_70, x_70));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_71, x_71));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_72, x_72));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_73, x_73));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_74, x_74));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_75, x_75));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_76, x_76));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_77, x_77));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_78, x_78));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_79, x_79));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_80, x_80));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_81, x_81));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_82, x_82));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_83, x_83));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_84, x_84));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_85, x_85));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_86, x_86));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_87, x_87));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_88, x_88));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_89, x_89));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_90, x_90));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_91, x_91));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_92, x_92));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_93, x_93));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_94, x_94));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_95, x_95));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_96, x_96));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_97, x_97));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_98, x_98));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_99, x_99));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_100, x_100));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_101, x_101));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_102, x_102));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_103, x_103));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_104, x_104));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_105, x_105));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_106, x_106));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_107, x_107));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_108, x_108));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_109, x_109));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_110, x_110));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_111, x_111));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_112, x_112));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_113, x_113));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_114, x_114));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_115, x_115));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_116, x_116));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_117, x_117));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_118, x_118));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_119, x_119));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_120, x_120));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_121, x_121));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_122, x_122));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_123, x_123));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_124, x_124));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_125, x_125));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_126, x_126));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_127, x_127));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_128, x_128));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_129, x_129));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_130, x_130));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_131, x_131));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_132, x_132));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_133, x_133));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_134, x_134));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_135, x_135));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_136, x_136));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_137, x_137));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_138, x_138));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_139, x_139));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_140, x_140));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_141, x_141));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_142, x_142));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_143, x_143));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_144, x_144));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_145, x_145));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_146, x_146));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_147, x_147));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_148, x_148));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_149, x_149));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_150, x_150));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_151, x_151));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_152, x_152));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_153, x_153));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_154, x_154));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_155, x_155));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_156, x_156));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_157, x_157));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_158, x_158));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_159, x_159));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_160, x_160));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_161, x_161));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_162, x_162));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_163, x_163));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_164, x_164));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_165, x_165));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_166, x_166));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_167, x_167));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_168, x_168));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_169, x_169));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_170, x_170));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_171, x_171));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_172, x_172));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_173, x_173));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_174, x_174));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_175, x_175));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_176, x_176));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_177, x_177));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_178, x_178));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_179, x_179));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_180, x_180));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_181, x_181));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_182, x_182));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_183, x_183));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_184, x_184));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_185, x_185));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_186, x_186));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_187, x_187));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_188, x_188));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_189, x_189));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_190, x_190));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_191, x_191));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_192, x_192));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_193, x_193));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_194, x_194));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_195, x_195));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_196, x_196));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_197, x_197));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_198, x_198));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_199, x_199));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_200, x_200));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_201, x_201));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_202, x_202));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_203, x_203));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_204, x_204));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_205, x_205));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_206, x_206));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_207, x_207));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_208, x_208));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_209, x_209));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_210, x_210));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_211, x_211));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_212, x_212));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_213, x_213));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_214, x_214));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_215, x_215));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_216, x_216));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_217, x_217));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_218, x_218));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_219, x_219));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_220, x_220));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_221, x_221));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_222, x_222));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_223, x_223));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_224, x_224));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_225, x_225));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_226, x_226));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_227, x_227));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_228, x_228));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_229, x_229));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_230, x_230));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_231, x_231));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_232, x_232));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_233, x_233));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_234, x_234));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_235, x_235));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_236, x_236));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_237, x_237));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_238, x_238));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_239, x_239));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_240, x_240));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_241, x_241));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_242, x_242));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_243, x_243));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_244, x_244));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_245, x_245));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_246, x_246));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_247, x_247));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_248, x_248));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_249, x_249));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_250, x_250));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_251, x_251));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_252, x_252));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_253, x_253));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_254, x_254));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_ir_7_255, x_255));
        r_sum[7] = sat_add(r_sum[7], b_hr_7);
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_hr_7_0, h_0));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_hr_7_1, h_1));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_hr_7_2, h_2));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_hr_7_3, h_3));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_hr_7_4, h_4));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_hr_7_5, h_5));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_hr_7_6, h_6));
        r_sum[7] = sat_add(r_sum[7], fx_mult_round(w_hr_7_7, h_7));

    end

    sigmoid #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) sigmoid_r0 (
        .reset(reset), .x(r_sum[0]), .y(r_act[0])
    );
    sigmoid #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) sigmoid_r1 (
        .reset(reset), .x(r_sum[1]), .y(r_act[1])
    );
    sigmoid #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) sigmoid_r2 (
        .reset(reset), .x(r_sum[2]), .y(r_act[2])
    );
    sigmoid #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) sigmoid_r3 (
        .reset(reset), .x(r_sum[3]), .y(r_act[3])
    );
    sigmoid #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) sigmoid_r4 (
        .reset(reset), .x(r_sum[4]), .y(r_act[4])
    );
    sigmoid #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) sigmoid_r5 (
        .reset(reset), .x(r_sum[5]), .y(r_act[5])
    );
    sigmoid #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) sigmoid_r6 (
        .reset(reset), .x(r_sum[6]), .y(r_act[6])
    );
    sigmoid #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) sigmoid_r7 (
        .reset(reset), .x(r_sum[7]), .y(r_act[7])
    );

    // Update gate: z_t = σ(W_iz*x + b_iz + W_hz*h + b_hz)
    // z gate computation
    logic signed [WIDTH-1:0] z_sum[8];
    logic signed [WIDTH-1:0] z_act[8];

    always_comb begin
        // z_sum[0]
        z_sum[0] = b_iz_0;
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_0, x_0));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_1, x_1));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_2, x_2));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_3, x_3));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_4, x_4));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_5, x_5));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_6, x_6));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_7, x_7));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_8, x_8));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_9, x_9));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_10, x_10));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_11, x_11));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_12, x_12));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_13, x_13));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_14, x_14));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_15, x_15));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_16, x_16));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_17, x_17));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_18, x_18));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_19, x_19));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_20, x_20));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_21, x_21));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_22, x_22));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_23, x_23));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_24, x_24));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_25, x_25));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_26, x_26));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_27, x_27));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_28, x_28));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_29, x_29));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_30, x_30));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_31, x_31));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_32, x_32));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_33, x_33));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_34, x_34));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_35, x_35));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_36, x_36));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_37, x_37));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_38, x_38));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_39, x_39));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_40, x_40));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_41, x_41));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_42, x_42));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_43, x_43));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_44, x_44));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_45, x_45));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_46, x_46));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_47, x_47));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_48, x_48));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_49, x_49));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_50, x_50));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_51, x_51));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_52, x_52));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_53, x_53));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_54, x_54));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_55, x_55));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_56, x_56));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_57, x_57));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_58, x_58));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_59, x_59));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_60, x_60));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_61, x_61));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_62, x_62));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_63, x_63));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_64, x_64));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_65, x_65));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_66, x_66));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_67, x_67));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_68, x_68));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_69, x_69));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_70, x_70));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_71, x_71));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_72, x_72));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_73, x_73));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_74, x_74));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_75, x_75));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_76, x_76));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_77, x_77));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_78, x_78));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_79, x_79));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_80, x_80));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_81, x_81));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_82, x_82));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_83, x_83));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_84, x_84));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_85, x_85));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_86, x_86));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_87, x_87));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_88, x_88));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_89, x_89));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_90, x_90));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_91, x_91));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_92, x_92));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_93, x_93));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_94, x_94));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_95, x_95));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_96, x_96));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_97, x_97));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_98, x_98));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_99, x_99));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_100, x_100));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_101, x_101));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_102, x_102));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_103, x_103));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_104, x_104));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_105, x_105));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_106, x_106));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_107, x_107));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_108, x_108));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_109, x_109));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_110, x_110));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_111, x_111));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_112, x_112));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_113, x_113));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_114, x_114));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_115, x_115));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_116, x_116));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_117, x_117));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_118, x_118));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_119, x_119));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_120, x_120));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_121, x_121));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_122, x_122));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_123, x_123));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_124, x_124));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_125, x_125));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_126, x_126));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_127, x_127));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_128, x_128));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_129, x_129));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_130, x_130));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_131, x_131));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_132, x_132));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_133, x_133));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_134, x_134));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_135, x_135));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_136, x_136));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_137, x_137));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_138, x_138));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_139, x_139));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_140, x_140));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_141, x_141));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_142, x_142));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_143, x_143));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_144, x_144));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_145, x_145));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_146, x_146));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_147, x_147));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_148, x_148));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_149, x_149));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_150, x_150));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_151, x_151));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_152, x_152));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_153, x_153));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_154, x_154));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_155, x_155));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_156, x_156));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_157, x_157));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_158, x_158));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_159, x_159));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_160, x_160));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_161, x_161));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_162, x_162));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_163, x_163));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_164, x_164));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_165, x_165));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_166, x_166));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_167, x_167));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_168, x_168));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_169, x_169));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_170, x_170));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_171, x_171));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_172, x_172));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_173, x_173));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_174, x_174));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_175, x_175));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_176, x_176));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_177, x_177));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_178, x_178));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_179, x_179));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_180, x_180));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_181, x_181));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_182, x_182));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_183, x_183));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_184, x_184));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_185, x_185));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_186, x_186));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_187, x_187));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_188, x_188));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_189, x_189));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_190, x_190));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_191, x_191));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_192, x_192));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_193, x_193));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_194, x_194));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_195, x_195));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_196, x_196));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_197, x_197));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_198, x_198));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_199, x_199));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_200, x_200));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_201, x_201));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_202, x_202));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_203, x_203));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_204, x_204));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_205, x_205));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_206, x_206));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_207, x_207));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_208, x_208));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_209, x_209));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_210, x_210));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_211, x_211));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_212, x_212));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_213, x_213));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_214, x_214));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_215, x_215));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_216, x_216));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_217, x_217));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_218, x_218));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_219, x_219));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_220, x_220));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_221, x_221));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_222, x_222));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_223, x_223));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_224, x_224));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_225, x_225));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_226, x_226));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_227, x_227));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_228, x_228));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_229, x_229));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_230, x_230));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_231, x_231));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_232, x_232));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_233, x_233));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_234, x_234));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_235, x_235));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_236, x_236));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_237, x_237));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_238, x_238));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_239, x_239));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_240, x_240));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_241, x_241));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_242, x_242));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_243, x_243));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_244, x_244));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_245, x_245));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_246, x_246));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_247, x_247));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_248, x_248));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_249, x_249));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_250, x_250));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_251, x_251));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_252, x_252));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_253, x_253));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_254, x_254));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_iz_0_255, x_255));
        z_sum[0] = sat_add(z_sum[0], b_hz_0);
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_hz_0_0, h_0));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_hz_0_1, h_1));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_hz_0_2, h_2));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_hz_0_3, h_3));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_hz_0_4, h_4));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_hz_0_5, h_5));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_hz_0_6, h_6));
        z_sum[0] = sat_add(z_sum[0], fx_mult_round(w_hz_0_7, h_7));

        // z_sum[1]
        z_sum[1] = b_iz_1;
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_0, x_0));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_1, x_1));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_2, x_2));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_3, x_3));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_4, x_4));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_5, x_5));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_6, x_6));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_7, x_7));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_8, x_8));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_9, x_9));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_10, x_10));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_11, x_11));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_12, x_12));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_13, x_13));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_14, x_14));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_15, x_15));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_16, x_16));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_17, x_17));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_18, x_18));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_19, x_19));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_20, x_20));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_21, x_21));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_22, x_22));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_23, x_23));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_24, x_24));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_25, x_25));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_26, x_26));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_27, x_27));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_28, x_28));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_29, x_29));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_30, x_30));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_31, x_31));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_32, x_32));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_33, x_33));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_34, x_34));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_35, x_35));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_36, x_36));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_37, x_37));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_38, x_38));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_39, x_39));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_40, x_40));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_41, x_41));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_42, x_42));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_43, x_43));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_44, x_44));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_45, x_45));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_46, x_46));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_47, x_47));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_48, x_48));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_49, x_49));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_50, x_50));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_51, x_51));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_52, x_52));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_53, x_53));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_54, x_54));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_55, x_55));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_56, x_56));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_57, x_57));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_58, x_58));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_59, x_59));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_60, x_60));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_61, x_61));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_62, x_62));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_63, x_63));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_64, x_64));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_65, x_65));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_66, x_66));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_67, x_67));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_68, x_68));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_69, x_69));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_70, x_70));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_71, x_71));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_72, x_72));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_73, x_73));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_74, x_74));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_75, x_75));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_76, x_76));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_77, x_77));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_78, x_78));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_79, x_79));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_80, x_80));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_81, x_81));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_82, x_82));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_83, x_83));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_84, x_84));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_85, x_85));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_86, x_86));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_87, x_87));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_88, x_88));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_89, x_89));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_90, x_90));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_91, x_91));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_92, x_92));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_93, x_93));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_94, x_94));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_95, x_95));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_96, x_96));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_97, x_97));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_98, x_98));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_99, x_99));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_100, x_100));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_101, x_101));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_102, x_102));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_103, x_103));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_104, x_104));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_105, x_105));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_106, x_106));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_107, x_107));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_108, x_108));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_109, x_109));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_110, x_110));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_111, x_111));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_112, x_112));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_113, x_113));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_114, x_114));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_115, x_115));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_116, x_116));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_117, x_117));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_118, x_118));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_119, x_119));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_120, x_120));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_121, x_121));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_122, x_122));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_123, x_123));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_124, x_124));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_125, x_125));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_126, x_126));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_127, x_127));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_128, x_128));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_129, x_129));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_130, x_130));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_131, x_131));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_132, x_132));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_133, x_133));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_134, x_134));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_135, x_135));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_136, x_136));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_137, x_137));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_138, x_138));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_139, x_139));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_140, x_140));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_141, x_141));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_142, x_142));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_143, x_143));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_144, x_144));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_145, x_145));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_146, x_146));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_147, x_147));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_148, x_148));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_149, x_149));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_150, x_150));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_151, x_151));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_152, x_152));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_153, x_153));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_154, x_154));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_155, x_155));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_156, x_156));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_157, x_157));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_158, x_158));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_159, x_159));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_160, x_160));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_161, x_161));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_162, x_162));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_163, x_163));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_164, x_164));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_165, x_165));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_166, x_166));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_167, x_167));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_168, x_168));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_169, x_169));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_170, x_170));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_171, x_171));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_172, x_172));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_173, x_173));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_174, x_174));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_175, x_175));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_176, x_176));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_177, x_177));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_178, x_178));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_179, x_179));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_180, x_180));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_181, x_181));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_182, x_182));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_183, x_183));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_184, x_184));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_185, x_185));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_186, x_186));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_187, x_187));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_188, x_188));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_189, x_189));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_190, x_190));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_191, x_191));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_192, x_192));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_193, x_193));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_194, x_194));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_195, x_195));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_196, x_196));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_197, x_197));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_198, x_198));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_199, x_199));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_200, x_200));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_201, x_201));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_202, x_202));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_203, x_203));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_204, x_204));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_205, x_205));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_206, x_206));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_207, x_207));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_208, x_208));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_209, x_209));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_210, x_210));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_211, x_211));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_212, x_212));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_213, x_213));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_214, x_214));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_215, x_215));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_216, x_216));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_217, x_217));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_218, x_218));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_219, x_219));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_220, x_220));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_221, x_221));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_222, x_222));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_223, x_223));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_224, x_224));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_225, x_225));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_226, x_226));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_227, x_227));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_228, x_228));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_229, x_229));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_230, x_230));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_231, x_231));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_232, x_232));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_233, x_233));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_234, x_234));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_235, x_235));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_236, x_236));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_237, x_237));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_238, x_238));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_239, x_239));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_240, x_240));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_241, x_241));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_242, x_242));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_243, x_243));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_244, x_244));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_245, x_245));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_246, x_246));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_247, x_247));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_248, x_248));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_249, x_249));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_250, x_250));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_251, x_251));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_252, x_252));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_253, x_253));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_254, x_254));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_iz_1_255, x_255));
        z_sum[1] = sat_add(z_sum[1], b_hz_1);
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_hz_1_0, h_0));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_hz_1_1, h_1));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_hz_1_2, h_2));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_hz_1_3, h_3));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_hz_1_4, h_4));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_hz_1_5, h_5));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_hz_1_6, h_6));
        z_sum[1] = sat_add(z_sum[1], fx_mult_round(w_hz_1_7, h_7));

        // z_sum[2]
        z_sum[2] = b_iz_2;
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_0, x_0));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_1, x_1));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_2, x_2));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_3, x_3));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_4, x_4));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_5, x_5));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_6, x_6));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_7, x_7));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_8, x_8));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_9, x_9));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_10, x_10));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_11, x_11));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_12, x_12));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_13, x_13));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_14, x_14));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_15, x_15));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_16, x_16));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_17, x_17));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_18, x_18));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_19, x_19));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_20, x_20));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_21, x_21));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_22, x_22));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_23, x_23));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_24, x_24));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_25, x_25));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_26, x_26));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_27, x_27));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_28, x_28));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_29, x_29));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_30, x_30));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_31, x_31));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_32, x_32));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_33, x_33));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_34, x_34));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_35, x_35));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_36, x_36));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_37, x_37));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_38, x_38));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_39, x_39));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_40, x_40));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_41, x_41));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_42, x_42));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_43, x_43));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_44, x_44));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_45, x_45));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_46, x_46));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_47, x_47));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_48, x_48));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_49, x_49));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_50, x_50));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_51, x_51));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_52, x_52));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_53, x_53));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_54, x_54));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_55, x_55));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_56, x_56));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_57, x_57));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_58, x_58));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_59, x_59));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_60, x_60));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_61, x_61));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_62, x_62));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_63, x_63));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_64, x_64));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_65, x_65));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_66, x_66));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_67, x_67));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_68, x_68));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_69, x_69));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_70, x_70));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_71, x_71));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_72, x_72));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_73, x_73));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_74, x_74));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_75, x_75));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_76, x_76));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_77, x_77));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_78, x_78));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_79, x_79));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_80, x_80));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_81, x_81));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_82, x_82));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_83, x_83));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_84, x_84));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_85, x_85));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_86, x_86));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_87, x_87));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_88, x_88));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_89, x_89));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_90, x_90));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_91, x_91));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_92, x_92));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_93, x_93));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_94, x_94));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_95, x_95));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_96, x_96));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_97, x_97));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_98, x_98));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_99, x_99));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_100, x_100));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_101, x_101));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_102, x_102));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_103, x_103));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_104, x_104));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_105, x_105));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_106, x_106));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_107, x_107));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_108, x_108));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_109, x_109));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_110, x_110));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_111, x_111));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_112, x_112));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_113, x_113));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_114, x_114));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_115, x_115));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_116, x_116));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_117, x_117));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_118, x_118));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_119, x_119));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_120, x_120));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_121, x_121));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_122, x_122));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_123, x_123));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_124, x_124));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_125, x_125));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_126, x_126));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_127, x_127));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_128, x_128));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_129, x_129));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_130, x_130));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_131, x_131));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_132, x_132));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_133, x_133));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_134, x_134));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_135, x_135));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_136, x_136));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_137, x_137));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_138, x_138));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_139, x_139));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_140, x_140));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_141, x_141));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_142, x_142));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_143, x_143));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_144, x_144));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_145, x_145));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_146, x_146));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_147, x_147));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_148, x_148));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_149, x_149));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_150, x_150));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_151, x_151));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_152, x_152));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_153, x_153));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_154, x_154));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_155, x_155));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_156, x_156));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_157, x_157));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_158, x_158));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_159, x_159));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_160, x_160));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_161, x_161));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_162, x_162));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_163, x_163));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_164, x_164));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_165, x_165));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_166, x_166));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_167, x_167));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_168, x_168));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_169, x_169));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_170, x_170));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_171, x_171));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_172, x_172));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_173, x_173));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_174, x_174));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_175, x_175));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_176, x_176));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_177, x_177));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_178, x_178));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_179, x_179));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_180, x_180));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_181, x_181));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_182, x_182));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_183, x_183));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_184, x_184));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_185, x_185));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_186, x_186));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_187, x_187));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_188, x_188));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_189, x_189));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_190, x_190));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_191, x_191));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_192, x_192));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_193, x_193));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_194, x_194));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_195, x_195));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_196, x_196));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_197, x_197));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_198, x_198));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_199, x_199));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_200, x_200));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_201, x_201));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_202, x_202));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_203, x_203));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_204, x_204));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_205, x_205));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_206, x_206));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_207, x_207));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_208, x_208));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_209, x_209));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_210, x_210));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_211, x_211));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_212, x_212));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_213, x_213));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_214, x_214));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_215, x_215));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_216, x_216));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_217, x_217));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_218, x_218));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_219, x_219));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_220, x_220));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_221, x_221));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_222, x_222));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_223, x_223));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_224, x_224));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_225, x_225));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_226, x_226));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_227, x_227));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_228, x_228));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_229, x_229));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_230, x_230));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_231, x_231));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_232, x_232));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_233, x_233));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_234, x_234));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_235, x_235));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_236, x_236));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_237, x_237));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_238, x_238));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_239, x_239));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_240, x_240));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_241, x_241));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_242, x_242));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_243, x_243));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_244, x_244));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_245, x_245));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_246, x_246));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_247, x_247));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_248, x_248));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_249, x_249));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_250, x_250));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_251, x_251));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_252, x_252));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_253, x_253));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_254, x_254));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_iz_2_255, x_255));
        z_sum[2] = sat_add(z_sum[2], b_hz_2);
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_hz_2_0, h_0));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_hz_2_1, h_1));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_hz_2_2, h_2));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_hz_2_3, h_3));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_hz_2_4, h_4));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_hz_2_5, h_5));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_hz_2_6, h_6));
        z_sum[2] = sat_add(z_sum[2], fx_mult_round(w_hz_2_7, h_7));

        // z_sum[3]
        z_sum[3] = b_iz_3;
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_0, x_0));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_1, x_1));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_2, x_2));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_3, x_3));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_4, x_4));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_5, x_5));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_6, x_6));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_7, x_7));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_8, x_8));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_9, x_9));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_10, x_10));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_11, x_11));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_12, x_12));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_13, x_13));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_14, x_14));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_15, x_15));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_16, x_16));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_17, x_17));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_18, x_18));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_19, x_19));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_20, x_20));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_21, x_21));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_22, x_22));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_23, x_23));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_24, x_24));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_25, x_25));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_26, x_26));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_27, x_27));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_28, x_28));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_29, x_29));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_30, x_30));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_31, x_31));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_32, x_32));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_33, x_33));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_34, x_34));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_35, x_35));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_36, x_36));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_37, x_37));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_38, x_38));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_39, x_39));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_40, x_40));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_41, x_41));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_42, x_42));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_43, x_43));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_44, x_44));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_45, x_45));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_46, x_46));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_47, x_47));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_48, x_48));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_49, x_49));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_50, x_50));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_51, x_51));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_52, x_52));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_53, x_53));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_54, x_54));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_55, x_55));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_56, x_56));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_57, x_57));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_58, x_58));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_59, x_59));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_60, x_60));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_61, x_61));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_62, x_62));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_63, x_63));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_64, x_64));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_65, x_65));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_66, x_66));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_67, x_67));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_68, x_68));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_69, x_69));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_70, x_70));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_71, x_71));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_72, x_72));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_73, x_73));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_74, x_74));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_75, x_75));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_76, x_76));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_77, x_77));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_78, x_78));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_79, x_79));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_80, x_80));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_81, x_81));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_82, x_82));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_83, x_83));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_84, x_84));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_85, x_85));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_86, x_86));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_87, x_87));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_88, x_88));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_89, x_89));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_90, x_90));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_91, x_91));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_92, x_92));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_93, x_93));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_94, x_94));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_95, x_95));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_96, x_96));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_97, x_97));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_98, x_98));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_99, x_99));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_100, x_100));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_101, x_101));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_102, x_102));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_103, x_103));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_104, x_104));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_105, x_105));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_106, x_106));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_107, x_107));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_108, x_108));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_109, x_109));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_110, x_110));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_111, x_111));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_112, x_112));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_113, x_113));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_114, x_114));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_115, x_115));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_116, x_116));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_117, x_117));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_118, x_118));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_119, x_119));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_120, x_120));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_121, x_121));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_122, x_122));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_123, x_123));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_124, x_124));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_125, x_125));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_126, x_126));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_127, x_127));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_128, x_128));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_129, x_129));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_130, x_130));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_131, x_131));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_132, x_132));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_133, x_133));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_134, x_134));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_135, x_135));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_136, x_136));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_137, x_137));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_138, x_138));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_139, x_139));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_140, x_140));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_141, x_141));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_142, x_142));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_143, x_143));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_144, x_144));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_145, x_145));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_146, x_146));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_147, x_147));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_148, x_148));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_149, x_149));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_150, x_150));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_151, x_151));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_152, x_152));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_153, x_153));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_154, x_154));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_155, x_155));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_156, x_156));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_157, x_157));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_158, x_158));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_159, x_159));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_160, x_160));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_161, x_161));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_162, x_162));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_163, x_163));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_164, x_164));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_165, x_165));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_166, x_166));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_167, x_167));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_168, x_168));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_169, x_169));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_170, x_170));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_171, x_171));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_172, x_172));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_173, x_173));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_174, x_174));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_175, x_175));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_176, x_176));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_177, x_177));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_178, x_178));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_179, x_179));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_180, x_180));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_181, x_181));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_182, x_182));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_183, x_183));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_184, x_184));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_185, x_185));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_186, x_186));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_187, x_187));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_188, x_188));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_189, x_189));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_190, x_190));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_191, x_191));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_192, x_192));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_193, x_193));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_194, x_194));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_195, x_195));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_196, x_196));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_197, x_197));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_198, x_198));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_199, x_199));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_200, x_200));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_201, x_201));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_202, x_202));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_203, x_203));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_204, x_204));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_205, x_205));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_206, x_206));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_207, x_207));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_208, x_208));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_209, x_209));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_210, x_210));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_211, x_211));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_212, x_212));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_213, x_213));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_214, x_214));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_215, x_215));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_216, x_216));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_217, x_217));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_218, x_218));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_219, x_219));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_220, x_220));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_221, x_221));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_222, x_222));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_223, x_223));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_224, x_224));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_225, x_225));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_226, x_226));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_227, x_227));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_228, x_228));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_229, x_229));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_230, x_230));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_231, x_231));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_232, x_232));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_233, x_233));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_234, x_234));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_235, x_235));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_236, x_236));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_237, x_237));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_238, x_238));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_239, x_239));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_240, x_240));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_241, x_241));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_242, x_242));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_243, x_243));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_244, x_244));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_245, x_245));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_246, x_246));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_247, x_247));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_248, x_248));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_249, x_249));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_250, x_250));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_251, x_251));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_252, x_252));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_253, x_253));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_254, x_254));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_iz_3_255, x_255));
        z_sum[3] = sat_add(z_sum[3], b_hz_3);
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_hz_3_0, h_0));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_hz_3_1, h_1));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_hz_3_2, h_2));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_hz_3_3, h_3));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_hz_3_4, h_4));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_hz_3_5, h_5));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_hz_3_6, h_6));
        z_sum[3] = sat_add(z_sum[3], fx_mult_round(w_hz_3_7, h_7));

        // z_sum[4]
        z_sum[4] = b_iz_4;
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_0, x_0));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_1, x_1));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_2, x_2));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_3, x_3));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_4, x_4));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_5, x_5));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_6, x_6));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_7, x_7));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_8, x_8));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_9, x_9));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_10, x_10));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_11, x_11));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_12, x_12));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_13, x_13));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_14, x_14));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_15, x_15));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_16, x_16));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_17, x_17));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_18, x_18));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_19, x_19));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_20, x_20));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_21, x_21));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_22, x_22));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_23, x_23));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_24, x_24));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_25, x_25));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_26, x_26));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_27, x_27));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_28, x_28));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_29, x_29));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_30, x_30));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_31, x_31));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_32, x_32));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_33, x_33));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_34, x_34));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_35, x_35));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_36, x_36));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_37, x_37));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_38, x_38));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_39, x_39));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_40, x_40));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_41, x_41));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_42, x_42));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_43, x_43));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_44, x_44));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_45, x_45));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_46, x_46));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_47, x_47));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_48, x_48));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_49, x_49));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_50, x_50));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_51, x_51));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_52, x_52));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_53, x_53));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_54, x_54));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_55, x_55));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_56, x_56));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_57, x_57));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_58, x_58));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_59, x_59));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_60, x_60));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_61, x_61));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_62, x_62));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_63, x_63));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_64, x_64));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_65, x_65));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_66, x_66));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_67, x_67));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_68, x_68));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_69, x_69));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_70, x_70));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_71, x_71));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_72, x_72));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_73, x_73));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_74, x_74));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_75, x_75));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_76, x_76));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_77, x_77));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_78, x_78));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_79, x_79));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_80, x_80));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_81, x_81));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_82, x_82));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_83, x_83));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_84, x_84));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_85, x_85));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_86, x_86));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_87, x_87));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_88, x_88));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_89, x_89));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_90, x_90));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_91, x_91));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_92, x_92));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_93, x_93));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_94, x_94));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_95, x_95));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_96, x_96));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_97, x_97));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_98, x_98));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_99, x_99));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_100, x_100));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_101, x_101));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_102, x_102));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_103, x_103));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_104, x_104));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_105, x_105));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_106, x_106));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_107, x_107));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_108, x_108));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_109, x_109));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_110, x_110));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_111, x_111));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_112, x_112));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_113, x_113));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_114, x_114));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_115, x_115));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_116, x_116));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_117, x_117));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_118, x_118));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_119, x_119));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_120, x_120));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_121, x_121));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_122, x_122));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_123, x_123));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_124, x_124));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_125, x_125));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_126, x_126));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_127, x_127));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_128, x_128));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_129, x_129));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_130, x_130));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_131, x_131));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_132, x_132));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_133, x_133));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_134, x_134));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_135, x_135));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_136, x_136));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_137, x_137));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_138, x_138));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_139, x_139));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_140, x_140));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_141, x_141));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_142, x_142));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_143, x_143));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_144, x_144));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_145, x_145));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_146, x_146));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_147, x_147));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_148, x_148));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_149, x_149));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_150, x_150));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_151, x_151));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_152, x_152));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_153, x_153));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_154, x_154));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_155, x_155));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_156, x_156));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_157, x_157));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_158, x_158));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_159, x_159));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_160, x_160));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_161, x_161));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_162, x_162));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_163, x_163));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_164, x_164));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_165, x_165));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_166, x_166));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_167, x_167));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_168, x_168));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_169, x_169));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_170, x_170));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_171, x_171));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_172, x_172));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_173, x_173));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_174, x_174));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_175, x_175));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_176, x_176));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_177, x_177));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_178, x_178));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_179, x_179));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_180, x_180));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_181, x_181));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_182, x_182));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_183, x_183));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_184, x_184));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_185, x_185));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_186, x_186));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_187, x_187));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_188, x_188));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_189, x_189));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_190, x_190));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_191, x_191));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_192, x_192));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_193, x_193));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_194, x_194));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_195, x_195));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_196, x_196));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_197, x_197));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_198, x_198));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_199, x_199));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_200, x_200));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_201, x_201));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_202, x_202));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_203, x_203));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_204, x_204));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_205, x_205));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_206, x_206));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_207, x_207));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_208, x_208));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_209, x_209));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_210, x_210));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_211, x_211));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_212, x_212));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_213, x_213));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_214, x_214));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_215, x_215));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_216, x_216));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_217, x_217));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_218, x_218));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_219, x_219));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_220, x_220));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_221, x_221));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_222, x_222));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_223, x_223));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_224, x_224));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_225, x_225));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_226, x_226));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_227, x_227));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_228, x_228));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_229, x_229));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_230, x_230));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_231, x_231));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_232, x_232));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_233, x_233));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_234, x_234));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_235, x_235));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_236, x_236));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_237, x_237));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_238, x_238));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_239, x_239));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_240, x_240));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_241, x_241));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_242, x_242));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_243, x_243));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_244, x_244));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_245, x_245));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_246, x_246));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_247, x_247));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_248, x_248));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_249, x_249));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_250, x_250));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_251, x_251));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_252, x_252));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_253, x_253));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_254, x_254));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_iz_4_255, x_255));
        z_sum[4] = sat_add(z_sum[4], b_hz_4);
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_hz_4_0, h_0));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_hz_4_1, h_1));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_hz_4_2, h_2));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_hz_4_3, h_3));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_hz_4_4, h_4));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_hz_4_5, h_5));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_hz_4_6, h_6));
        z_sum[4] = sat_add(z_sum[4], fx_mult_round(w_hz_4_7, h_7));

        // z_sum[5]
        z_sum[5] = b_iz_5;
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_0, x_0));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_1, x_1));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_2, x_2));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_3, x_3));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_4, x_4));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_5, x_5));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_6, x_6));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_7, x_7));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_8, x_8));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_9, x_9));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_10, x_10));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_11, x_11));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_12, x_12));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_13, x_13));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_14, x_14));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_15, x_15));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_16, x_16));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_17, x_17));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_18, x_18));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_19, x_19));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_20, x_20));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_21, x_21));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_22, x_22));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_23, x_23));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_24, x_24));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_25, x_25));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_26, x_26));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_27, x_27));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_28, x_28));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_29, x_29));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_30, x_30));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_31, x_31));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_32, x_32));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_33, x_33));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_34, x_34));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_35, x_35));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_36, x_36));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_37, x_37));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_38, x_38));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_39, x_39));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_40, x_40));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_41, x_41));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_42, x_42));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_43, x_43));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_44, x_44));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_45, x_45));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_46, x_46));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_47, x_47));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_48, x_48));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_49, x_49));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_50, x_50));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_51, x_51));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_52, x_52));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_53, x_53));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_54, x_54));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_55, x_55));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_56, x_56));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_57, x_57));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_58, x_58));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_59, x_59));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_60, x_60));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_61, x_61));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_62, x_62));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_63, x_63));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_64, x_64));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_65, x_65));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_66, x_66));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_67, x_67));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_68, x_68));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_69, x_69));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_70, x_70));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_71, x_71));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_72, x_72));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_73, x_73));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_74, x_74));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_75, x_75));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_76, x_76));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_77, x_77));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_78, x_78));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_79, x_79));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_80, x_80));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_81, x_81));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_82, x_82));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_83, x_83));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_84, x_84));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_85, x_85));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_86, x_86));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_87, x_87));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_88, x_88));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_89, x_89));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_90, x_90));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_91, x_91));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_92, x_92));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_93, x_93));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_94, x_94));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_95, x_95));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_96, x_96));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_97, x_97));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_98, x_98));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_99, x_99));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_100, x_100));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_101, x_101));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_102, x_102));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_103, x_103));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_104, x_104));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_105, x_105));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_106, x_106));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_107, x_107));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_108, x_108));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_109, x_109));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_110, x_110));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_111, x_111));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_112, x_112));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_113, x_113));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_114, x_114));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_115, x_115));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_116, x_116));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_117, x_117));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_118, x_118));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_119, x_119));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_120, x_120));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_121, x_121));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_122, x_122));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_123, x_123));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_124, x_124));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_125, x_125));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_126, x_126));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_127, x_127));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_128, x_128));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_129, x_129));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_130, x_130));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_131, x_131));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_132, x_132));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_133, x_133));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_134, x_134));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_135, x_135));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_136, x_136));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_137, x_137));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_138, x_138));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_139, x_139));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_140, x_140));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_141, x_141));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_142, x_142));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_143, x_143));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_144, x_144));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_145, x_145));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_146, x_146));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_147, x_147));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_148, x_148));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_149, x_149));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_150, x_150));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_151, x_151));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_152, x_152));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_153, x_153));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_154, x_154));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_155, x_155));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_156, x_156));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_157, x_157));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_158, x_158));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_159, x_159));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_160, x_160));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_161, x_161));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_162, x_162));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_163, x_163));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_164, x_164));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_165, x_165));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_166, x_166));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_167, x_167));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_168, x_168));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_169, x_169));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_170, x_170));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_171, x_171));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_172, x_172));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_173, x_173));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_174, x_174));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_175, x_175));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_176, x_176));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_177, x_177));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_178, x_178));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_179, x_179));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_180, x_180));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_181, x_181));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_182, x_182));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_183, x_183));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_184, x_184));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_185, x_185));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_186, x_186));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_187, x_187));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_188, x_188));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_189, x_189));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_190, x_190));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_191, x_191));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_192, x_192));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_193, x_193));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_194, x_194));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_195, x_195));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_196, x_196));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_197, x_197));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_198, x_198));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_199, x_199));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_200, x_200));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_201, x_201));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_202, x_202));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_203, x_203));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_204, x_204));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_205, x_205));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_206, x_206));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_207, x_207));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_208, x_208));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_209, x_209));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_210, x_210));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_211, x_211));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_212, x_212));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_213, x_213));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_214, x_214));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_215, x_215));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_216, x_216));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_217, x_217));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_218, x_218));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_219, x_219));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_220, x_220));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_221, x_221));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_222, x_222));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_223, x_223));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_224, x_224));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_225, x_225));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_226, x_226));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_227, x_227));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_228, x_228));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_229, x_229));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_230, x_230));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_231, x_231));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_232, x_232));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_233, x_233));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_234, x_234));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_235, x_235));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_236, x_236));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_237, x_237));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_238, x_238));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_239, x_239));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_240, x_240));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_241, x_241));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_242, x_242));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_243, x_243));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_244, x_244));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_245, x_245));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_246, x_246));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_247, x_247));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_248, x_248));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_249, x_249));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_250, x_250));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_251, x_251));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_252, x_252));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_253, x_253));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_254, x_254));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_iz_5_255, x_255));
        z_sum[5] = sat_add(z_sum[5], b_hz_5);
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_hz_5_0, h_0));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_hz_5_1, h_1));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_hz_5_2, h_2));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_hz_5_3, h_3));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_hz_5_4, h_4));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_hz_5_5, h_5));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_hz_5_6, h_6));
        z_sum[5] = sat_add(z_sum[5], fx_mult_round(w_hz_5_7, h_7));

        // z_sum[6]
        z_sum[6] = b_iz_6;
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_0, x_0));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_1, x_1));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_2, x_2));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_3, x_3));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_4, x_4));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_5, x_5));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_6, x_6));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_7, x_7));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_8, x_8));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_9, x_9));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_10, x_10));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_11, x_11));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_12, x_12));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_13, x_13));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_14, x_14));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_15, x_15));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_16, x_16));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_17, x_17));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_18, x_18));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_19, x_19));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_20, x_20));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_21, x_21));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_22, x_22));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_23, x_23));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_24, x_24));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_25, x_25));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_26, x_26));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_27, x_27));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_28, x_28));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_29, x_29));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_30, x_30));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_31, x_31));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_32, x_32));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_33, x_33));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_34, x_34));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_35, x_35));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_36, x_36));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_37, x_37));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_38, x_38));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_39, x_39));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_40, x_40));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_41, x_41));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_42, x_42));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_43, x_43));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_44, x_44));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_45, x_45));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_46, x_46));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_47, x_47));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_48, x_48));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_49, x_49));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_50, x_50));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_51, x_51));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_52, x_52));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_53, x_53));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_54, x_54));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_55, x_55));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_56, x_56));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_57, x_57));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_58, x_58));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_59, x_59));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_60, x_60));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_61, x_61));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_62, x_62));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_63, x_63));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_64, x_64));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_65, x_65));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_66, x_66));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_67, x_67));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_68, x_68));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_69, x_69));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_70, x_70));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_71, x_71));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_72, x_72));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_73, x_73));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_74, x_74));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_75, x_75));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_76, x_76));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_77, x_77));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_78, x_78));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_79, x_79));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_80, x_80));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_81, x_81));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_82, x_82));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_83, x_83));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_84, x_84));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_85, x_85));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_86, x_86));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_87, x_87));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_88, x_88));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_89, x_89));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_90, x_90));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_91, x_91));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_92, x_92));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_93, x_93));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_94, x_94));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_95, x_95));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_96, x_96));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_97, x_97));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_98, x_98));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_99, x_99));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_100, x_100));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_101, x_101));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_102, x_102));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_103, x_103));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_104, x_104));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_105, x_105));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_106, x_106));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_107, x_107));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_108, x_108));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_109, x_109));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_110, x_110));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_111, x_111));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_112, x_112));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_113, x_113));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_114, x_114));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_115, x_115));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_116, x_116));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_117, x_117));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_118, x_118));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_119, x_119));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_120, x_120));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_121, x_121));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_122, x_122));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_123, x_123));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_124, x_124));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_125, x_125));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_126, x_126));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_127, x_127));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_128, x_128));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_129, x_129));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_130, x_130));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_131, x_131));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_132, x_132));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_133, x_133));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_134, x_134));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_135, x_135));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_136, x_136));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_137, x_137));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_138, x_138));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_139, x_139));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_140, x_140));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_141, x_141));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_142, x_142));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_143, x_143));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_144, x_144));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_145, x_145));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_146, x_146));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_147, x_147));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_148, x_148));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_149, x_149));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_150, x_150));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_151, x_151));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_152, x_152));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_153, x_153));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_154, x_154));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_155, x_155));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_156, x_156));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_157, x_157));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_158, x_158));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_159, x_159));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_160, x_160));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_161, x_161));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_162, x_162));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_163, x_163));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_164, x_164));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_165, x_165));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_166, x_166));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_167, x_167));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_168, x_168));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_169, x_169));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_170, x_170));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_171, x_171));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_172, x_172));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_173, x_173));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_174, x_174));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_175, x_175));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_176, x_176));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_177, x_177));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_178, x_178));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_179, x_179));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_180, x_180));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_181, x_181));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_182, x_182));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_183, x_183));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_184, x_184));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_185, x_185));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_186, x_186));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_187, x_187));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_188, x_188));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_189, x_189));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_190, x_190));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_191, x_191));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_192, x_192));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_193, x_193));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_194, x_194));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_195, x_195));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_196, x_196));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_197, x_197));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_198, x_198));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_199, x_199));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_200, x_200));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_201, x_201));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_202, x_202));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_203, x_203));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_204, x_204));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_205, x_205));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_206, x_206));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_207, x_207));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_208, x_208));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_209, x_209));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_210, x_210));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_211, x_211));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_212, x_212));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_213, x_213));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_214, x_214));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_215, x_215));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_216, x_216));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_217, x_217));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_218, x_218));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_219, x_219));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_220, x_220));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_221, x_221));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_222, x_222));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_223, x_223));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_224, x_224));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_225, x_225));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_226, x_226));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_227, x_227));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_228, x_228));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_229, x_229));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_230, x_230));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_231, x_231));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_232, x_232));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_233, x_233));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_234, x_234));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_235, x_235));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_236, x_236));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_237, x_237));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_238, x_238));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_239, x_239));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_240, x_240));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_241, x_241));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_242, x_242));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_243, x_243));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_244, x_244));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_245, x_245));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_246, x_246));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_247, x_247));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_248, x_248));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_249, x_249));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_250, x_250));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_251, x_251));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_252, x_252));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_253, x_253));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_254, x_254));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_iz_6_255, x_255));
        z_sum[6] = sat_add(z_sum[6], b_hz_6);
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_hz_6_0, h_0));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_hz_6_1, h_1));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_hz_6_2, h_2));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_hz_6_3, h_3));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_hz_6_4, h_4));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_hz_6_5, h_5));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_hz_6_6, h_6));
        z_sum[6] = sat_add(z_sum[6], fx_mult_round(w_hz_6_7, h_7));

        // z_sum[7]
        z_sum[7] = b_iz_7;
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_0, x_0));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_1, x_1));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_2, x_2));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_3, x_3));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_4, x_4));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_5, x_5));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_6, x_6));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_7, x_7));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_8, x_8));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_9, x_9));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_10, x_10));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_11, x_11));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_12, x_12));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_13, x_13));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_14, x_14));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_15, x_15));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_16, x_16));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_17, x_17));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_18, x_18));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_19, x_19));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_20, x_20));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_21, x_21));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_22, x_22));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_23, x_23));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_24, x_24));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_25, x_25));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_26, x_26));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_27, x_27));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_28, x_28));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_29, x_29));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_30, x_30));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_31, x_31));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_32, x_32));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_33, x_33));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_34, x_34));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_35, x_35));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_36, x_36));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_37, x_37));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_38, x_38));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_39, x_39));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_40, x_40));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_41, x_41));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_42, x_42));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_43, x_43));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_44, x_44));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_45, x_45));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_46, x_46));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_47, x_47));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_48, x_48));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_49, x_49));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_50, x_50));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_51, x_51));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_52, x_52));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_53, x_53));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_54, x_54));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_55, x_55));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_56, x_56));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_57, x_57));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_58, x_58));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_59, x_59));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_60, x_60));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_61, x_61));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_62, x_62));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_63, x_63));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_64, x_64));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_65, x_65));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_66, x_66));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_67, x_67));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_68, x_68));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_69, x_69));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_70, x_70));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_71, x_71));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_72, x_72));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_73, x_73));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_74, x_74));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_75, x_75));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_76, x_76));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_77, x_77));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_78, x_78));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_79, x_79));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_80, x_80));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_81, x_81));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_82, x_82));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_83, x_83));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_84, x_84));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_85, x_85));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_86, x_86));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_87, x_87));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_88, x_88));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_89, x_89));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_90, x_90));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_91, x_91));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_92, x_92));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_93, x_93));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_94, x_94));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_95, x_95));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_96, x_96));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_97, x_97));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_98, x_98));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_99, x_99));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_100, x_100));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_101, x_101));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_102, x_102));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_103, x_103));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_104, x_104));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_105, x_105));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_106, x_106));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_107, x_107));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_108, x_108));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_109, x_109));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_110, x_110));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_111, x_111));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_112, x_112));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_113, x_113));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_114, x_114));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_115, x_115));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_116, x_116));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_117, x_117));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_118, x_118));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_119, x_119));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_120, x_120));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_121, x_121));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_122, x_122));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_123, x_123));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_124, x_124));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_125, x_125));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_126, x_126));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_127, x_127));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_128, x_128));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_129, x_129));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_130, x_130));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_131, x_131));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_132, x_132));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_133, x_133));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_134, x_134));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_135, x_135));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_136, x_136));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_137, x_137));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_138, x_138));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_139, x_139));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_140, x_140));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_141, x_141));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_142, x_142));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_143, x_143));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_144, x_144));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_145, x_145));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_146, x_146));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_147, x_147));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_148, x_148));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_149, x_149));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_150, x_150));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_151, x_151));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_152, x_152));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_153, x_153));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_154, x_154));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_155, x_155));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_156, x_156));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_157, x_157));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_158, x_158));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_159, x_159));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_160, x_160));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_161, x_161));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_162, x_162));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_163, x_163));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_164, x_164));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_165, x_165));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_166, x_166));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_167, x_167));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_168, x_168));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_169, x_169));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_170, x_170));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_171, x_171));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_172, x_172));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_173, x_173));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_174, x_174));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_175, x_175));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_176, x_176));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_177, x_177));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_178, x_178));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_179, x_179));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_180, x_180));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_181, x_181));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_182, x_182));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_183, x_183));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_184, x_184));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_185, x_185));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_186, x_186));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_187, x_187));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_188, x_188));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_189, x_189));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_190, x_190));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_191, x_191));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_192, x_192));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_193, x_193));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_194, x_194));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_195, x_195));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_196, x_196));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_197, x_197));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_198, x_198));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_199, x_199));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_200, x_200));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_201, x_201));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_202, x_202));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_203, x_203));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_204, x_204));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_205, x_205));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_206, x_206));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_207, x_207));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_208, x_208));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_209, x_209));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_210, x_210));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_211, x_211));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_212, x_212));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_213, x_213));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_214, x_214));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_215, x_215));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_216, x_216));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_217, x_217));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_218, x_218));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_219, x_219));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_220, x_220));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_221, x_221));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_222, x_222));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_223, x_223));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_224, x_224));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_225, x_225));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_226, x_226));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_227, x_227));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_228, x_228));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_229, x_229));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_230, x_230));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_231, x_231));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_232, x_232));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_233, x_233));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_234, x_234));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_235, x_235));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_236, x_236));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_237, x_237));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_238, x_238));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_239, x_239));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_240, x_240));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_241, x_241));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_242, x_242));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_243, x_243));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_244, x_244));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_245, x_245));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_246, x_246));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_247, x_247));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_248, x_248));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_249, x_249));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_250, x_250));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_251, x_251));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_252, x_252));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_253, x_253));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_254, x_254));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_iz_7_255, x_255));
        z_sum[7] = sat_add(z_sum[7], b_hz_7);
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_hz_7_0, h_0));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_hz_7_1, h_1));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_hz_7_2, h_2));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_hz_7_3, h_3));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_hz_7_4, h_4));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_hz_7_5, h_5));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_hz_7_6, h_6));
        z_sum[7] = sat_add(z_sum[7], fx_mult_round(w_hz_7_7, h_7));

    end

    sigmoid #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) sigmoid_z0 (
        .reset(reset), .x(z_sum[0]), .y(z_act[0])
    );
    sigmoid #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) sigmoid_z1 (
        .reset(reset), .x(z_sum[1]), .y(z_act[1])
    );
    sigmoid #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) sigmoid_z2 (
        .reset(reset), .x(z_sum[2]), .y(z_act[2])
    );
    sigmoid #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) sigmoid_z3 (
        .reset(reset), .x(z_sum[3]), .y(z_act[3])
    );
    sigmoid #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) sigmoid_z4 (
        .reset(reset), .x(z_sum[4]), .y(z_act[4])
    );
    sigmoid #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) sigmoid_z5 (
        .reset(reset), .x(z_sum[5]), .y(z_act[5])
    );
    sigmoid #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) sigmoid_z6 (
        .reset(reset), .x(z_sum[6]), .y(z_act[6])
    );
    sigmoid #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) sigmoid_z7 (
        .reset(reset), .x(z_sum[7]), .y(z_act[7])
    );

    // Candidate hidden state: n_t = tanh(W_in*x + b_in + r_t ⊙ (W_hn*h + b_hn))
    // Candidate hidden state computation
    logic signed [WIDTH-1:0] wn_h[8];
    logic signed [WIDTH-1:0] gated_h[8];
    logic signed [WIDTH-1:0] n_sum[8];
    logic signed [WIDTH-1:0] n_act[8];

    always_comb begin
        // wn_h[0] = W_hn*h + b_hn
        wn_h[0] = b_hn_0;
        wn_h[0] = sat_add(wn_h[0], fx_mult_round(w_hn_0_0, h_0));
        wn_h[0] = sat_add(wn_h[0], fx_mult_round(w_hn_0_1, h_1));
        wn_h[0] = sat_add(wn_h[0], fx_mult_round(w_hn_0_2, h_2));
        wn_h[0] = sat_add(wn_h[0], fx_mult_round(w_hn_0_3, h_3));
        wn_h[0] = sat_add(wn_h[0], fx_mult_round(w_hn_0_4, h_4));
        wn_h[0] = sat_add(wn_h[0], fx_mult_round(w_hn_0_5, h_5));
        wn_h[0] = sat_add(wn_h[0], fx_mult_round(w_hn_0_6, h_6));
        wn_h[0] = sat_add(wn_h[0], fx_mult_round(w_hn_0_7, h_7));

        // gated_h[0] = r_t ⊙ wn_h
        gated_h[0] = fx_mult_round(r_act[0], wn_h[0]);

        // n_sum[0] = W_in*x + b_in + gated_h
        n_sum[0] = b_in_0;
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_0, x_0));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_1, x_1));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_2, x_2));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_3, x_3));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_4, x_4));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_5, x_5));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_6, x_6));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_7, x_7));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_8, x_8));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_9, x_9));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_10, x_10));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_11, x_11));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_12, x_12));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_13, x_13));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_14, x_14));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_15, x_15));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_16, x_16));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_17, x_17));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_18, x_18));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_19, x_19));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_20, x_20));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_21, x_21));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_22, x_22));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_23, x_23));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_24, x_24));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_25, x_25));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_26, x_26));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_27, x_27));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_28, x_28));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_29, x_29));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_30, x_30));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_31, x_31));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_32, x_32));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_33, x_33));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_34, x_34));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_35, x_35));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_36, x_36));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_37, x_37));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_38, x_38));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_39, x_39));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_40, x_40));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_41, x_41));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_42, x_42));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_43, x_43));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_44, x_44));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_45, x_45));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_46, x_46));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_47, x_47));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_48, x_48));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_49, x_49));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_50, x_50));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_51, x_51));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_52, x_52));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_53, x_53));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_54, x_54));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_55, x_55));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_56, x_56));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_57, x_57));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_58, x_58));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_59, x_59));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_60, x_60));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_61, x_61));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_62, x_62));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_63, x_63));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_64, x_64));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_65, x_65));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_66, x_66));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_67, x_67));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_68, x_68));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_69, x_69));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_70, x_70));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_71, x_71));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_72, x_72));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_73, x_73));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_74, x_74));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_75, x_75));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_76, x_76));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_77, x_77));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_78, x_78));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_79, x_79));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_80, x_80));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_81, x_81));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_82, x_82));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_83, x_83));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_84, x_84));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_85, x_85));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_86, x_86));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_87, x_87));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_88, x_88));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_89, x_89));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_90, x_90));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_91, x_91));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_92, x_92));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_93, x_93));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_94, x_94));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_95, x_95));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_96, x_96));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_97, x_97));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_98, x_98));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_99, x_99));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_100, x_100));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_101, x_101));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_102, x_102));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_103, x_103));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_104, x_104));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_105, x_105));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_106, x_106));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_107, x_107));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_108, x_108));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_109, x_109));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_110, x_110));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_111, x_111));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_112, x_112));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_113, x_113));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_114, x_114));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_115, x_115));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_116, x_116));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_117, x_117));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_118, x_118));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_119, x_119));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_120, x_120));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_121, x_121));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_122, x_122));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_123, x_123));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_124, x_124));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_125, x_125));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_126, x_126));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_127, x_127));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_128, x_128));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_129, x_129));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_130, x_130));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_131, x_131));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_132, x_132));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_133, x_133));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_134, x_134));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_135, x_135));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_136, x_136));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_137, x_137));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_138, x_138));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_139, x_139));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_140, x_140));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_141, x_141));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_142, x_142));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_143, x_143));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_144, x_144));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_145, x_145));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_146, x_146));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_147, x_147));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_148, x_148));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_149, x_149));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_150, x_150));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_151, x_151));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_152, x_152));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_153, x_153));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_154, x_154));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_155, x_155));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_156, x_156));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_157, x_157));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_158, x_158));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_159, x_159));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_160, x_160));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_161, x_161));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_162, x_162));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_163, x_163));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_164, x_164));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_165, x_165));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_166, x_166));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_167, x_167));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_168, x_168));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_169, x_169));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_170, x_170));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_171, x_171));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_172, x_172));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_173, x_173));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_174, x_174));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_175, x_175));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_176, x_176));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_177, x_177));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_178, x_178));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_179, x_179));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_180, x_180));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_181, x_181));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_182, x_182));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_183, x_183));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_184, x_184));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_185, x_185));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_186, x_186));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_187, x_187));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_188, x_188));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_189, x_189));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_190, x_190));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_191, x_191));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_192, x_192));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_193, x_193));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_194, x_194));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_195, x_195));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_196, x_196));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_197, x_197));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_198, x_198));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_199, x_199));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_200, x_200));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_201, x_201));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_202, x_202));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_203, x_203));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_204, x_204));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_205, x_205));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_206, x_206));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_207, x_207));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_208, x_208));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_209, x_209));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_210, x_210));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_211, x_211));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_212, x_212));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_213, x_213));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_214, x_214));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_215, x_215));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_216, x_216));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_217, x_217));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_218, x_218));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_219, x_219));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_220, x_220));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_221, x_221));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_222, x_222));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_223, x_223));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_224, x_224));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_225, x_225));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_226, x_226));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_227, x_227));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_228, x_228));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_229, x_229));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_230, x_230));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_231, x_231));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_232, x_232));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_233, x_233));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_234, x_234));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_235, x_235));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_236, x_236));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_237, x_237));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_238, x_238));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_239, x_239));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_240, x_240));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_241, x_241));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_242, x_242));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_243, x_243));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_244, x_244));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_245, x_245));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_246, x_246));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_247, x_247));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_248, x_248));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_249, x_249));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_250, x_250));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_251, x_251));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_252, x_252));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_253, x_253));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_254, x_254));
        n_sum[0] = sat_add(n_sum[0], fx_mult_round(w_in_0_255, x_255));
        n_sum[0] = sat_add(n_sum[0], gated_h[0]);

        // wn_h[1] = W_hn*h + b_hn
        wn_h[1] = b_hn_1;
        wn_h[1] = sat_add(wn_h[1], fx_mult_round(w_hn_1_0, h_0));
        wn_h[1] = sat_add(wn_h[1], fx_mult_round(w_hn_1_1, h_1));
        wn_h[1] = sat_add(wn_h[1], fx_mult_round(w_hn_1_2, h_2));
        wn_h[1] = sat_add(wn_h[1], fx_mult_round(w_hn_1_3, h_3));
        wn_h[1] = sat_add(wn_h[1], fx_mult_round(w_hn_1_4, h_4));
        wn_h[1] = sat_add(wn_h[1], fx_mult_round(w_hn_1_5, h_5));
        wn_h[1] = sat_add(wn_h[1], fx_mult_round(w_hn_1_6, h_6));
        wn_h[1] = sat_add(wn_h[1], fx_mult_round(w_hn_1_7, h_7));

        // gated_h[1] = r_t ⊙ wn_h
        gated_h[1] = fx_mult_round(r_act[1], wn_h[1]);

        // n_sum[1] = W_in*x + b_in + gated_h
        n_sum[1] = b_in_1;
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_0, x_0));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_1, x_1));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_2, x_2));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_3, x_3));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_4, x_4));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_5, x_5));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_6, x_6));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_7, x_7));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_8, x_8));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_9, x_9));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_10, x_10));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_11, x_11));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_12, x_12));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_13, x_13));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_14, x_14));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_15, x_15));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_16, x_16));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_17, x_17));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_18, x_18));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_19, x_19));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_20, x_20));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_21, x_21));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_22, x_22));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_23, x_23));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_24, x_24));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_25, x_25));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_26, x_26));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_27, x_27));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_28, x_28));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_29, x_29));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_30, x_30));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_31, x_31));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_32, x_32));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_33, x_33));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_34, x_34));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_35, x_35));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_36, x_36));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_37, x_37));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_38, x_38));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_39, x_39));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_40, x_40));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_41, x_41));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_42, x_42));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_43, x_43));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_44, x_44));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_45, x_45));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_46, x_46));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_47, x_47));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_48, x_48));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_49, x_49));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_50, x_50));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_51, x_51));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_52, x_52));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_53, x_53));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_54, x_54));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_55, x_55));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_56, x_56));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_57, x_57));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_58, x_58));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_59, x_59));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_60, x_60));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_61, x_61));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_62, x_62));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_63, x_63));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_64, x_64));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_65, x_65));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_66, x_66));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_67, x_67));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_68, x_68));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_69, x_69));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_70, x_70));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_71, x_71));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_72, x_72));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_73, x_73));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_74, x_74));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_75, x_75));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_76, x_76));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_77, x_77));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_78, x_78));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_79, x_79));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_80, x_80));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_81, x_81));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_82, x_82));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_83, x_83));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_84, x_84));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_85, x_85));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_86, x_86));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_87, x_87));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_88, x_88));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_89, x_89));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_90, x_90));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_91, x_91));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_92, x_92));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_93, x_93));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_94, x_94));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_95, x_95));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_96, x_96));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_97, x_97));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_98, x_98));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_99, x_99));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_100, x_100));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_101, x_101));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_102, x_102));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_103, x_103));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_104, x_104));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_105, x_105));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_106, x_106));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_107, x_107));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_108, x_108));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_109, x_109));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_110, x_110));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_111, x_111));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_112, x_112));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_113, x_113));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_114, x_114));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_115, x_115));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_116, x_116));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_117, x_117));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_118, x_118));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_119, x_119));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_120, x_120));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_121, x_121));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_122, x_122));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_123, x_123));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_124, x_124));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_125, x_125));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_126, x_126));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_127, x_127));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_128, x_128));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_129, x_129));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_130, x_130));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_131, x_131));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_132, x_132));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_133, x_133));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_134, x_134));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_135, x_135));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_136, x_136));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_137, x_137));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_138, x_138));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_139, x_139));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_140, x_140));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_141, x_141));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_142, x_142));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_143, x_143));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_144, x_144));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_145, x_145));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_146, x_146));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_147, x_147));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_148, x_148));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_149, x_149));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_150, x_150));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_151, x_151));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_152, x_152));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_153, x_153));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_154, x_154));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_155, x_155));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_156, x_156));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_157, x_157));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_158, x_158));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_159, x_159));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_160, x_160));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_161, x_161));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_162, x_162));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_163, x_163));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_164, x_164));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_165, x_165));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_166, x_166));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_167, x_167));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_168, x_168));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_169, x_169));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_170, x_170));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_171, x_171));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_172, x_172));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_173, x_173));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_174, x_174));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_175, x_175));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_176, x_176));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_177, x_177));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_178, x_178));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_179, x_179));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_180, x_180));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_181, x_181));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_182, x_182));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_183, x_183));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_184, x_184));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_185, x_185));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_186, x_186));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_187, x_187));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_188, x_188));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_189, x_189));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_190, x_190));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_191, x_191));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_192, x_192));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_193, x_193));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_194, x_194));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_195, x_195));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_196, x_196));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_197, x_197));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_198, x_198));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_199, x_199));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_200, x_200));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_201, x_201));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_202, x_202));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_203, x_203));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_204, x_204));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_205, x_205));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_206, x_206));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_207, x_207));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_208, x_208));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_209, x_209));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_210, x_210));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_211, x_211));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_212, x_212));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_213, x_213));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_214, x_214));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_215, x_215));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_216, x_216));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_217, x_217));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_218, x_218));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_219, x_219));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_220, x_220));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_221, x_221));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_222, x_222));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_223, x_223));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_224, x_224));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_225, x_225));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_226, x_226));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_227, x_227));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_228, x_228));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_229, x_229));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_230, x_230));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_231, x_231));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_232, x_232));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_233, x_233));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_234, x_234));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_235, x_235));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_236, x_236));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_237, x_237));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_238, x_238));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_239, x_239));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_240, x_240));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_241, x_241));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_242, x_242));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_243, x_243));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_244, x_244));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_245, x_245));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_246, x_246));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_247, x_247));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_248, x_248));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_249, x_249));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_250, x_250));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_251, x_251));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_252, x_252));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_253, x_253));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_254, x_254));
        n_sum[1] = sat_add(n_sum[1], fx_mult_round(w_in_1_255, x_255));
        n_sum[1] = sat_add(n_sum[1], gated_h[1]);

        // wn_h[2] = W_hn*h + b_hn
        wn_h[2] = b_hn_2;
        wn_h[2] = sat_add(wn_h[2], fx_mult_round(w_hn_2_0, h_0));
        wn_h[2] = sat_add(wn_h[2], fx_mult_round(w_hn_2_1, h_1));
        wn_h[2] = sat_add(wn_h[2], fx_mult_round(w_hn_2_2, h_2));
        wn_h[2] = sat_add(wn_h[2], fx_mult_round(w_hn_2_3, h_3));
        wn_h[2] = sat_add(wn_h[2], fx_mult_round(w_hn_2_4, h_4));
        wn_h[2] = sat_add(wn_h[2], fx_mult_round(w_hn_2_5, h_5));
        wn_h[2] = sat_add(wn_h[2], fx_mult_round(w_hn_2_6, h_6));
        wn_h[2] = sat_add(wn_h[2], fx_mult_round(w_hn_2_7, h_7));

        // gated_h[2] = r_t ⊙ wn_h
        gated_h[2] = fx_mult_round(r_act[2], wn_h[2]);

        // n_sum[2] = W_in*x + b_in + gated_h
        n_sum[2] = b_in_2;
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_0, x_0));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_1, x_1));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_2, x_2));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_3, x_3));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_4, x_4));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_5, x_5));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_6, x_6));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_7, x_7));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_8, x_8));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_9, x_9));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_10, x_10));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_11, x_11));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_12, x_12));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_13, x_13));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_14, x_14));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_15, x_15));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_16, x_16));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_17, x_17));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_18, x_18));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_19, x_19));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_20, x_20));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_21, x_21));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_22, x_22));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_23, x_23));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_24, x_24));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_25, x_25));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_26, x_26));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_27, x_27));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_28, x_28));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_29, x_29));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_30, x_30));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_31, x_31));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_32, x_32));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_33, x_33));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_34, x_34));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_35, x_35));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_36, x_36));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_37, x_37));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_38, x_38));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_39, x_39));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_40, x_40));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_41, x_41));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_42, x_42));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_43, x_43));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_44, x_44));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_45, x_45));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_46, x_46));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_47, x_47));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_48, x_48));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_49, x_49));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_50, x_50));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_51, x_51));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_52, x_52));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_53, x_53));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_54, x_54));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_55, x_55));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_56, x_56));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_57, x_57));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_58, x_58));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_59, x_59));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_60, x_60));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_61, x_61));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_62, x_62));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_63, x_63));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_64, x_64));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_65, x_65));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_66, x_66));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_67, x_67));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_68, x_68));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_69, x_69));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_70, x_70));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_71, x_71));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_72, x_72));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_73, x_73));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_74, x_74));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_75, x_75));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_76, x_76));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_77, x_77));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_78, x_78));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_79, x_79));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_80, x_80));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_81, x_81));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_82, x_82));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_83, x_83));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_84, x_84));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_85, x_85));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_86, x_86));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_87, x_87));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_88, x_88));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_89, x_89));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_90, x_90));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_91, x_91));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_92, x_92));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_93, x_93));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_94, x_94));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_95, x_95));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_96, x_96));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_97, x_97));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_98, x_98));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_99, x_99));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_100, x_100));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_101, x_101));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_102, x_102));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_103, x_103));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_104, x_104));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_105, x_105));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_106, x_106));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_107, x_107));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_108, x_108));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_109, x_109));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_110, x_110));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_111, x_111));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_112, x_112));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_113, x_113));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_114, x_114));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_115, x_115));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_116, x_116));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_117, x_117));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_118, x_118));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_119, x_119));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_120, x_120));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_121, x_121));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_122, x_122));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_123, x_123));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_124, x_124));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_125, x_125));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_126, x_126));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_127, x_127));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_128, x_128));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_129, x_129));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_130, x_130));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_131, x_131));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_132, x_132));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_133, x_133));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_134, x_134));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_135, x_135));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_136, x_136));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_137, x_137));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_138, x_138));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_139, x_139));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_140, x_140));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_141, x_141));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_142, x_142));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_143, x_143));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_144, x_144));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_145, x_145));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_146, x_146));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_147, x_147));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_148, x_148));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_149, x_149));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_150, x_150));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_151, x_151));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_152, x_152));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_153, x_153));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_154, x_154));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_155, x_155));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_156, x_156));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_157, x_157));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_158, x_158));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_159, x_159));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_160, x_160));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_161, x_161));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_162, x_162));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_163, x_163));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_164, x_164));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_165, x_165));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_166, x_166));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_167, x_167));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_168, x_168));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_169, x_169));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_170, x_170));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_171, x_171));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_172, x_172));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_173, x_173));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_174, x_174));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_175, x_175));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_176, x_176));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_177, x_177));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_178, x_178));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_179, x_179));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_180, x_180));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_181, x_181));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_182, x_182));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_183, x_183));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_184, x_184));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_185, x_185));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_186, x_186));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_187, x_187));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_188, x_188));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_189, x_189));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_190, x_190));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_191, x_191));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_192, x_192));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_193, x_193));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_194, x_194));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_195, x_195));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_196, x_196));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_197, x_197));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_198, x_198));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_199, x_199));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_200, x_200));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_201, x_201));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_202, x_202));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_203, x_203));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_204, x_204));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_205, x_205));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_206, x_206));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_207, x_207));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_208, x_208));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_209, x_209));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_210, x_210));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_211, x_211));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_212, x_212));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_213, x_213));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_214, x_214));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_215, x_215));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_216, x_216));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_217, x_217));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_218, x_218));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_219, x_219));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_220, x_220));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_221, x_221));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_222, x_222));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_223, x_223));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_224, x_224));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_225, x_225));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_226, x_226));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_227, x_227));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_228, x_228));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_229, x_229));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_230, x_230));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_231, x_231));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_232, x_232));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_233, x_233));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_234, x_234));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_235, x_235));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_236, x_236));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_237, x_237));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_238, x_238));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_239, x_239));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_240, x_240));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_241, x_241));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_242, x_242));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_243, x_243));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_244, x_244));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_245, x_245));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_246, x_246));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_247, x_247));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_248, x_248));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_249, x_249));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_250, x_250));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_251, x_251));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_252, x_252));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_253, x_253));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_254, x_254));
        n_sum[2] = sat_add(n_sum[2], fx_mult_round(w_in_2_255, x_255));
        n_sum[2] = sat_add(n_sum[2], gated_h[2]);

        // wn_h[3] = W_hn*h + b_hn
        wn_h[3] = b_hn_3;
        wn_h[3] = sat_add(wn_h[3], fx_mult_round(w_hn_3_0, h_0));
        wn_h[3] = sat_add(wn_h[3], fx_mult_round(w_hn_3_1, h_1));
        wn_h[3] = sat_add(wn_h[3], fx_mult_round(w_hn_3_2, h_2));
        wn_h[3] = sat_add(wn_h[3], fx_mult_round(w_hn_3_3, h_3));
        wn_h[3] = sat_add(wn_h[3], fx_mult_round(w_hn_3_4, h_4));
        wn_h[3] = sat_add(wn_h[3], fx_mult_round(w_hn_3_5, h_5));
        wn_h[3] = sat_add(wn_h[3], fx_mult_round(w_hn_3_6, h_6));
        wn_h[3] = sat_add(wn_h[3], fx_mult_round(w_hn_3_7, h_7));

        // gated_h[3] = r_t ⊙ wn_h
        gated_h[3] = fx_mult_round(r_act[3], wn_h[3]);

        // n_sum[3] = W_in*x + b_in + gated_h
        n_sum[3] = b_in_3;
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_0, x_0));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_1, x_1));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_2, x_2));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_3, x_3));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_4, x_4));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_5, x_5));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_6, x_6));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_7, x_7));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_8, x_8));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_9, x_9));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_10, x_10));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_11, x_11));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_12, x_12));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_13, x_13));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_14, x_14));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_15, x_15));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_16, x_16));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_17, x_17));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_18, x_18));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_19, x_19));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_20, x_20));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_21, x_21));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_22, x_22));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_23, x_23));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_24, x_24));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_25, x_25));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_26, x_26));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_27, x_27));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_28, x_28));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_29, x_29));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_30, x_30));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_31, x_31));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_32, x_32));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_33, x_33));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_34, x_34));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_35, x_35));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_36, x_36));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_37, x_37));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_38, x_38));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_39, x_39));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_40, x_40));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_41, x_41));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_42, x_42));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_43, x_43));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_44, x_44));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_45, x_45));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_46, x_46));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_47, x_47));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_48, x_48));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_49, x_49));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_50, x_50));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_51, x_51));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_52, x_52));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_53, x_53));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_54, x_54));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_55, x_55));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_56, x_56));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_57, x_57));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_58, x_58));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_59, x_59));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_60, x_60));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_61, x_61));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_62, x_62));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_63, x_63));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_64, x_64));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_65, x_65));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_66, x_66));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_67, x_67));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_68, x_68));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_69, x_69));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_70, x_70));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_71, x_71));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_72, x_72));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_73, x_73));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_74, x_74));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_75, x_75));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_76, x_76));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_77, x_77));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_78, x_78));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_79, x_79));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_80, x_80));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_81, x_81));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_82, x_82));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_83, x_83));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_84, x_84));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_85, x_85));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_86, x_86));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_87, x_87));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_88, x_88));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_89, x_89));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_90, x_90));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_91, x_91));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_92, x_92));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_93, x_93));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_94, x_94));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_95, x_95));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_96, x_96));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_97, x_97));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_98, x_98));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_99, x_99));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_100, x_100));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_101, x_101));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_102, x_102));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_103, x_103));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_104, x_104));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_105, x_105));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_106, x_106));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_107, x_107));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_108, x_108));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_109, x_109));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_110, x_110));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_111, x_111));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_112, x_112));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_113, x_113));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_114, x_114));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_115, x_115));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_116, x_116));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_117, x_117));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_118, x_118));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_119, x_119));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_120, x_120));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_121, x_121));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_122, x_122));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_123, x_123));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_124, x_124));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_125, x_125));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_126, x_126));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_127, x_127));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_128, x_128));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_129, x_129));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_130, x_130));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_131, x_131));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_132, x_132));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_133, x_133));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_134, x_134));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_135, x_135));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_136, x_136));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_137, x_137));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_138, x_138));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_139, x_139));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_140, x_140));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_141, x_141));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_142, x_142));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_143, x_143));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_144, x_144));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_145, x_145));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_146, x_146));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_147, x_147));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_148, x_148));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_149, x_149));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_150, x_150));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_151, x_151));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_152, x_152));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_153, x_153));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_154, x_154));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_155, x_155));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_156, x_156));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_157, x_157));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_158, x_158));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_159, x_159));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_160, x_160));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_161, x_161));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_162, x_162));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_163, x_163));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_164, x_164));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_165, x_165));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_166, x_166));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_167, x_167));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_168, x_168));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_169, x_169));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_170, x_170));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_171, x_171));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_172, x_172));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_173, x_173));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_174, x_174));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_175, x_175));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_176, x_176));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_177, x_177));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_178, x_178));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_179, x_179));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_180, x_180));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_181, x_181));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_182, x_182));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_183, x_183));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_184, x_184));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_185, x_185));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_186, x_186));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_187, x_187));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_188, x_188));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_189, x_189));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_190, x_190));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_191, x_191));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_192, x_192));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_193, x_193));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_194, x_194));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_195, x_195));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_196, x_196));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_197, x_197));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_198, x_198));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_199, x_199));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_200, x_200));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_201, x_201));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_202, x_202));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_203, x_203));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_204, x_204));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_205, x_205));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_206, x_206));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_207, x_207));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_208, x_208));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_209, x_209));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_210, x_210));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_211, x_211));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_212, x_212));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_213, x_213));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_214, x_214));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_215, x_215));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_216, x_216));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_217, x_217));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_218, x_218));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_219, x_219));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_220, x_220));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_221, x_221));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_222, x_222));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_223, x_223));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_224, x_224));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_225, x_225));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_226, x_226));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_227, x_227));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_228, x_228));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_229, x_229));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_230, x_230));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_231, x_231));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_232, x_232));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_233, x_233));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_234, x_234));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_235, x_235));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_236, x_236));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_237, x_237));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_238, x_238));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_239, x_239));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_240, x_240));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_241, x_241));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_242, x_242));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_243, x_243));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_244, x_244));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_245, x_245));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_246, x_246));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_247, x_247));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_248, x_248));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_249, x_249));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_250, x_250));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_251, x_251));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_252, x_252));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_253, x_253));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_254, x_254));
        n_sum[3] = sat_add(n_sum[3], fx_mult_round(w_in_3_255, x_255));
        n_sum[3] = sat_add(n_sum[3], gated_h[3]);

        // wn_h[4] = W_hn*h + b_hn
        wn_h[4] = b_hn_4;
        wn_h[4] = sat_add(wn_h[4], fx_mult_round(w_hn_4_0, h_0));
        wn_h[4] = sat_add(wn_h[4], fx_mult_round(w_hn_4_1, h_1));
        wn_h[4] = sat_add(wn_h[4], fx_mult_round(w_hn_4_2, h_2));
        wn_h[4] = sat_add(wn_h[4], fx_mult_round(w_hn_4_3, h_3));
        wn_h[4] = sat_add(wn_h[4], fx_mult_round(w_hn_4_4, h_4));
        wn_h[4] = sat_add(wn_h[4], fx_mult_round(w_hn_4_5, h_5));
        wn_h[4] = sat_add(wn_h[4], fx_mult_round(w_hn_4_6, h_6));
        wn_h[4] = sat_add(wn_h[4], fx_mult_round(w_hn_4_7, h_7));

        // gated_h[4] = r_t ⊙ wn_h
        gated_h[4] = fx_mult_round(r_act[4], wn_h[4]);

        // n_sum[4] = W_in*x + b_in + gated_h
        n_sum[4] = b_in_4;
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_0, x_0));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_1, x_1));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_2, x_2));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_3, x_3));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_4, x_4));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_5, x_5));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_6, x_6));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_7, x_7));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_8, x_8));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_9, x_9));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_10, x_10));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_11, x_11));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_12, x_12));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_13, x_13));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_14, x_14));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_15, x_15));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_16, x_16));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_17, x_17));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_18, x_18));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_19, x_19));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_20, x_20));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_21, x_21));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_22, x_22));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_23, x_23));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_24, x_24));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_25, x_25));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_26, x_26));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_27, x_27));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_28, x_28));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_29, x_29));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_30, x_30));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_31, x_31));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_32, x_32));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_33, x_33));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_34, x_34));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_35, x_35));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_36, x_36));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_37, x_37));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_38, x_38));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_39, x_39));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_40, x_40));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_41, x_41));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_42, x_42));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_43, x_43));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_44, x_44));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_45, x_45));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_46, x_46));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_47, x_47));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_48, x_48));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_49, x_49));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_50, x_50));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_51, x_51));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_52, x_52));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_53, x_53));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_54, x_54));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_55, x_55));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_56, x_56));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_57, x_57));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_58, x_58));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_59, x_59));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_60, x_60));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_61, x_61));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_62, x_62));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_63, x_63));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_64, x_64));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_65, x_65));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_66, x_66));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_67, x_67));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_68, x_68));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_69, x_69));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_70, x_70));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_71, x_71));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_72, x_72));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_73, x_73));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_74, x_74));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_75, x_75));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_76, x_76));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_77, x_77));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_78, x_78));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_79, x_79));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_80, x_80));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_81, x_81));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_82, x_82));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_83, x_83));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_84, x_84));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_85, x_85));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_86, x_86));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_87, x_87));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_88, x_88));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_89, x_89));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_90, x_90));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_91, x_91));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_92, x_92));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_93, x_93));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_94, x_94));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_95, x_95));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_96, x_96));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_97, x_97));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_98, x_98));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_99, x_99));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_100, x_100));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_101, x_101));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_102, x_102));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_103, x_103));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_104, x_104));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_105, x_105));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_106, x_106));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_107, x_107));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_108, x_108));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_109, x_109));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_110, x_110));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_111, x_111));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_112, x_112));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_113, x_113));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_114, x_114));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_115, x_115));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_116, x_116));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_117, x_117));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_118, x_118));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_119, x_119));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_120, x_120));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_121, x_121));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_122, x_122));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_123, x_123));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_124, x_124));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_125, x_125));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_126, x_126));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_127, x_127));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_128, x_128));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_129, x_129));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_130, x_130));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_131, x_131));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_132, x_132));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_133, x_133));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_134, x_134));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_135, x_135));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_136, x_136));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_137, x_137));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_138, x_138));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_139, x_139));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_140, x_140));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_141, x_141));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_142, x_142));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_143, x_143));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_144, x_144));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_145, x_145));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_146, x_146));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_147, x_147));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_148, x_148));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_149, x_149));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_150, x_150));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_151, x_151));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_152, x_152));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_153, x_153));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_154, x_154));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_155, x_155));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_156, x_156));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_157, x_157));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_158, x_158));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_159, x_159));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_160, x_160));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_161, x_161));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_162, x_162));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_163, x_163));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_164, x_164));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_165, x_165));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_166, x_166));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_167, x_167));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_168, x_168));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_169, x_169));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_170, x_170));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_171, x_171));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_172, x_172));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_173, x_173));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_174, x_174));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_175, x_175));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_176, x_176));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_177, x_177));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_178, x_178));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_179, x_179));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_180, x_180));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_181, x_181));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_182, x_182));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_183, x_183));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_184, x_184));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_185, x_185));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_186, x_186));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_187, x_187));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_188, x_188));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_189, x_189));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_190, x_190));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_191, x_191));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_192, x_192));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_193, x_193));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_194, x_194));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_195, x_195));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_196, x_196));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_197, x_197));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_198, x_198));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_199, x_199));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_200, x_200));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_201, x_201));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_202, x_202));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_203, x_203));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_204, x_204));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_205, x_205));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_206, x_206));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_207, x_207));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_208, x_208));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_209, x_209));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_210, x_210));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_211, x_211));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_212, x_212));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_213, x_213));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_214, x_214));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_215, x_215));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_216, x_216));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_217, x_217));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_218, x_218));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_219, x_219));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_220, x_220));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_221, x_221));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_222, x_222));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_223, x_223));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_224, x_224));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_225, x_225));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_226, x_226));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_227, x_227));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_228, x_228));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_229, x_229));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_230, x_230));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_231, x_231));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_232, x_232));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_233, x_233));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_234, x_234));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_235, x_235));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_236, x_236));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_237, x_237));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_238, x_238));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_239, x_239));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_240, x_240));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_241, x_241));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_242, x_242));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_243, x_243));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_244, x_244));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_245, x_245));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_246, x_246));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_247, x_247));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_248, x_248));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_249, x_249));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_250, x_250));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_251, x_251));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_252, x_252));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_253, x_253));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_254, x_254));
        n_sum[4] = sat_add(n_sum[4], fx_mult_round(w_in_4_255, x_255));
        n_sum[4] = sat_add(n_sum[4], gated_h[4]);

        // wn_h[5] = W_hn*h + b_hn
        wn_h[5] = b_hn_5;
        wn_h[5] = sat_add(wn_h[5], fx_mult_round(w_hn_5_0, h_0));
        wn_h[5] = sat_add(wn_h[5], fx_mult_round(w_hn_5_1, h_1));
        wn_h[5] = sat_add(wn_h[5], fx_mult_round(w_hn_5_2, h_2));
        wn_h[5] = sat_add(wn_h[5], fx_mult_round(w_hn_5_3, h_3));
        wn_h[5] = sat_add(wn_h[5], fx_mult_round(w_hn_5_4, h_4));
        wn_h[5] = sat_add(wn_h[5], fx_mult_round(w_hn_5_5, h_5));
        wn_h[5] = sat_add(wn_h[5], fx_mult_round(w_hn_5_6, h_6));
        wn_h[5] = sat_add(wn_h[5], fx_mult_round(w_hn_5_7, h_7));

        // gated_h[5] = r_t ⊙ wn_h
        gated_h[5] = fx_mult_round(r_act[5], wn_h[5]);

        // n_sum[5] = W_in*x + b_in + gated_h
        n_sum[5] = b_in_5;
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_0, x_0));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_1, x_1));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_2, x_2));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_3, x_3));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_4, x_4));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_5, x_5));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_6, x_6));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_7, x_7));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_8, x_8));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_9, x_9));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_10, x_10));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_11, x_11));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_12, x_12));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_13, x_13));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_14, x_14));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_15, x_15));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_16, x_16));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_17, x_17));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_18, x_18));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_19, x_19));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_20, x_20));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_21, x_21));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_22, x_22));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_23, x_23));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_24, x_24));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_25, x_25));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_26, x_26));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_27, x_27));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_28, x_28));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_29, x_29));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_30, x_30));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_31, x_31));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_32, x_32));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_33, x_33));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_34, x_34));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_35, x_35));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_36, x_36));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_37, x_37));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_38, x_38));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_39, x_39));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_40, x_40));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_41, x_41));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_42, x_42));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_43, x_43));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_44, x_44));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_45, x_45));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_46, x_46));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_47, x_47));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_48, x_48));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_49, x_49));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_50, x_50));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_51, x_51));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_52, x_52));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_53, x_53));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_54, x_54));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_55, x_55));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_56, x_56));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_57, x_57));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_58, x_58));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_59, x_59));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_60, x_60));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_61, x_61));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_62, x_62));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_63, x_63));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_64, x_64));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_65, x_65));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_66, x_66));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_67, x_67));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_68, x_68));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_69, x_69));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_70, x_70));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_71, x_71));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_72, x_72));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_73, x_73));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_74, x_74));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_75, x_75));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_76, x_76));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_77, x_77));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_78, x_78));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_79, x_79));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_80, x_80));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_81, x_81));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_82, x_82));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_83, x_83));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_84, x_84));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_85, x_85));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_86, x_86));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_87, x_87));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_88, x_88));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_89, x_89));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_90, x_90));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_91, x_91));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_92, x_92));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_93, x_93));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_94, x_94));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_95, x_95));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_96, x_96));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_97, x_97));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_98, x_98));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_99, x_99));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_100, x_100));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_101, x_101));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_102, x_102));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_103, x_103));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_104, x_104));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_105, x_105));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_106, x_106));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_107, x_107));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_108, x_108));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_109, x_109));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_110, x_110));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_111, x_111));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_112, x_112));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_113, x_113));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_114, x_114));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_115, x_115));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_116, x_116));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_117, x_117));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_118, x_118));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_119, x_119));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_120, x_120));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_121, x_121));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_122, x_122));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_123, x_123));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_124, x_124));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_125, x_125));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_126, x_126));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_127, x_127));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_128, x_128));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_129, x_129));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_130, x_130));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_131, x_131));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_132, x_132));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_133, x_133));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_134, x_134));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_135, x_135));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_136, x_136));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_137, x_137));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_138, x_138));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_139, x_139));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_140, x_140));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_141, x_141));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_142, x_142));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_143, x_143));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_144, x_144));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_145, x_145));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_146, x_146));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_147, x_147));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_148, x_148));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_149, x_149));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_150, x_150));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_151, x_151));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_152, x_152));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_153, x_153));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_154, x_154));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_155, x_155));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_156, x_156));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_157, x_157));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_158, x_158));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_159, x_159));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_160, x_160));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_161, x_161));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_162, x_162));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_163, x_163));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_164, x_164));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_165, x_165));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_166, x_166));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_167, x_167));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_168, x_168));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_169, x_169));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_170, x_170));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_171, x_171));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_172, x_172));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_173, x_173));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_174, x_174));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_175, x_175));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_176, x_176));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_177, x_177));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_178, x_178));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_179, x_179));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_180, x_180));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_181, x_181));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_182, x_182));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_183, x_183));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_184, x_184));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_185, x_185));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_186, x_186));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_187, x_187));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_188, x_188));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_189, x_189));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_190, x_190));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_191, x_191));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_192, x_192));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_193, x_193));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_194, x_194));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_195, x_195));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_196, x_196));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_197, x_197));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_198, x_198));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_199, x_199));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_200, x_200));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_201, x_201));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_202, x_202));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_203, x_203));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_204, x_204));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_205, x_205));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_206, x_206));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_207, x_207));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_208, x_208));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_209, x_209));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_210, x_210));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_211, x_211));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_212, x_212));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_213, x_213));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_214, x_214));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_215, x_215));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_216, x_216));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_217, x_217));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_218, x_218));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_219, x_219));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_220, x_220));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_221, x_221));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_222, x_222));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_223, x_223));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_224, x_224));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_225, x_225));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_226, x_226));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_227, x_227));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_228, x_228));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_229, x_229));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_230, x_230));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_231, x_231));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_232, x_232));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_233, x_233));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_234, x_234));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_235, x_235));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_236, x_236));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_237, x_237));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_238, x_238));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_239, x_239));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_240, x_240));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_241, x_241));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_242, x_242));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_243, x_243));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_244, x_244));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_245, x_245));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_246, x_246));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_247, x_247));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_248, x_248));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_249, x_249));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_250, x_250));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_251, x_251));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_252, x_252));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_253, x_253));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_254, x_254));
        n_sum[5] = sat_add(n_sum[5], fx_mult_round(w_in_5_255, x_255));
        n_sum[5] = sat_add(n_sum[5], gated_h[5]);

        // wn_h[6] = W_hn*h + b_hn
        wn_h[6] = b_hn_6;
        wn_h[6] = sat_add(wn_h[6], fx_mult_round(w_hn_6_0, h_0));
        wn_h[6] = sat_add(wn_h[6], fx_mult_round(w_hn_6_1, h_1));
        wn_h[6] = sat_add(wn_h[6], fx_mult_round(w_hn_6_2, h_2));
        wn_h[6] = sat_add(wn_h[6], fx_mult_round(w_hn_6_3, h_3));
        wn_h[6] = sat_add(wn_h[6], fx_mult_round(w_hn_6_4, h_4));
        wn_h[6] = sat_add(wn_h[6], fx_mult_round(w_hn_6_5, h_5));
        wn_h[6] = sat_add(wn_h[6], fx_mult_round(w_hn_6_6, h_6));
        wn_h[6] = sat_add(wn_h[6], fx_mult_round(w_hn_6_7, h_7));

        // gated_h[6] = r_t ⊙ wn_h
        gated_h[6] = fx_mult_round(r_act[6], wn_h[6]);

        // n_sum[6] = W_in*x + b_in + gated_h
        n_sum[6] = b_in_6;
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_0, x_0));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_1, x_1));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_2, x_2));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_3, x_3));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_4, x_4));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_5, x_5));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_6, x_6));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_7, x_7));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_8, x_8));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_9, x_9));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_10, x_10));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_11, x_11));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_12, x_12));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_13, x_13));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_14, x_14));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_15, x_15));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_16, x_16));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_17, x_17));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_18, x_18));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_19, x_19));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_20, x_20));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_21, x_21));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_22, x_22));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_23, x_23));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_24, x_24));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_25, x_25));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_26, x_26));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_27, x_27));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_28, x_28));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_29, x_29));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_30, x_30));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_31, x_31));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_32, x_32));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_33, x_33));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_34, x_34));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_35, x_35));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_36, x_36));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_37, x_37));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_38, x_38));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_39, x_39));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_40, x_40));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_41, x_41));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_42, x_42));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_43, x_43));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_44, x_44));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_45, x_45));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_46, x_46));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_47, x_47));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_48, x_48));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_49, x_49));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_50, x_50));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_51, x_51));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_52, x_52));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_53, x_53));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_54, x_54));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_55, x_55));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_56, x_56));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_57, x_57));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_58, x_58));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_59, x_59));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_60, x_60));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_61, x_61));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_62, x_62));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_63, x_63));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_64, x_64));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_65, x_65));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_66, x_66));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_67, x_67));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_68, x_68));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_69, x_69));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_70, x_70));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_71, x_71));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_72, x_72));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_73, x_73));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_74, x_74));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_75, x_75));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_76, x_76));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_77, x_77));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_78, x_78));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_79, x_79));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_80, x_80));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_81, x_81));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_82, x_82));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_83, x_83));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_84, x_84));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_85, x_85));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_86, x_86));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_87, x_87));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_88, x_88));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_89, x_89));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_90, x_90));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_91, x_91));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_92, x_92));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_93, x_93));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_94, x_94));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_95, x_95));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_96, x_96));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_97, x_97));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_98, x_98));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_99, x_99));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_100, x_100));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_101, x_101));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_102, x_102));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_103, x_103));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_104, x_104));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_105, x_105));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_106, x_106));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_107, x_107));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_108, x_108));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_109, x_109));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_110, x_110));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_111, x_111));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_112, x_112));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_113, x_113));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_114, x_114));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_115, x_115));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_116, x_116));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_117, x_117));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_118, x_118));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_119, x_119));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_120, x_120));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_121, x_121));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_122, x_122));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_123, x_123));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_124, x_124));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_125, x_125));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_126, x_126));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_127, x_127));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_128, x_128));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_129, x_129));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_130, x_130));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_131, x_131));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_132, x_132));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_133, x_133));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_134, x_134));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_135, x_135));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_136, x_136));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_137, x_137));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_138, x_138));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_139, x_139));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_140, x_140));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_141, x_141));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_142, x_142));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_143, x_143));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_144, x_144));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_145, x_145));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_146, x_146));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_147, x_147));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_148, x_148));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_149, x_149));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_150, x_150));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_151, x_151));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_152, x_152));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_153, x_153));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_154, x_154));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_155, x_155));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_156, x_156));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_157, x_157));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_158, x_158));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_159, x_159));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_160, x_160));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_161, x_161));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_162, x_162));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_163, x_163));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_164, x_164));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_165, x_165));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_166, x_166));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_167, x_167));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_168, x_168));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_169, x_169));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_170, x_170));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_171, x_171));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_172, x_172));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_173, x_173));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_174, x_174));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_175, x_175));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_176, x_176));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_177, x_177));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_178, x_178));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_179, x_179));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_180, x_180));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_181, x_181));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_182, x_182));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_183, x_183));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_184, x_184));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_185, x_185));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_186, x_186));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_187, x_187));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_188, x_188));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_189, x_189));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_190, x_190));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_191, x_191));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_192, x_192));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_193, x_193));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_194, x_194));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_195, x_195));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_196, x_196));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_197, x_197));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_198, x_198));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_199, x_199));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_200, x_200));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_201, x_201));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_202, x_202));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_203, x_203));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_204, x_204));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_205, x_205));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_206, x_206));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_207, x_207));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_208, x_208));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_209, x_209));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_210, x_210));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_211, x_211));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_212, x_212));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_213, x_213));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_214, x_214));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_215, x_215));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_216, x_216));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_217, x_217));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_218, x_218));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_219, x_219));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_220, x_220));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_221, x_221));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_222, x_222));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_223, x_223));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_224, x_224));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_225, x_225));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_226, x_226));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_227, x_227));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_228, x_228));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_229, x_229));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_230, x_230));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_231, x_231));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_232, x_232));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_233, x_233));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_234, x_234));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_235, x_235));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_236, x_236));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_237, x_237));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_238, x_238));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_239, x_239));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_240, x_240));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_241, x_241));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_242, x_242));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_243, x_243));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_244, x_244));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_245, x_245));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_246, x_246));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_247, x_247));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_248, x_248));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_249, x_249));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_250, x_250));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_251, x_251));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_252, x_252));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_253, x_253));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_254, x_254));
        n_sum[6] = sat_add(n_sum[6], fx_mult_round(w_in_6_255, x_255));
        n_sum[6] = sat_add(n_sum[6], gated_h[6]);

        // wn_h[7] = W_hn*h + b_hn
        wn_h[7] = b_hn_7;
        wn_h[7] = sat_add(wn_h[7], fx_mult_round(w_hn_7_0, h_0));
        wn_h[7] = sat_add(wn_h[7], fx_mult_round(w_hn_7_1, h_1));
        wn_h[7] = sat_add(wn_h[7], fx_mult_round(w_hn_7_2, h_2));
        wn_h[7] = sat_add(wn_h[7], fx_mult_round(w_hn_7_3, h_3));
        wn_h[7] = sat_add(wn_h[7], fx_mult_round(w_hn_7_4, h_4));
        wn_h[7] = sat_add(wn_h[7], fx_mult_round(w_hn_7_5, h_5));
        wn_h[7] = sat_add(wn_h[7], fx_mult_round(w_hn_7_6, h_6));
        wn_h[7] = sat_add(wn_h[7], fx_mult_round(w_hn_7_7, h_7));

        // gated_h[7] = r_t ⊙ wn_h
        gated_h[7] = fx_mult_round(r_act[7], wn_h[7]);

        // n_sum[7] = W_in*x + b_in + gated_h
        n_sum[7] = b_in_7;
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_0, x_0));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_1, x_1));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_2, x_2));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_3, x_3));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_4, x_4));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_5, x_5));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_6, x_6));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_7, x_7));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_8, x_8));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_9, x_9));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_10, x_10));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_11, x_11));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_12, x_12));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_13, x_13));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_14, x_14));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_15, x_15));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_16, x_16));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_17, x_17));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_18, x_18));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_19, x_19));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_20, x_20));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_21, x_21));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_22, x_22));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_23, x_23));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_24, x_24));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_25, x_25));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_26, x_26));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_27, x_27));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_28, x_28));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_29, x_29));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_30, x_30));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_31, x_31));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_32, x_32));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_33, x_33));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_34, x_34));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_35, x_35));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_36, x_36));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_37, x_37));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_38, x_38));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_39, x_39));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_40, x_40));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_41, x_41));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_42, x_42));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_43, x_43));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_44, x_44));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_45, x_45));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_46, x_46));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_47, x_47));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_48, x_48));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_49, x_49));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_50, x_50));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_51, x_51));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_52, x_52));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_53, x_53));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_54, x_54));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_55, x_55));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_56, x_56));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_57, x_57));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_58, x_58));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_59, x_59));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_60, x_60));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_61, x_61));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_62, x_62));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_63, x_63));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_64, x_64));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_65, x_65));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_66, x_66));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_67, x_67));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_68, x_68));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_69, x_69));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_70, x_70));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_71, x_71));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_72, x_72));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_73, x_73));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_74, x_74));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_75, x_75));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_76, x_76));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_77, x_77));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_78, x_78));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_79, x_79));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_80, x_80));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_81, x_81));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_82, x_82));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_83, x_83));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_84, x_84));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_85, x_85));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_86, x_86));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_87, x_87));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_88, x_88));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_89, x_89));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_90, x_90));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_91, x_91));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_92, x_92));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_93, x_93));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_94, x_94));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_95, x_95));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_96, x_96));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_97, x_97));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_98, x_98));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_99, x_99));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_100, x_100));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_101, x_101));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_102, x_102));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_103, x_103));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_104, x_104));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_105, x_105));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_106, x_106));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_107, x_107));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_108, x_108));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_109, x_109));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_110, x_110));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_111, x_111));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_112, x_112));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_113, x_113));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_114, x_114));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_115, x_115));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_116, x_116));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_117, x_117));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_118, x_118));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_119, x_119));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_120, x_120));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_121, x_121));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_122, x_122));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_123, x_123));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_124, x_124));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_125, x_125));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_126, x_126));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_127, x_127));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_128, x_128));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_129, x_129));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_130, x_130));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_131, x_131));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_132, x_132));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_133, x_133));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_134, x_134));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_135, x_135));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_136, x_136));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_137, x_137));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_138, x_138));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_139, x_139));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_140, x_140));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_141, x_141));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_142, x_142));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_143, x_143));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_144, x_144));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_145, x_145));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_146, x_146));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_147, x_147));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_148, x_148));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_149, x_149));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_150, x_150));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_151, x_151));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_152, x_152));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_153, x_153));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_154, x_154));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_155, x_155));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_156, x_156));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_157, x_157));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_158, x_158));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_159, x_159));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_160, x_160));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_161, x_161));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_162, x_162));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_163, x_163));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_164, x_164));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_165, x_165));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_166, x_166));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_167, x_167));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_168, x_168));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_169, x_169));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_170, x_170));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_171, x_171));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_172, x_172));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_173, x_173));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_174, x_174));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_175, x_175));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_176, x_176));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_177, x_177));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_178, x_178));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_179, x_179));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_180, x_180));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_181, x_181));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_182, x_182));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_183, x_183));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_184, x_184));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_185, x_185));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_186, x_186));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_187, x_187));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_188, x_188));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_189, x_189));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_190, x_190));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_191, x_191));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_192, x_192));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_193, x_193));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_194, x_194));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_195, x_195));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_196, x_196));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_197, x_197));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_198, x_198));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_199, x_199));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_200, x_200));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_201, x_201));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_202, x_202));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_203, x_203));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_204, x_204));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_205, x_205));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_206, x_206));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_207, x_207));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_208, x_208));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_209, x_209));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_210, x_210));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_211, x_211));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_212, x_212));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_213, x_213));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_214, x_214));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_215, x_215));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_216, x_216));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_217, x_217));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_218, x_218));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_219, x_219));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_220, x_220));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_221, x_221));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_222, x_222));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_223, x_223));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_224, x_224));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_225, x_225));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_226, x_226));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_227, x_227));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_228, x_228));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_229, x_229));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_230, x_230));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_231, x_231));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_232, x_232));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_233, x_233));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_234, x_234));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_235, x_235));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_236, x_236));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_237, x_237));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_238, x_238));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_239, x_239));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_240, x_240));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_241, x_241));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_242, x_242));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_243, x_243));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_244, x_244));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_245, x_245));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_246, x_246));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_247, x_247));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_248, x_248));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_249, x_249));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_250, x_250));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_251, x_251));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_252, x_252));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_253, x_253));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_254, x_254));
        n_sum[7] = sat_add(n_sum[7], fx_mult_round(w_in_7_255, x_255));
        n_sum[7] = sat_add(n_sum[7], gated_h[7]);

    end

    tanh #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) tanh_n0 (
         .reset(reset), .x(n_sum[0]), .y(n_act[0])
    );
    tanh #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) tanh_n1 (
         .reset(reset), .x(n_sum[1]), .y(n_act[1])
    );
    tanh #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) tanh_n2 (
         .reset(reset), .x(n_sum[2]), .y(n_act[2])
    );
    tanh #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) tanh_n3 (
         .reset(reset), .x(n_sum[3]), .y(n_act[3])
    );
    tanh #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) tanh_n4 (
         .reset(reset), .x(n_sum[4]), .y(n_act[4])
    );
    tanh #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) tanh_n5 (
         .reset(reset), .x(n_sum[5]), .y(n_act[5])
    );
    tanh #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) tanh_n6 (
         .reset(reset), .x(n_sum[6]), .y(n_act[6])
    );
    tanh #(.INT_WIDTH(INT_WIDTH), .FRAC_WIDTH(FRAC_WIDTH)) tanh_n7 (
         .reset(reset), .x(n_sum[7]), .y(n_act[7])
    );

    // Final hidden state update
    // Hidden state update: h_t = (1 - z_t) ⊙ n_t + z_t ⊙ h_{t-1}
    logic signed [WIDTH-1:0] one_minus_z[8];
    logic signed [WIDTH-1:0] part1[8], part2[8];
    logic signed [WIDTH-1:0] h_new[8];

    always_comb begin
        one_minus_z[0] = sat_add(ONE, -z_act[0]);
        part1[0] = fx_mult_round(one_minus_z[0], n_act[0]);
        part2[0] = fx_mult_round(z_act[0], h_0);
        h_new[0] = sat_add(part1[0], part2[0]);
        one_minus_z[1] = sat_add(ONE, -z_act[1]);
        part1[1] = fx_mult_round(one_minus_z[1], n_act[1]);
        part2[1] = fx_mult_round(z_act[1], h_1);
        h_new[1] = sat_add(part1[1], part2[1]);
        one_minus_z[2] = sat_add(ONE, -z_act[2]);
        part1[2] = fx_mult_round(one_minus_z[2], n_act[2]);
        part2[2] = fx_mult_round(z_act[2], h_2);
        h_new[2] = sat_add(part1[2], part2[2]);
        one_minus_z[3] = sat_add(ONE, -z_act[3]);
        part1[3] = fx_mult_round(one_minus_z[3], n_act[3]);
        part2[3] = fx_mult_round(z_act[3], h_3);
        h_new[3] = sat_add(part1[3], part2[3]);
        one_minus_z[4] = sat_add(ONE, -z_act[4]);
        part1[4] = fx_mult_round(one_minus_z[4], n_act[4]);
        part2[4] = fx_mult_round(z_act[4], h_4);
        h_new[4] = sat_add(part1[4], part2[4]);
        one_minus_z[5] = sat_add(ONE, -z_act[5]);
        part1[5] = fx_mult_round(one_minus_z[5], n_act[5]);
        part2[5] = fx_mult_round(z_act[5], h_5);
        h_new[5] = sat_add(part1[5], part2[5]);
        one_minus_z[6] = sat_add(ONE, -z_act[6]);
        part1[6] = fx_mult_round(one_minus_z[6], n_act[6]);
        part2[6] = fx_mult_round(z_act[6], h_6);
        h_new[6] = sat_add(part1[6], part2[6]);
        one_minus_z[7] = sat_add(ONE, -z_act[7]);
        part1[7] = fx_mult_round(one_minus_z[7], n_act[7]);
        part2[7] = fx_mult_round(z_act[7], h_7);
        h_new[7] = sat_add(part1[7], part2[7]);
    end

    // Register outputs
    always_ff @(posedge clk or posedge reset) begin
        if (reset) begin
            y_0 <= '0;
            y_1 <= '0;
            y_2 <= '0;
            y_3 <= '0;
            y_4 <= '0;
            y_5 <= '0;
            y_6 <= '0;
            y_7 <= '0;
        end else begin
            y_0 <= h_new[0];
            y_1 <= h_new[1];
            y_2 <= h_new[2];
            y_3 <= h_new[3];
            y_4 <= h_new[4];
            y_5 <= h_new[5];
            y_6 <= h_new[6];
            y_7 <= h_new[7];
        end
    end

endmodule
