`timescale 1ns / 1ps

module gru_tb;

// Parameters
parameter int INT_WIDTH  = 4;
parameter int FRAC_WIDTH = 5;
parameter int WIDTH      = INT_WIDTH + FRAC_WIDTH;
parameter real CLK_PERIOD = 10.0;

// Clock and reset
logic clk;
logic reset;

// Inputs
logic signed [WIDTH-1:0] x_0 = 0;
logic signed [WIDTH-1:0] x_1 = 0;
logic signed [WIDTH-1:0] x_2 = 0;
logic signed [WIDTH-1:0] x_3 = 0;
logic signed [WIDTH-1:0] x_4 = 0;
logic signed [WIDTH-1:0] x_5 = 0;
logic signed [WIDTH-1:0] x_6 = 0;
logic signed [WIDTH-1:0] x_7 = 0;
logic signed [WIDTH-1:0] x_8 = 0;
logic signed [WIDTH-1:0] x_9 = 0;
logic signed [WIDTH-1:0] x_10 = 0;
logic signed [WIDTH-1:0] x_11 = 0;
logic signed [WIDTH-1:0] x_12 = 0;
logic signed [WIDTH-1:0] x_13 = 0;
logic signed [WIDTH-1:0] x_14 = 0;
logic signed [WIDTH-1:0] x_15 = 0;
logic signed [WIDTH-1:0] x_16 = 0;
logic signed [WIDTH-1:0] x_17 = 0;
logic signed [WIDTH-1:0] x_18 = 0;
logic signed [WIDTH-1:0] x_19 = 0;
logic signed [WIDTH-1:0] x_20 = 0;
logic signed [WIDTH-1:0] x_21 = 0;
logic signed [WIDTH-1:0] x_22 = 0;
logic signed [WIDTH-1:0] x_23 = 0;
logic signed [WIDTH-1:0] x_24 = 0;
logic signed [WIDTH-1:0] x_25 = 0;
logic signed [WIDTH-1:0] x_26 = 0;
logic signed [WIDTH-1:0] x_27 = 0;
logic signed [WIDTH-1:0] x_28 = 0;
logic signed [WIDTH-1:0] x_29 = 0;
logic signed [WIDTH-1:0] x_30 = 0;
logic signed [WIDTH-1:0] x_31 = 0;
logic signed [WIDTH-1:0] x_32 = 0;
logic signed [WIDTH-1:0] x_33 = 0;
logic signed [WIDTH-1:0] x_34 = 0;
logic signed [WIDTH-1:0] x_35 = 0;
logic signed [WIDTH-1:0] x_36 = 0;
logic signed [WIDTH-1:0] x_37 = 0;
logic signed [WIDTH-1:0] x_38 = 0;
logic signed [WIDTH-1:0] x_39 = 0;
logic signed [WIDTH-1:0] x_40 = 0;
logic signed [WIDTH-1:0] x_41 = 0;
logic signed [WIDTH-1:0] x_42 = 0;
logic signed [WIDTH-1:0] x_43 = 0;
logic signed [WIDTH-1:0] x_44 = 0;
logic signed [WIDTH-1:0] x_45 = 0;
logic signed [WIDTH-1:0] x_46 = 0;
logic signed [WIDTH-1:0] x_47 = 0;
logic signed [WIDTH-1:0] x_48 = 0;
logic signed [WIDTH-1:0] x_49 = 0;
logic signed [WIDTH-1:0] x_50 = 0;
logic signed [WIDTH-1:0] x_51 = 0;
logic signed [WIDTH-1:0] x_52 = 0;
logic signed [WIDTH-1:0] x_53 = 0;
logic signed [WIDTH-1:0] x_54 = 0;
logic signed [WIDTH-1:0] x_55 = 0;
logic signed [WIDTH-1:0] x_56 = 0;
logic signed [WIDTH-1:0] x_57 = 0;
logic signed [WIDTH-1:0] x_58 = 0;
logic signed [WIDTH-1:0] x_59 = 0;
logic signed [WIDTH-1:0] x_60 = 0;
logic signed [WIDTH-1:0] x_61 = 0;
logic signed [WIDTH-1:0] x_62 = 0;
logic signed [WIDTH-1:0] x_63 = 0;
logic signed [WIDTH-1:0] x_64 = 0;
logic signed [WIDTH-1:0] x_65 = 0;
logic signed [WIDTH-1:0] x_66 = 0;
logic signed [WIDTH-1:0] x_67 = 0;
logic signed [WIDTH-1:0] x_68 = 0;
logic signed [WIDTH-1:0] x_69 = 0;
logic signed [WIDTH-1:0] x_70 = 0;
logic signed [WIDTH-1:0] x_71 = 0;
logic signed [WIDTH-1:0] x_72 = 0;
logic signed [WIDTH-1:0] x_73 = 0;
logic signed [WIDTH-1:0] x_74 = 0;
logic signed [WIDTH-1:0] x_75 = 0;
logic signed [WIDTH-1:0] x_76 = 0;
logic signed [WIDTH-1:0] x_77 = 0;
logic signed [WIDTH-1:0] x_78 = 0;
logic signed [WIDTH-1:0] x_79 = 0;
logic signed [WIDTH-1:0] x_80 = 0;
logic signed [WIDTH-1:0] x_81 = 0;
logic signed [WIDTH-1:0] x_82 = 0;
logic signed [WIDTH-1:0] x_83 = 0;
logic signed [WIDTH-1:0] x_84 = 0;
logic signed [WIDTH-1:0] x_85 = 0;
logic signed [WIDTH-1:0] x_86 = 0;
logic signed [WIDTH-1:0] x_87 = 0;
logic signed [WIDTH-1:0] x_88 = 0;
logic signed [WIDTH-1:0] x_89 = 0;
logic signed [WIDTH-1:0] x_90 = 0;
logic signed [WIDTH-1:0] x_91 = 0;
logic signed [WIDTH-1:0] x_92 = 0;
logic signed [WIDTH-1:0] x_93 = 0;
logic signed [WIDTH-1:0] x_94 = 0;
logic signed [WIDTH-1:0] x_95 = 0;
logic signed [WIDTH-1:0] x_96 = 0;
logic signed [WIDTH-1:0] x_97 = 0;
logic signed [WIDTH-1:0] x_98 = 0;
logic signed [WIDTH-1:0] x_99 = 0;
logic signed [WIDTH-1:0] x_100 = 0;
logic signed [WIDTH-1:0] x_101 = 0;
logic signed [WIDTH-1:0] x_102 = 0;
logic signed [WIDTH-1:0] x_103 = 0;
logic signed [WIDTH-1:0] x_104 = 0;
logic signed [WIDTH-1:0] x_105 = 0;
logic signed [WIDTH-1:0] x_106 = 0;
logic signed [WIDTH-1:0] x_107 = 0;
logic signed [WIDTH-1:0] x_108 = 0;
logic signed [WIDTH-1:0] x_109 = 0;
logic signed [WIDTH-1:0] x_110 = 0;
logic signed [WIDTH-1:0] x_111 = 0;
logic signed [WIDTH-1:0] x_112 = 0;
logic signed [WIDTH-1:0] x_113 = 0;
logic signed [WIDTH-1:0] x_114 = 0;
logic signed [WIDTH-1:0] x_115 = 0;
logic signed [WIDTH-1:0] x_116 = 0;
logic signed [WIDTH-1:0] x_117 = 0;
logic signed [WIDTH-1:0] x_118 = 0;
logic signed [WIDTH-1:0] x_119 = 0;
logic signed [WIDTH-1:0] x_120 = 0;
logic signed [WIDTH-1:0] x_121 = 0;
logic signed [WIDTH-1:0] x_122 = 0;
logic signed [WIDTH-1:0] x_123 = 0;
logic signed [WIDTH-1:0] x_124 = 0;
logic signed [WIDTH-1:0] x_125 = 0;
logic signed [WIDTH-1:0] x_126 = 0;
logic signed [WIDTH-1:0] x_127 = 0;
logic signed [WIDTH-1:0] x_128 = 0;
logic signed [WIDTH-1:0] x_129 = 0;
logic signed [WIDTH-1:0] x_130 = 0;
logic signed [WIDTH-1:0] x_131 = 0;
logic signed [WIDTH-1:0] x_132 = 0;
logic signed [WIDTH-1:0] x_133 = 0;
logic signed [WIDTH-1:0] x_134 = 0;
logic signed [WIDTH-1:0] x_135 = 0;
logic signed [WIDTH-1:0] x_136 = 0;
logic signed [WIDTH-1:0] x_137 = 0;
logic signed [WIDTH-1:0] x_138 = 0;
logic signed [WIDTH-1:0] x_139 = 0;
logic signed [WIDTH-1:0] x_140 = 0;
logic signed [WIDTH-1:0] x_141 = 0;
logic signed [WIDTH-1:0] x_142 = 0;
logic signed [WIDTH-1:0] x_143 = 0;
logic signed [WIDTH-1:0] x_144 = 0;
logic signed [WIDTH-1:0] x_145 = 0;
logic signed [WIDTH-1:0] x_146 = 0;
logic signed [WIDTH-1:0] x_147 = 0;
logic signed [WIDTH-1:0] x_148 = 0;
logic signed [WIDTH-1:0] x_149 = 0;
logic signed [WIDTH-1:0] x_150 = 0;
logic signed [WIDTH-1:0] x_151 = 0;
logic signed [WIDTH-1:0] x_152 = 0;
logic signed [WIDTH-1:0] x_153 = 0;
logic signed [WIDTH-1:0] x_154 = 0;
logic signed [WIDTH-1:0] x_155 = 0;
logic signed [WIDTH-1:0] x_156 = 0;
logic signed [WIDTH-1:0] x_157 = 0;
logic signed [WIDTH-1:0] x_158 = 0;
logic signed [WIDTH-1:0] x_159 = 0;
logic signed [WIDTH-1:0] x_160 = 0;
logic signed [WIDTH-1:0] x_161 = 0;
logic signed [WIDTH-1:0] x_162 = 0;
logic signed [WIDTH-1:0] x_163 = 0;
logic signed [WIDTH-1:0] x_164 = 0;
logic signed [WIDTH-1:0] x_165 = 0;
logic signed [WIDTH-1:0] x_166 = 0;
logic signed [WIDTH-1:0] x_167 = 0;
logic signed [WIDTH-1:0] x_168 = 0;
logic signed [WIDTH-1:0] x_169 = 0;
logic signed [WIDTH-1:0] x_170 = 0;
logic signed [WIDTH-1:0] x_171 = 0;
logic signed [WIDTH-1:0] x_172 = 0;
logic signed [WIDTH-1:0] x_173 = 0;
logic signed [WIDTH-1:0] x_174 = 0;
logic signed [WIDTH-1:0] x_175 = 0;
logic signed [WIDTH-1:0] x_176 = 0;
logic signed [WIDTH-1:0] x_177 = 0;
logic signed [WIDTH-1:0] x_178 = 0;
logic signed [WIDTH-1:0] x_179 = 0;
logic signed [WIDTH-1:0] x_180 = 0;
logic signed [WIDTH-1:0] x_181 = 0;
logic signed [WIDTH-1:0] x_182 = 0;
logic signed [WIDTH-1:0] x_183 = 0;
logic signed [WIDTH-1:0] x_184 = 0;
logic signed [WIDTH-1:0] x_185 = 0;
logic signed [WIDTH-1:0] x_186 = 0;
logic signed [WIDTH-1:0] x_187 = 0;
logic signed [WIDTH-1:0] x_188 = 0;
logic signed [WIDTH-1:0] x_189 = 0;
logic signed [WIDTH-1:0] x_190 = 0;
logic signed [WIDTH-1:0] x_191 = 0;
logic signed [WIDTH-1:0] x_192 = 0;
logic signed [WIDTH-1:0] x_193 = 0;
logic signed [WIDTH-1:0] x_194 = 0;
logic signed [WIDTH-1:0] x_195 = 0;
logic signed [WIDTH-1:0] x_196 = 0;
logic signed [WIDTH-1:0] x_197 = 0;
logic signed [WIDTH-1:0] x_198 = 0;
logic signed [WIDTH-1:0] x_199 = 0;
logic signed [WIDTH-1:0] x_200 = 0;
logic signed [WIDTH-1:0] x_201 = 0;
logic signed [WIDTH-1:0] x_202 = 0;
logic signed [WIDTH-1:0] x_203 = 0;
logic signed [WIDTH-1:0] x_204 = 0;
logic signed [WIDTH-1:0] x_205 = 0;
logic signed [WIDTH-1:0] x_206 = 0;
logic signed [WIDTH-1:0] x_207 = 0;
logic signed [WIDTH-1:0] x_208 = 0;
logic signed [WIDTH-1:0] x_209 = 0;
logic signed [WIDTH-1:0] x_210 = 0;
logic signed [WIDTH-1:0] x_211 = 0;
logic signed [WIDTH-1:0] x_212 = 0;
logic signed [WIDTH-1:0] x_213 = 0;
logic signed [WIDTH-1:0] x_214 = 0;
logic signed [WIDTH-1:0] x_215 = 0;
logic signed [WIDTH-1:0] x_216 = 0;
logic signed [WIDTH-1:0] x_217 = 0;
logic signed [WIDTH-1:0] x_218 = 0;
logic signed [WIDTH-1:0] x_219 = 0;
logic signed [WIDTH-1:0] x_220 = 0;
logic signed [WIDTH-1:0] x_221 = 0;
logic signed [WIDTH-1:0] x_222 = 0;
logic signed [WIDTH-1:0] x_223 = 0;
logic signed [WIDTH-1:0] x_224 = 0;
logic signed [WIDTH-1:0] x_225 = 0;
logic signed [WIDTH-1:0] x_226 = 0;
logic signed [WIDTH-1:0] x_227 = 0;
logic signed [WIDTH-1:0] x_228 = 0;
logic signed [WIDTH-1:0] x_229 = 0;
logic signed [WIDTH-1:0] x_230 = 0;
logic signed [WIDTH-1:0] x_231 = 0;
logic signed [WIDTH-1:0] x_232 = 0;
logic signed [WIDTH-1:0] x_233 = 0;
logic signed [WIDTH-1:0] x_234 = 0;
logic signed [WIDTH-1:0] x_235 = 0;
logic signed [WIDTH-1:0] x_236 = 0;
logic signed [WIDTH-1:0] x_237 = 0;
logic signed [WIDTH-1:0] x_238 = 0;
logic signed [WIDTH-1:0] x_239 = 0;
logic signed [WIDTH-1:0] x_240 = 0;
logic signed [WIDTH-1:0] x_241 = 0;
logic signed [WIDTH-1:0] x_242 = 0;
logic signed [WIDTH-1:0] x_243 = 0;
logic signed [WIDTH-1:0] x_244 = 0;
logic signed [WIDTH-1:0] x_245 = 0;
logic signed [WIDTH-1:0] x_246 = 0;
logic signed [WIDTH-1:0] x_247 = 0;
logic signed [WIDTH-1:0] x_248 = 0;
logic signed [WIDTH-1:0] x_249 = 0;
logic signed [WIDTH-1:0] x_250 = 0;
logic signed [WIDTH-1:0] x_251 = 0;
logic signed [WIDTH-1:0] x_252 = 0;
logic signed [WIDTH-1:0] x_253 = 0;
logic signed [WIDTH-1:0] x_254 = 0;
logic signed [WIDTH-1:0] x_255 = 0;

logic signed [WIDTH-1:0] h_0 = 0;
logic signed [WIDTH-1:0] h_1 = 0;
logic signed [WIDTH-1:0] h_2 = 0;
logic signed [WIDTH-1:0] h_3 = 0;
logic signed [WIDTH-1:0] h_4 = 0;
logic signed [WIDTH-1:0] h_5 = 0;
logic signed [WIDTH-1:0] h_6 = 0;
logic signed [WIDTH-1:0] h_7 = 0;

// Input weights (h×d for each gate)
logic signed [WIDTH-1:0] w_ir_0_0 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_1 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_0_2 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_3 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_4 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_5 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_0_6 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_7 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_8 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_0_9 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_10 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_0_11 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_12 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_0_13 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_14 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_15 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_0_16 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_17 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_0_18 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_19 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_0_20 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_21 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_22 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_23 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_24 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_0_25 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_26 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_27 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_28 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_0_29 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_0_30 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_31 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_32 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_33 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_34 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_35 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_36 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_0_37 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_38 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_39 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_40 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_0_41 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_0_42 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_43 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_44 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_45 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_0_46 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_0_47 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_0_48 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_49 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_50 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_51 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_52 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_0_53 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_54 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_55 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_56 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_0_57 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_58 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_59 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_60 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_0_61 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_0_62 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_0_63 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_64 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_0_65 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_66 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_0_67 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_0_68 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_69 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_70 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_71 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_72 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_73 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_74 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_75 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_76 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_77 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_78 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_0_79 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_80 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_81 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_82 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_83 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_84 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_85 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_86 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_87 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_88 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_89 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_0_90 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_0_91 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_0_92 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_0_93 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_94 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_95 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_96 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_0_97 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_98 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_99 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_100 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_101 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_102 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_103 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_104 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_105 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_106 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_107 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_108 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_109 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_110 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_111 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_112 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_113 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_0_114 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_115 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_0_116 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_117 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_118 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_119 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_120 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_121 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_0_122 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_123 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_0_124 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_125 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_126 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_0_127 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_128 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_129 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_130 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_0_131 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_0_132 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_133 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_134 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_135 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_0_136 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_137 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_138 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_139 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_0_140 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_141 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_142 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_143 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_144 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_0_145 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_0_146 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_147 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_148 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_149 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_150 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_151 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_0_152 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_153 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_154 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_155 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_0_156 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_157 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_0_158 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_159 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_160 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_161 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_162 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_163 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_164 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_165 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_166 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_167 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_168 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_169 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_170 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_171 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_172 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_173 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_174 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_175 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_176 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_177 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_178 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_0_179 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_180 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_181 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_182 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_0_183 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_184 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_185 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_0_186 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_0_187 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_188 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_0_189 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_190 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_0_191 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_0_192 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_193 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_0_194 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_195 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_0_196 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_0_197 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_198 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_199 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_200 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_201 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_0_202 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_0_203 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_204 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_0_205 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_206 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_207 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_208 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_209 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_210 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_211 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_212 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_213 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_214 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_215 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_216 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_0_217 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_218 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_219 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_220 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_221 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_222 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_0_223 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_0_224 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_225 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_0_226 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_227 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_228 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_229 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_0_230 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_231 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_232 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_233 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_0_234 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_0_235 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_236 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_237 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_238 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_0_239 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_240 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_241 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_242 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_0_243 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_244 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_245 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_0_246 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_247 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_0_248 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_249 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_250 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_0_251 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_252 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_253 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_254 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_0_255 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_0 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_1 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_2 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_3 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_4 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_5 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_1_6 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_7 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_1_8 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_1_9 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_10 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_1_11 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_12 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_13 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_1_14 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_15 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_16 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_17 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_18 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_19 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_1_20 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_21 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_1_22 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_1_23 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_1_24 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_1_25 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_1_26 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_27 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_1_28 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_1_29 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_30 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_1_31 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_32 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_1_33 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_1_34 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_35 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_36 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_1_37 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_1_38 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_39 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_40 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_41 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_42 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_43 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_44 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_1_45 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_46 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_47 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_48 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_49 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_50 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_1_51 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_52 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_1_53 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_1_54 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_1_55 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_1_56 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_1_57 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_1_58 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_1_59 = 'b000001110;
logic signed [WIDTH-1:0] w_ir_1_60 = 'b000001010;
logic signed [WIDTH-1:0] w_ir_1_61 = 'b000001011;
logic signed [WIDTH-1:0] w_ir_1_62 = 'b000001101;
logic signed [WIDTH-1:0] w_ir_1_63 = 'b000001100;
logic signed [WIDTH-1:0] w_ir_1_64 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_65 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_66 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_67 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_68 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_69 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_1_70 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_1_71 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_1_72 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_1_73 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_74 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_75 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_76 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_77 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_78 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_79 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_80 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_1_81 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_1_82 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_83 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_1_84 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_85 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_86 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_1_87 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_88 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_89 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_90 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_91 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_1_92 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_93 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_94 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_95 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_1_96 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_97 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_1_98 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_99 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_1_100 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_101 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_1_102 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_1_103 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_1_104 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_105 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_106 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_107 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_108 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_109 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_110 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_111 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_1_112 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_113 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_114 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_115 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_116 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_117 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_118 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_119 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_120 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_121 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_1_122 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_123 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_124 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_1_125 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_1_126 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_127 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_1_128 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_1_129 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_130 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_1_131 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_132 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_1_133 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_134 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_1_135 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_1_136 = 'b000001011;
logic signed [WIDTH-1:0] w_ir_1_137 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_1_138 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_1_139 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_140 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_141 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_142 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_143 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_1_144 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_145 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_1_146 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_147 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_148 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_149 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_1_150 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_1_151 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_152 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_1_153 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_1_154 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_1_155 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_156 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_1_157 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_1_158 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_1_159 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_1_160 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_161 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_1_162 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_1_163 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_1_164 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_165 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_166 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_1_167 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_168 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_1_169 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_170 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_1_171 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_172 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_1_173 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_174 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_1_175 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_1_176 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_1_177 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_178 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_1_179 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_180 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_1_181 = 'b111110010;
logic signed [WIDTH-1:0] w_ir_1_182 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_183 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_184 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_1_185 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_186 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_1_187 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_1_188 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_189 = 'b111110100;
logic signed [WIDTH-1:0] w_ir_1_190 = 'b111110001;
logic signed [WIDTH-1:0] w_ir_1_191 = 'b111110000;
logic signed [WIDTH-1:0] w_ir_1_192 = 'b111110101;
logic signed [WIDTH-1:0] w_ir_1_193 = 'b111110101;
logic signed [WIDTH-1:0] w_ir_1_194 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_1_195 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_196 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_1_197 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_1_198 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_1_199 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_200 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_1_201 = 'b111110100;
logic signed [WIDTH-1:0] w_ir_1_202 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_203 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_1_204 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_1_205 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_1_206 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_1_207 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_208 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_209 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_210 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_211 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_1_212 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_213 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_214 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_1_215 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_216 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_1_217 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_1_218 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_1_219 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_220 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_1_221 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_1_222 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_1_223 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_1_224 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_1_225 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_226 = 'b111110100;
logic signed [WIDTH-1:0] w_ir_1_227 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_1_228 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_1_229 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_230 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_1_231 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_1_232 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_233 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_1_234 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_1_235 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_1_236 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_1_237 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_238 = 'b000010010;
logic signed [WIDTH-1:0] w_ir_1_239 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_1_240 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_241 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_1_242 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_1_243 = 'b000001100;
logic signed [WIDTH-1:0] w_ir_1_244 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_1_245 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_1_246 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_1_247 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_248 = 'b000010010;
logic signed [WIDTH-1:0] w_ir_1_249 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_250 = 'b000010011;
logic signed [WIDTH-1:0] w_ir_1_251 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_1_252 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_1_253 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_1_254 = 'b000001100;
logic signed [WIDTH-1:0] w_ir_1_255 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_2_0 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_2_1 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_2 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_3 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_4 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_5 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_6 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_2_7 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_2_8 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_9 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_2_10 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_11 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_2_12 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_13 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_14 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_15 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_16 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_17 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_2_18 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_2_19 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_20 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_21 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_22 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_2_23 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_24 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_25 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_26 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_2_27 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_28 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_29 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_30 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_2_31 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_32 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_33 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_2_34 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_2_35 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_2_36 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_2_37 = 'b111110110;
logic signed [WIDTH-1:0] w_ir_2_38 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_39 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_40 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_41 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_2_42 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_2_43 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_44 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_45 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_2_46 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_2_47 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_2_48 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_49 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_2_50 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_51 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_52 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_53 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_2_54 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_2_55 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_2_56 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_2_57 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_58 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_2_59 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_60 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_2_61 = 'b111110010;
logic signed [WIDTH-1:0] w_ir_2_62 = 'b111110000;
logic signed [WIDTH-1:0] w_ir_2_63 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_2_64 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_2_65 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_66 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_67 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_68 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_69 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_2_70 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_2_71 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_2_72 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_73 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_2_74 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_75 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_2_76 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_2_77 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_2_78 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_79 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_2_80 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_2_81 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_82 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_2_83 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_2_84 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_2_85 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_2_86 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_87 = 'b000001010;
logic signed [WIDTH-1:0] w_ir_2_88 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_89 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_2_90 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_2_91 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_2_92 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_2_93 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_2_94 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_95 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_2_96 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_2_97 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_98 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_2_99 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_2_100 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_2_101 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_102 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_103 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_2_104 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_2_105 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_2_106 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_2_107 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_2_108 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_109 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_2_110 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_111 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_112 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_2_113 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_114 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_2_115 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_116 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_2_117 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_2_118 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_2_119 = 'b000001010;
logic signed [WIDTH-1:0] w_ir_2_120 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_2_121 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_122 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_123 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_2_124 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_2_125 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_126 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_2_127 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_2_128 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_2_129 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_130 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_131 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_132 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_2_133 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_2_134 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_2_135 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_2_136 = 'b111110100;
logic signed [WIDTH-1:0] w_ir_2_137 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_138 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_139 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_2_140 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_2_141 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_2_142 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_143 = 'b111110101;
logic signed [WIDTH-1:0] w_ir_2_144 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_145 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_2_146 = 'b111110100;
logic signed [WIDTH-1:0] w_ir_2_147 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_2_148 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_2_149 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_2_150 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_2_151 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_2_152 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_2_153 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_2_154 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_2_155 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_156 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_2_157 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_2_158 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_159 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_160 = 'b000001011;
logic signed [WIDTH-1:0] w_ir_2_161 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_2_162 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_2_163 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_2_164 = 'b000001010;
logic signed [WIDTH-1:0] w_ir_2_165 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_2_166 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_2_167 = 'b111110101;
logic signed [WIDTH-1:0] w_ir_2_168 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_169 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_170 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_2_171 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_172 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_2_173 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_2_174 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_175 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_176 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_2_177 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_178 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_2_179 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_2_180 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_2_181 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_2_182 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_183 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_2_184 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_2_185 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_2_186 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_2_187 = 'b000001010;
logic signed [WIDTH-1:0] w_ir_2_188 = 'b000001111;
logic signed [WIDTH-1:0] w_ir_2_189 = 'b000001010;
logic signed [WIDTH-1:0] w_ir_2_190 = 'b000010001;
logic signed [WIDTH-1:0] w_ir_2_191 = 'b000001101;
logic signed [WIDTH-1:0] w_ir_2_192 = 'b111110101;
logic signed [WIDTH-1:0] w_ir_2_193 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_2_194 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_195 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_2_196 = 'b111110110;
logic signed [WIDTH-1:0] w_ir_2_197 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_198 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_2_199 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_2_200 = 'b111110010;
logic signed [WIDTH-1:0] w_ir_2_201 = 'b111110101;
logic signed [WIDTH-1:0] w_ir_2_202 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_2_203 = 'b111110101;
logic signed [WIDTH-1:0] w_ir_2_204 = 'b111110101;
logic signed [WIDTH-1:0] w_ir_2_205 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_2_206 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_207 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_208 = 'b000001011;
logic signed [WIDTH-1:0] w_ir_2_209 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_210 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_211 = 'b000001101;
logic signed [WIDTH-1:0] w_ir_2_212 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_213 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_2_214 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_2_215 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_2_216 = 'b111110110;
logic signed [WIDTH-1:0] w_ir_2_217 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_218 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_2_219 = 'b111110110;
logic signed [WIDTH-1:0] w_ir_2_220 = 'b000001101;
logic signed [WIDTH-1:0] w_ir_2_221 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_222 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_223 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_2_224 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_225 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_226 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_2_227 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_228 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_2_229 = 'b111110110;
logic signed [WIDTH-1:0] w_ir_2_230 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_231 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_232 = 'b111110100;
logic signed [WIDTH-1:0] w_ir_2_233 = 'b111110110;
logic signed [WIDTH-1:0] w_ir_2_234 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_2_235 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_236 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_2_237 = 'b000001100;
logic signed [WIDTH-1:0] w_ir_2_238 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_239 = 'b000001010;
logic signed [WIDTH-1:0] w_ir_2_240 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_241 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_242 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_2_243 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_2_244 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_245 = 'b111110110;
logic signed [WIDTH-1:0] w_ir_2_246 = 'b000001100;
logic signed [WIDTH-1:0] w_ir_2_247 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_248 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_2_249 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_2_250 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_2_251 = 'b000001011;
logic signed [WIDTH-1:0] w_ir_2_252 = 'b000001011;
logic signed [WIDTH-1:0] w_ir_2_253 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_2_254 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_255 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_3_0 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_3_1 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_3_2 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_3 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_4 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_5 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_3_6 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_7 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_8 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_3_9 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_10 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_3_11 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_12 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_3_13 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_14 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_15 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_3_16 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_17 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_3_18 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_19 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_3_20 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_21 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_22 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_3_23 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_3_24 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_3_25 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_26 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_27 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_3_28 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_3_29 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_3_30 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_31 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_3_32 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_33 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_34 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_35 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_36 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_3_37 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_3_38 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_39 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_40 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_3_41 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_3_42 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_43 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_44 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_45 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_46 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_3_47 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_3_48 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_49 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_50 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_51 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_52 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_3_53 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_54 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_55 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_56 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_3_57 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_58 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_59 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_60 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_3_61 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_3_62 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_3_63 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_64 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_65 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_66 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_3_67 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_3_68 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_69 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_70 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_71 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_72 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_73 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_74 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_75 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_76 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_77 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_78 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_3_79 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_80 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_81 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_82 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_83 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_84 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_85 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_86 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_87 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_88 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_89 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_3_90 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_3_91 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_3_92 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_3_93 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_94 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_95 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_96 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_97 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_98 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_99 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_100 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_101 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_102 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_103 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_104 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_105 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_106 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_107 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_108 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_109 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_110 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_111 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_112 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_113 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_3_114 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_115 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_3_116 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_117 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_118 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_119 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_120 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_121 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_3_122 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_123 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_124 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_125 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_126 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_3_127 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_128 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_129 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_130 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_3_131 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_132 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_133 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_134 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_135 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_3_136 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_137 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_138 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_139 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_3_140 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_141 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_142 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_143 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_3_144 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_3_145 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_3_146 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_147 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_148 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_149 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_150 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_151 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_3_152 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_3_153 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_154 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_155 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_3_156 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_157 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_3_158 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_159 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_160 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_161 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_3_162 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_163 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_164 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_165 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_166 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_167 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_168 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_169 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_170 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_171 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_172 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_173 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_174 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_175 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_176 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_177 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_178 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_179 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_3_180 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_3_181 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_182 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_3_183 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_184 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_185 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_3_186 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_187 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_188 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_3_189 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_190 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_3_191 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_3_192 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_193 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_3_194 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_195 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_3_196 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_3_197 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_198 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_199 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_200 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_201 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_3_202 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_203 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_204 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_205 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_206 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_207 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_208 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_209 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_210 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_211 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_212 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_213 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_214 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_3_215 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_216 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_3_217 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_218 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_219 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_220 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_221 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_222 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_223 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_3_224 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_225 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_3_226 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_227 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_228 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_229 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_3_230 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_3_231 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_232 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_233 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_3_234 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_3_235 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_236 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_237 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_238 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_3_239 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_240 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_241 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_242 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_243 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_244 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_245 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_246 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_247 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_3_248 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_249 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_250 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_251 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_252 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_253 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_254 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_3_255 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_4_0 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_1 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_4_2 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_3 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_4_4 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_5 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_4_6 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_4_7 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_4_8 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_4_9 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_4_10 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_4_11 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_4_12 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_13 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_4_14 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_4_15 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_16 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_4_17 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_4_18 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_4_19 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_4_20 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_21 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_4_22 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_4_23 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_4_24 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_4_25 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_4_26 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_27 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_4_28 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_4_29 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_30 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_4_31 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_4_32 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_4_33 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_4_34 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_4_35 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_4_36 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_4_37 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_4_38 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_4_39 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_4_40 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_4_41 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_4_42 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_43 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_4_44 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_4_45 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_46 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_47 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_48 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_49 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_4_50 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_4_51 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_4_52 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_4_53 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_4_54 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_4_55 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_4_56 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_4_57 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_4_58 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_4_59 = 'b000001110;
logic signed [WIDTH-1:0] w_ir_4_60 = 'b000001010;
logic signed [WIDTH-1:0] w_ir_4_61 = 'b000001011;
logic signed [WIDTH-1:0] w_ir_4_62 = 'b000001101;
logic signed [WIDTH-1:0] w_ir_4_63 = 'b000001100;
logic signed [WIDTH-1:0] w_ir_4_64 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_4_65 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_4_66 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_4_67 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_68 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_69 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_4_70 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_4_71 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_4_72 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_4_73 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_4_74 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_75 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_76 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_4_77 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_78 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_4_79 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_4_80 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_4_81 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_4_82 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_4_83 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_4_84 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_85 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_86 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_4_87 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_4_88 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_89 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_4_90 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_91 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_4_92 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_4_93 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_4_94 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_4_95 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_4_96 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_97 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_4_98 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_4_99 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_4_100 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_4_101 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_4_102 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_4_103 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_4_104 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_4_105 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_106 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_107 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_4_108 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_4_109 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_4_110 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_111 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_4_112 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_4_113 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_4_114 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_4_115 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_4_116 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_4_117 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_4_118 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_4_119 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_120 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_4_121 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_4_122 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_4_123 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_4_124 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_4_125 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_4_126 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_4_127 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_4_128 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_4_129 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_4_130 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_4_131 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_4_132 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_4_133 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_4_134 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_4_135 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_4_136 = 'b000001011;
logic signed [WIDTH-1:0] w_ir_4_137 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_4_138 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_4_139 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_140 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_141 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_4_142 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_4_143 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_4_144 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_4_145 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_4_146 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_147 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_148 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_149 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_4_150 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_4_151 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_152 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_4_153 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_4_154 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_4_155 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_4_156 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_4_157 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_4_158 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_4_159 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_4_160 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_161 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_4_162 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_4_163 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_4_164 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_165 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_4_166 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_4_167 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_168 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_4_169 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_4_170 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_4_171 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_4_172 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_4_173 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_4_174 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_4_175 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_4_176 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_4_177 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_4_178 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_4_179 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_180 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_4_181 = 'b111110010;
logic signed [WIDTH-1:0] w_ir_4_182 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_4_183 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_4_184 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_4_185 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_4_186 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_4_187 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_4_188 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_4_189 = 'b111110100;
logic signed [WIDTH-1:0] w_ir_4_190 = 'b111110001;
logic signed [WIDTH-1:0] w_ir_4_191 = 'b111110000;
logic signed [WIDTH-1:0] w_ir_4_192 = 'b111110101;
logic signed [WIDTH-1:0] w_ir_4_193 = 'b111110101;
logic signed [WIDTH-1:0] w_ir_4_194 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_4_195 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_4_196 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_4_197 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_4_198 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_4_199 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_4_200 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_4_201 = 'b111110100;
logic signed [WIDTH-1:0] w_ir_4_202 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_4_203 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_4_204 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_4_205 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_4_206 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_4_207 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_208 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_4_209 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_4_210 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_4_211 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_4_212 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_4_213 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_4_214 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_4_215 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_4_216 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_4_217 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_4_218 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_4_219 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_4_220 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_4_221 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_4_222 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_4_223 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_4_224 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_4_225 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_4_226 = 'b111110100;
logic signed [WIDTH-1:0] w_ir_4_227 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_4_228 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_4_229 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_230 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_4_231 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_4_232 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_4_233 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_4_234 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_4_235 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_4_236 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_4_237 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_4_238 = 'b000010010;
logic signed [WIDTH-1:0] w_ir_4_239 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_4_240 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_4_241 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_4_242 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_4_243 = 'b000001100;
logic signed [WIDTH-1:0] w_ir_4_244 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_4_245 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_4_246 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_4_247 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_4_248 = 'b000010010;
logic signed [WIDTH-1:0] w_ir_4_249 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_4_250 = 'b000010011;
logic signed [WIDTH-1:0] w_ir_4_251 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_4_252 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_4_253 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_4_254 = 'b000001100;
logic signed [WIDTH-1:0] w_ir_4_255 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_5_0 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_5_1 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_5_2 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_3 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_4 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_5_5 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_6 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_5_7 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_5_8 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_9 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_5_10 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_5_11 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_5_12 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_13 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_14 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_15 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_5_16 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_5_17 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_5_18 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_5_19 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_20 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_5_21 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_5_22 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_5_23 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_5_24 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_5_25 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_5_26 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_5_27 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_5_28 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_29 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_5_30 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_5_31 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_32 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_5_33 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_5_34 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_5_35 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_5_36 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_5_37 = 'b111110110;
logic signed [WIDTH-1:0] w_ir_5_38 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_5_39 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_5_40 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_5_41 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_5_42 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_5_43 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_44 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_5_45 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_5_46 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_5_47 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_5_48 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_5_49 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_5_50 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_5_51 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_5_52 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_53 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_5_54 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_5_55 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_5_56 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_5_57 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_58 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_5_59 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_60 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_5_61 = 'b111110010;
logic signed [WIDTH-1:0] w_ir_5_62 = 'b111110000;
logic signed [WIDTH-1:0] w_ir_5_63 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_5_64 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_5_65 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_5_66 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_5_67 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_5_68 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_5_69 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_5_70 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_5_71 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_5_72 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_5_73 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_5_74 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_75 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_5_76 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_5_77 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_5_78 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_79 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_5_80 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_5_81 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_82 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_5_83 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_5_84 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_5_85 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_5_86 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_87 = 'b000001010;
logic signed [WIDTH-1:0] w_ir_5_88 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_89 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_5_90 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_5_91 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_5_92 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_5_93 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_5_94 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_95 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_5_96 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_5_97 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_98 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_5_99 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_5_100 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_5_101 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_5_102 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_5_103 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_5_104 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_5_105 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_5_106 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_5_107 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_5_108 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_5_109 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_5_110 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_5_111 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_112 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_5_113 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_5_114 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_5_115 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_116 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_5_117 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_5_118 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_5_119 = 'b000001010;
logic signed [WIDTH-1:0] w_ir_5_120 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_5_121 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_122 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_5_123 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_5_124 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_5_125 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_5_126 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_5_127 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_5_128 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_5_129 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_130 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_5_131 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_5_132 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_5_133 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_5_134 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_5_135 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_5_136 = 'b111110100;
logic signed [WIDTH-1:0] w_ir_5_137 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_138 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_5_139 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_5_140 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_5_141 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_5_142 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_5_143 = 'b111110101;
logic signed [WIDTH-1:0] w_ir_5_144 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_145 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_5_146 = 'b111110100;
logic signed [WIDTH-1:0] w_ir_5_147 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_5_148 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_5_149 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_5_150 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_5_151 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_5_152 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_5_153 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_5_154 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_5_155 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_156 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_5_157 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_5_158 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_5_159 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_5_160 = 'b000001011;
logic signed [WIDTH-1:0] w_ir_5_161 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_5_162 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_5_163 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_5_164 = 'b000001010;
logic signed [WIDTH-1:0] w_ir_5_165 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_5_166 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_5_167 = 'b111110101;
logic signed [WIDTH-1:0] w_ir_5_168 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_169 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_5_170 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_5_171 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_5_172 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_5_173 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_5_174 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_175 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_176 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_5_177 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_5_178 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_5_179 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_5_180 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_5_181 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_5_182 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_5_183 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_5_184 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_5_185 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_5_186 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_5_187 = 'b000001010;
logic signed [WIDTH-1:0] w_ir_5_188 = 'b000001111;
logic signed [WIDTH-1:0] w_ir_5_189 = 'b000001010;
logic signed [WIDTH-1:0] w_ir_5_190 = 'b000010001;
logic signed [WIDTH-1:0] w_ir_5_191 = 'b000001101;
logic signed [WIDTH-1:0] w_ir_5_192 = 'b111110101;
logic signed [WIDTH-1:0] w_ir_5_193 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_5_194 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_5_195 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_5_196 = 'b111110110;
logic signed [WIDTH-1:0] w_ir_5_197 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_5_198 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_5_199 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_5_200 = 'b111110010;
logic signed [WIDTH-1:0] w_ir_5_201 = 'b111110101;
logic signed [WIDTH-1:0] w_ir_5_202 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_5_203 = 'b111110101;
logic signed [WIDTH-1:0] w_ir_5_204 = 'b111110101;
logic signed [WIDTH-1:0] w_ir_5_205 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_5_206 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_207 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_208 = 'b000001011;
logic signed [WIDTH-1:0] w_ir_5_209 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_210 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_5_211 = 'b000001101;
logic signed [WIDTH-1:0] w_ir_5_212 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_213 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_5_214 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_5_215 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_5_216 = 'b111110110;
logic signed [WIDTH-1:0] w_ir_5_217 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_218 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_5_219 = 'b111110110;
logic signed [WIDTH-1:0] w_ir_5_220 = 'b000001101;
logic signed [WIDTH-1:0] w_ir_5_221 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_222 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_5_223 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_5_224 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_225 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_226 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_5_227 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_228 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_5_229 = 'b111110110;
logic signed [WIDTH-1:0] w_ir_5_230 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_5_231 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_5_232 = 'b111110100;
logic signed [WIDTH-1:0] w_ir_5_233 = 'b111110110;
logic signed [WIDTH-1:0] w_ir_5_234 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_5_235 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_5_236 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_5_237 = 'b000001100;
logic signed [WIDTH-1:0] w_ir_5_238 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_5_239 = 'b000001010;
logic signed [WIDTH-1:0] w_ir_5_240 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_5_241 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_5_242 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_5_243 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_5_244 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_5_245 = 'b111110110;
logic signed [WIDTH-1:0] w_ir_5_246 = 'b000001100;
logic signed [WIDTH-1:0] w_ir_5_247 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_5_248 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_5_249 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_5_250 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_5_251 = 'b000001011;
logic signed [WIDTH-1:0] w_ir_5_252 = 'b000001011;
logic signed [WIDTH-1:0] w_ir_5_253 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_5_254 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_5_255 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_6_0 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_6_1 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_6_2 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_3 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_4 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_5 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_6_6 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_7 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_8 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_6_9 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_10 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_6_11 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_12 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_6_13 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_14 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_15 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_6_16 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_17 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_6_18 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_19 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_6_20 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_21 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_22 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_6_23 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_6_24 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_6_25 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_26 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_27 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_6_28 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_6_29 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_6_30 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_31 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_6_32 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_33 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_34 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_35 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_36 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_6_37 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_6_38 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_39 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_40 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_6_41 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_6_42 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_43 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_44 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_45 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_6_46 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_6_47 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_6_48 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_49 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_50 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_51 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_52 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_6_53 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_54 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_55 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_56 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_6_57 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_58 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_59 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_60 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_6_61 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_6_62 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_6_63 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_64 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_6_65 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_66 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_6_67 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_6_68 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_69 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_70 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_71 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_72 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_73 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_74 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_75 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_76 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_77 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_78 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_6_79 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_80 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_81 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_82 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_83 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_84 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_85 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_86 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_87 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_88 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_89 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_6_90 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_6_91 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_6_92 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_6_93 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_94 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_95 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_96 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_6_97 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_98 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_99 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_100 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_101 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_102 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_103 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_104 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_105 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_106 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_107 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_108 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_109 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_110 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_111 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_112 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_113 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_6_114 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_115 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_6_116 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_117 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_118 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_119 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_120 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_121 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_6_122 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_123 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_6_124 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_125 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_126 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_6_127 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_128 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_129 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_130 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_6_131 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_6_132 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_133 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_134 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_135 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_6_136 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_137 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_138 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_139 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_6_140 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_141 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_142 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_143 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_6_144 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_6_145 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_6_146 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_147 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_148 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_149 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_150 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_151 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_6_152 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_6_153 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_154 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_155 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_6_156 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_157 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_6_158 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_159 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_160 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_161 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_6_162 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_163 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_164 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_165 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_166 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_167 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_168 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_169 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_170 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_171 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_172 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_173 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_174 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_175 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_176 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_177 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_178 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_6_179 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_6_180 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_6_181 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_182 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_6_183 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_184 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_185 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_6_186 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_6_187 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_188 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_6_189 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_190 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_6_191 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_6_192 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_193 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_6_194 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_195 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_6_196 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_6_197 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_198 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_199 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_200 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_201 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_6_202 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_6_203 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_204 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_6_205 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_206 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_207 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_208 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_209 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_210 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_211 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_212 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_213 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_214 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_6_215 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_216 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_6_217 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_218 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_219 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_220 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_221 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_222 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_6_223 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_6_224 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_225 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_6_226 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_6_227 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_228 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_229 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_6_230 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_6_231 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_232 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_6_233 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_6_234 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_6_235 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_6_236 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_237 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_238 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_6_239 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_240 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_241 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_6_242 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_6_243 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_244 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_245 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_6_246 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_6_247 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_6_248 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_249 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_6_250 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_6_251 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_252 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_253 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_6_254 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_6_255 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_7_0 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_1 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_7_2 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_3 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_7_4 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_5 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_7_6 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_7_7 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_7_8 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_7_9 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_7_10 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_7_11 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_7_12 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_13 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_7_14 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_7_15 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_16 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_7_17 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_7_18 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_7_19 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_7_20 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_21 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_7_22 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_7_23 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_7_24 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_7_25 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_7_26 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_27 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_7_28 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_7_29 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_30 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_7_31 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_7_32 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_7_33 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_7_34 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_7_35 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_7_36 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_7_37 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_7_38 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_7_39 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_7_40 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_7_41 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_7_42 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_43 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_7_44 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_7_45 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_46 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_47 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_48 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_49 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_7_50 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_7_51 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_7_52 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_7_53 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_7_54 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_7_55 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_7_56 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_7_57 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_7_58 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_7_59 = 'b000001110;
logic signed [WIDTH-1:0] w_ir_7_60 = 'b000001010;
logic signed [WIDTH-1:0] w_ir_7_61 = 'b000001011;
logic signed [WIDTH-1:0] w_ir_7_62 = 'b000001101;
logic signed [WIDTH-1:0] w_ir_7_63 = 'b000001100;
logic signed [WIDTH-1:0] w_ir_7_64 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_7_65 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_7_66 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_7_67 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_68 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_69 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_7_70 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_7_71 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_7_72 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_7_73 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_7_74 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_75 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_76 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_7_77 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_78 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_7_79 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_7_80 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_7_81 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_7_82 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_7_83 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_7_84 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_85 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_86 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_7_87 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_7_88 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_89 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_7_90 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_91 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_7_92 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_7_93 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_7_94 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_7_95 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_7_96 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_97 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_7_98 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_7_99 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_7_100 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_7_101 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_7_102 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_7_103 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_7_104 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_7_105 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_106 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_107 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_7_108 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_7_109 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_7_110 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_111 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_7_112 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_7_113 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_7_114 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_7_115 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_7_116 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_7_117 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_7_118 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_7_119 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_120 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_7_121 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_7_122 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_7_123 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_7_124 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_7_125 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_7_126 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_7_127 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_7_128 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_7_129 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_7_130 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_7_131 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_7_132 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_7_133 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_7_134 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_7_135 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_7_136 = 'b000001011;
logic signed [WIDTH-1:0] w_ir_7_137 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_7_138 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_7_139 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_140 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_141 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_7_142 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_7_143 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_7_144 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_7_145 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_7_146 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_147 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_148 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_149 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_7_150 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_7_151 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_152 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_7_153 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_7_154 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_7_155 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_7_156 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_7_157 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_7_158 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_7_159 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_7_160 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_161 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_7_162 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_7_163 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_7_164 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_165 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_7_166 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_7_167 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_168 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_7_169 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_7_170 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_7_171 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_7_172 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_7_173 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_7_174 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_7_175 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_7_176 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_7_177 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_7_178 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_7_179 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_180 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_7_181 = 'b111110010;
logic signed [WIDTH-1:0] w_ir_7_182 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_7_183 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_7_184 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_7_185 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_7_186 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_7_187 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_7_188 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_7_189 = 'b111110100;
logic signed [WIDTH-1:0] w_ir_7_190 = 'b111110001;
logic signed [WIDTH-1:0] w_ir_7_191 = 'b111110000;
logic signed [WIDTH-1:0] w_ir_7_192 = 'b111110101;
logic signed [WIDTH-1:0] w_ir_7_193 = 'b111110101;
logic signed [WIDTH-1:0] w_ir_7_194 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_7_195 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_7_196 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_7_197 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_7_198 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_7_199 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_7_200 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_7_201 = 'b111110100;
logic signed [WIDTH-1:0] w_ir_7_202 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_7_203 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_7_204 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_7_205 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_7_206 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_7_207 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_208 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_7_209 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_7_210 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_7_211 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_7_212 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_7_213 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_7_214 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_7_215 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_7_216 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_7_217 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_7_218 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_7_219 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_7_220 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_7_221 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_7_222 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_7_223 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_7_224 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_7_225 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_7_226 = 'b111110100;
logic signed [WIDTH-1:0] w_ir_7_227 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_7_228 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_7_229 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_230 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_7_231 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_7_232 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_7_233 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_7_234 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_7_235 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_7_236 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_7_237 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_7_238 = 'b000010010;
logic signed [WIDTH-1:0] w_ir_7_239 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_7_240 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_7_241 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_7_242 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_7_243 = 'b000001100;
logic signed [WIDTH-1:0] w_ir_7_244 = 'b111110111;
logic signed [WIDTH-1:0] w_ir_7_245 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_7_246 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_7_247 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_7_248 = 'b000010010;
logic signed [WIDTH-1:0] w_ir_7_249 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_7_250 = 'b000010011;
logic signed [WIDTH-1:0] w_ir_7_251 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_7_252 = 'b111111000;
logic signed [WIDTH-1:0] w_ir_7_253 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_7_254 = 'b000001100;
logic signed [WIDTH-1:0] w_ir_7_255 = 'b111111000;

logic signed [WIDTH-1:0] w_iz_0_0 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_0_1 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_0_2 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_3 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_4 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_5 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_6 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_0_7 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_0_8 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_9 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_0_10 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_0_11 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_0_12 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_13 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_14 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_15 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_0_16 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_17 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_0_18 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_0_19 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_20 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_21 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_0_22 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_0_23 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_0_24 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_25 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_26 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_0_27 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_0_28 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_29 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_30 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_0_31 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_32 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_33 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_0_34 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_0_35 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_36 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_37 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_0_38 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_0_39 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_40 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_41 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_0_42 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_0_43 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_44 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_45 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_0_46 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_0_47 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_0_48 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_0_49 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_0_50 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_51 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_0_52 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_53 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_0_54 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_0_55 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_56 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_0_57 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_58 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_0_59 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_60 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_0_61 = 'b111110010;
logic signed [WIDTH-1:0] w_iz_0_62 = 'b111110000;
logic signed [WIDTH-1:0] w_iz_0_63 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_0_64 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_0_65 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_0_66 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_0_67 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_68 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_0_69 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_0_70 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_0_71 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_0_72 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_73 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_0_74 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_75 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_0_76 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_0_77 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_0_78 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_79 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_0_80 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_0_81 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_82 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_0_83 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_0_84 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_0_85 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_0_86 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_87 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_0_88 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_89 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_0_90 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_91 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_0_92 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_93 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_0_94 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_95 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_0_96 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_0_97 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_98 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_0_99 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_0_100 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_0_101 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_0_102 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_103 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_0_104 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_0_105 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_0_106 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_0_107 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_0_108 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_109 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_0_110 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_0_111 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_112 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_0_113 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_114 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_115 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_116 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_0_117 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_0_118 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_0_119 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_0_120 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_0_121 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_122 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_123 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_0_124 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_0_125 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_126 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_127 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_128 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_0_129 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_130 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_131 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_0_132 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_0_133 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_0_134 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_0_135 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_0_136 = 'b111110100;
logic signed [WIDTH-1:0] w_iz_0_137 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_138 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_139 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_0_140 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_0_141 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_0_142 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_143 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_0_144 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_145 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_0_146 = 'b111110100;
logic signed [WIDTH-1:0] w_iz_0_147 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_0_148 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_0_149 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_0_150 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_0_151 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_0_152 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_0_153 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_0_154 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_0_155 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_156 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_0_157 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_0_158 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_159 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_160 = 'b000001011;
logic signed [WIDTH-1:0] w_iz_0_161 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_0_162 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_0_163 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_0_164 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_0_165 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_0_166 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_0_167 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_0_168 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_169 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_170 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_0_171 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_0_172 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_173 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_0_174 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_175 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_176 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_177 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_178 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_0_179 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_180 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_0_181 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_0_182 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_183 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_0_184 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_185 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_0_186 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_0_187 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_0_188 = 'b000001111;
logic signed [WIDTH-1:0] w_iz_0_189 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_0_190 = 'b000010001;
logic signed [WIDTH-1:0] w_iz_0_191 = 'b000001101;
logic signed [WIDTH-1:0] w_iz_0_192 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_0_193 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_0_194 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_0_195 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_0_196 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_0_197 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_0_198 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_0_199 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_0_200 = 'b111110010;
logic signed [WIDTH-1:0] w_iz_0_201 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_0_202 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_0_203 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_0_204 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_0_205 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_0_206 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_207 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_208 = 'b000001011;
logic signed [WIDTH-1:0] w_iz_0_209 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_210 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_211 = 'b000001101;
logic signed [WIDTH-1:0] w_iz_0_212 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_213 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_0_214 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_215 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_0_216 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_0_217 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_218 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_0_219 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_0_220 = 'b000001101;
logic signed [WIDTH-1:0] w_iz_0_221 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_222 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_0_223 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_0_224 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_225 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_226 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_0_227 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_228 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_0_229 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_0_230 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_231 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_232 = 'b111110100;
logic signed [WIDTH-1:0] w_iz_0_233 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_0_234 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_0_235 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_0_236 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_0_237 = 'b000001100;
logic signed [WIDTH-1:0] w_iz_0_238 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_239 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_0_240 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_0_241 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_242 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_0_243 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_0_244 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_245 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_0_246 = 'b000001100;
logic signed [WIDTH-1:0] w_iz_0_247 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_0_248 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_0_249 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_0_250 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_0_251 = 'b000001011;
logic signed [WIDTH-1:0] w_iz_0_252 = 'b000001011;
logic signed [WIDTH-1:0] w_iz_0_253 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_0_254 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_0_255 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_1_0 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_1_1 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_1_2 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_3 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_4 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_5 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_1_6 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_7 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_8 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_1_9 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_10 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_1_11 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_12 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_1_13 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_14 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_15 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_1_16 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_17 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_1_18 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_19 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_1_20 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_21 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_22 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_1_23 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_1_24 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_1_25 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_26 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_27 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_1_28 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_1_29 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_1_30 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_31 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_1_32 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_33 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_34 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_35 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_36 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_1_37 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_1_38 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_39 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_40 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_1_41 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_1_42 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_43 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_44 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_45 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_46 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_1_47 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_1_48 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_49 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_50 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_51 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_52 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_1_53 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_54 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_55 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_56 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_1_57 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_58 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_59 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_60 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_1_61 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_1_62 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_1_63 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_64 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_65 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_66 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_1_67 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_1_68 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_69 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_70 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_71 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_72 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_73 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_74 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_75 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_76 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_77 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_78 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_1_79 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_80 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_81 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_82 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_83 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_84 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_85 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_86 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_87 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_88 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_89 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_1_90 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_1_91 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_1_92 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_1_93 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_94 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_95 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_96 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_97 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_98 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_99 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_100 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_101 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_102 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_103 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_104 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_105 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_106 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_107 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_108 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_109 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_110 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_111 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_112 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_113 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_1_114 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_115 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_1_116 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_117 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_118 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_119 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_120 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_121 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_1_122 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_123 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_124 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_125 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_126 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_1_127 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_128 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_129 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_130 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_1_131 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_132 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_133 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_134 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_135 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_1_136 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_137 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_138 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_139 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_1_140 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_141 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_142 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_143 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_1_144 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_1_145 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_1_146 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_147 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_148 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_149 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_150 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_151 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_1_152 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_1_153 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_154 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_155 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_1_156 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_157 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_1_158 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_159 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_160 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_161 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_1_162 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_163 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_164 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_165 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_166 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_167 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_168 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_169 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_170 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_171 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_172 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_173 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_174 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_175 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_176 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_177 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_178 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_179 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_1_180 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_1_181 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_182 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_1_183 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_184 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_185 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_1_186 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_187 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_188 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_1_189 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_190 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_1_191 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_1_192 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_193 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_1_194 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_195 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_1_196 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_1_197 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_198 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_199 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_200 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_201 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_1_202 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_203 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_204 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_205 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_206 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_207 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_208 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_209 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_210 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_211 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_212 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_213 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_214 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_1_215 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_216 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_1_217 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_218 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_219 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_220 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_221 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_222 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_223 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_1_224 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_225 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_1_226 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_227 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_228 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_229 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_1_230 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_1_231 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_232 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_233 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_1_234 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_1_235 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_236 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_237 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_238 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_1_239 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_240 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_241 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_242 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_243 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_244 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_245 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_246 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_247 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_1_248 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_249 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_250 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_251 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_252 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_253 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_254 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_1_255 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_0 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_1 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_2 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_3 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_4 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_5 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_2_6 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_7 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_8 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_2_9 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_10 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_2_11 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_12 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_13 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_2_14 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_2_15 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_16 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_17 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_18 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_19 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_20 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_21 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_2_22 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_2_23 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_2_24 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_2_25 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_2_26 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_27 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_2_28 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_2_29 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_30 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_2_31 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_32 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_2_33 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_2_34 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_35 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_36 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_2_37 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_38 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_39 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_2_40 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_2_41 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_42 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_43 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_44 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_2_45 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_46 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_47 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_48 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_49 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_50 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_2_51 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_52 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_2_53 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_2_54 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_2_55 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_2_56 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_2_57 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_2_58 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_2_59 = 'b000001110;
logic signed [WIDTH-1:0] w_iz_2_60 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_2_61 = 'b000001011;
logic signed [WIDTH-1:0] w_iz_2_62 = 'b000001101;
logic signed [WIDTH-1:0] w_iz_2_63 = 'b000001100;
logic signed [WIDTH-1:0] w_iz_2_64 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_2_65 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_2_66 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_2_67 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_68 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_69 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_70 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_2_71 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_2_72 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_2_73 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_74 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_75 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_76 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_77 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_78 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_79 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_80 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_2_81 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_82 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_2_83 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_2_84 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_85 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_86 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_2_87 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_2_88 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_89 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_90 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_91 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_2_92 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_2_93 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_94 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_95 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_2_96 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_97 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_2_98 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_99 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_2_100 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_101 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_2_102 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_2_103 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_2_104 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_105 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_106 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_107 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_108 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_2_109 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_110 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_111 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_2_112 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_2_113 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_2_114 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_2_115 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_2_116 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_117 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_118 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_2_119 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_120 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_2_121 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_122 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_123 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_124 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_2_125 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_2_126 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_127 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_2_128 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_2_129 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_130 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_2_131 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_132 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_2_133 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_2_134 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_2_135 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_2_136 = 'b000001011;
logic signed [WIDTH-1:0] w_iz_2_137 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_2_138 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_2_139 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_140 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_141 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_2_142 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_143 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_2_144 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_145 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_2_146 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_147 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_148 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_149 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_150 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_2_151 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_152 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_153 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_2_154 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_2_155 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_156 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_2_157 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_2_158 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_159 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_2_160 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_161 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_2_162 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_2_163 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_2_164 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_165 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_2_166 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_2_167 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_168 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_2_169 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_170 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_2_171 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_2_172 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_2_173 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_174 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_2_175 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_2_176 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_2_177 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_178 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_2_179 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_180 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_2_181 = 'b111110010;
logic signed [WIDTH-1:0] w_iz_2_182 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_183 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_2_184 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_185 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_186 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_187 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_2_188 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_189 = 'b111110100;
logic signed [WIDTH-1:0] w_iz_2_190 = 'b111110001;
logic signed [WIDTH-1:0] w_iz_2_191 = 'b111110000;
logic signed [WIDTH-1:0] w_iz_2_192 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_2_193 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_2_194 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_2_195 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_196 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_2_197 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_2_198 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_2_199 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_2_200 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_201 = 'b111110100;
logic signed [WIDTH-1:0] w_iz_2_202 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_203 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_2_204 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_2_205 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_2_206 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_2_207 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_208 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_2_209 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_210 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_2_211 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_2_212 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_213 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_214 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_2_215 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_216 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_2_217 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_2_218 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_2_219 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_220 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_2_221 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_2_222 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_2_223 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_2_224 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_225 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_226 = 'b111110100;
logic signed [WIDTH-1:0] w_iz_2_227 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_2_228 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_2_229 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_230 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_2_231 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_2_232 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_233 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_2_234 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_2_235 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_2_236 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_237 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_2_238 = 'b000010010;
logic signed [WIDTH-1:0] w_iz_2_239 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_240 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_241 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_242 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_2_243 = 'b000001100;
logic signed [WIDTH-1:0] w_iz_2_244 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_2_245 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_2_246 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_2_247 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_2_248 = 'b000010010;
logic signed [WIDTH-1:0] w_iz_2_249 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_2_250 = 'b000010011;
logic signed [WIDTH-1:0] w_iz_2_251 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_2_252 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_2_253 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_2_254 = 'b000001100;
logic signed [WIDTH-1:0] w_iz_2_255 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_3_0 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_3_1 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_3_2 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_3 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_4 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_3_5 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_6 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_3_7 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_3_8 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_9 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_3_10 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_3_11 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_3_12 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_13 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_14 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_15 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_3_16 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_3_17 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_3_18 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_3_19 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_20 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_3_21 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_3_22 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_3_23 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_3_24 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_3_25 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_3_26 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_3_27 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_3_28 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_29 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_3_30 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_3_31 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_32 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_3_33 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_3_34 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_3_35 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_3_36 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_3_37 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_3_38 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_3_39 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_3_40 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_3_41 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_3_42 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_3_43 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_44 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_3_45 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_3_46 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_3_47 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_3_48 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_3_49 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_3_50 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_3_51 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_3_52 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_53 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_3_54 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_3_55 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_3_56 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_3_57 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_58 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_3_59 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_60 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_3_61 = 'b111110010;
logic signed [WIDTH-1:0] w_iz_3_62 = 'b111110000;
logic signed [WIDTH-1:0] w_iz_3_63 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_3_64 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_3_65 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_3_66 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_3_67 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_3_68 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_3_69 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_3_70 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_3_71 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_3_72 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_3_73 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_3_74 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_75 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_3_76 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_3_77 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_3_78 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_79 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_3_80 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_3_81 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_82 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_3_83 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_3_84 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_3_85 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_3_86 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_87 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_3_88 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_89 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_3_90 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_3_91 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_3_92 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_3_93 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_3_94 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_95 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_3_96 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_3_97 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_98 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_3_99 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_3_100 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_3_101 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_3_102 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_3_103 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_3_104 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_3_105 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_3_106 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_3_107 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_3_108 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_3_109 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_3_110 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_3_111 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_112 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_3_113 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_3_114 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_3_115 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_116 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_3_117 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_3_118 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_3_119 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_3_120 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_3_121 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_122 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_3_123 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_3_124 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_3_125 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_3_126 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_3_127 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_3_128 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_3_129 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_130 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_3_131 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_3_132 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_3_133 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_3_134 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_3_135 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_3_136 = 'b111110100;
logic signed [WIDTH-1:0] w_iz_3_137 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_138 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_3_139 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_3_140 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_3_141 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_3_142 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_3_143 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_3_144 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_145 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_3_146 = 'b111110100;
logic signed [WIDTH-1:0] w_iz_3_147 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_3_148 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_3_149 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_3_150 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_3_151 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_3_152 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_3_153 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_3_154 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_3_155 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_156 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_3_157 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_3_158 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_3_159 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_3_160 = 'b000001011;
logic signed [WIDTH-1:0] w_iz_3_161 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_3_162 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_3_163 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_3_164 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_3_165 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_3_166 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_3_167 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_3_168 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_169 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_3_170 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_3_171 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_3_172 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_3_173 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_3_174 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_175 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_176 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_3_177 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_3_178 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_3_179 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_3_180 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_3_181 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_3_182 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_3_183 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_3_184 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_3_185 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_3_186 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_3_187 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_3_188 = 'b000001111;
logic signed [WIDTH-1:0] w_iz_3_189 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_3_190 = 'b000010001;
logic signed [WIDTH-1:0] w_iz_3_191 = 'b000001101;
logic signed [WIDTH-1:0] w_iz_3_192 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_3_193 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_3_194 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_3_195 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_3_196 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_3_197 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_3_198 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_3_199 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_3_200 = 'b111110010;
logic signed [WIDTH-1:0] w_iz_3_201 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_3_202 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_3_203 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_3_204 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_3_205 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_3_206 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_207 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_208 = 'b000001011;
logic signed [WIDTH-1:0] w_iz_3_209 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_210 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_3_211 = 'b000001101;
logic signed [WIDTH-1:0] w_iz_3_212 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_213 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_3_214 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_3_215 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_3_216 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_3_217 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_218 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_3_219 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_3_220 = 'b000001101;
logic signed [WIDTH-1:0] w_iz_3_221 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_222 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_3_223 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_3_224 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_225 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_226 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_3_227 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_228 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_3_229 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_3_230 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_231 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_3_232 = 'b111110100;
logic signed [WIDTH-1:0] w_iz_3_233 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_3_234 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_3_235 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_3_236 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_3_237 = 'b000001100;
logic signed [WIDTH-1:0] w_iz_3_238 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_3_239 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_3_240 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_3_241 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_3_242 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_3_243 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_3_244 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_245 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_3_246 = 'b000001100;
logic signed [WIDTH-1:0] w_iz_3_247 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_3_248 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_3_249 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_3_250 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_3_251 = 'b000001011;
logic signed [WIDTH-1:0] w_iz_3_252 = 'b000001011;
logic signed [WIDTH-1:0] w_iz_3_253 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_3_254 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_3_255 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_4_0 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_4_1 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_4_2 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_3 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_4 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_5 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_4_6 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_7 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_8 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_4_9 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_10 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_4_11 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_12 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_4_13 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_14 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_15 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_4_16 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_17 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_4_18 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_19 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_4_20 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_21 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_22 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_4_23 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_4_24 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_4_25 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_26 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_27 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_4_28 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_4_29 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_4_30 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_31 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_4_32 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_33 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_34 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_35 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_36 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_4_37 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_4_38 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_39 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_40 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_4_41 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_4_42 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_43 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_44 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_45 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_4_46 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_4_47 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_4_48 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_49 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_50 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_51 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_52 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_4_53 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_54 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_55 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_56 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_4_57 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_58 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_59 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_60 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_4_61 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_4_62 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_4_63 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_64 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_4_65 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_66 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_4_67 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_4_68 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_69 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_70 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_71 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_72 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_73 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_74 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_75 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_76 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_77 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_78 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_4_79 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_80 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_81 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_82 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_83 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_84 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_85 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_86 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_87 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_88 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_89 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_4_90 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_4_91 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_4_92 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_4_93 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_94 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_95 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_96 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_4_97 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_98 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_99 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_100 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_101 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_102 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_103 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_104 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_105 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_106 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_107 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_108 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_109 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_110 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_111 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_112 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_113 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_4_114 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_115 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_4_116 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_117 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_118 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_119 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_120 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_121 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_4_122 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_123 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_4_124 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_125 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_126 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_4_127 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_128 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_129 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_130 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_4_131 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_4_132 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_133 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_134 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_135 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_4_136 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_137 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_138 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_139 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_4_140 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_141 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_142 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_143 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_4_144 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_4_145 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_4_146 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_147 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_148 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_149 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_150 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_151 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_4_152 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_4_153 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_154 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_155 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_4_156 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_157 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_4_158 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_159 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_160 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_161 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_4_162 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_163 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_164 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_165 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_166 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_167 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_168 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_169 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_170 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_171 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_172 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_173 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_174 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_175 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_176 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_177 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_178 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_4_179 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_4_180 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_4_181 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_182 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_4_183 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_184 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_185 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_4_186 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_4_187 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_188 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_4_189 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_190 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_4_191 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_4_192 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_193 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_4_194 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_195 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_4_196 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_4_197 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_198 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_199 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_200 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_201 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_4_202 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_4_203 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_204 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_4_205 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_206 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_207 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_208 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_209 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_210 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_211 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_212 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_213 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_214 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_4_215 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_216 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_4_217 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_218 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_219 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_220 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_221 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_222 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_4_223 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_4_224 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_225 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_4_226 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_4_227 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_228 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_229 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_4_230 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_4_231 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_232 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_4_233 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_4_234 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_4_235 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_4_236 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_237 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_238 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_4_239 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_240 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_241 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_4_242 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_4_243 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_244 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_245 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_4_246 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_4_247 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_4_248 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_249 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_4_250 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_4_251 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_252 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_253 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_4_254 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_4_255 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_5_0 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_1 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_5_2 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_3 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_5_4 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_5 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_5_6 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_5_7 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_5_8 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_5_9 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_5_10 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_5_11 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_5_12 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_13 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_5_14 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_5_15 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_16 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_5_17 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_5_18 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_5_19 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_5_20 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_21 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_5_22 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_5_23 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_5_24 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_5_25 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_5_26 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_27 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_5_28 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_5_29 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_30 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_5_31 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_5_32 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_5_33 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_5_34 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_5_35 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_5_36 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_5_37 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_5_38 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_5_39 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_5_40 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_5_41 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_5_42 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_43 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_5_44 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_5_45 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_46 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_47 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_48 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_49 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_5_50 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_5_51 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_5_52 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_5_53 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_5_54 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_5_55 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_5_56 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_5_57 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_5_58 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_5_59 = 'b000001110;
logic signed [WIDTH-1:0] w_iz_5_60 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_5_61 = 'b000001011;
logic signed [WIDTH-1:0] w_iz_5_62 = 'b000001101;
logic signed [WIDTH-1:0] w_iz_5_63 = 'b000001100;
logic signed [WIDTH-1:0] w_iz_5_64 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_5_65 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_5_66 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_5_67 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_68 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_69 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_5_70 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_5_71 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_5_72 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_5_73 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_5_74 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_75 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_76 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_5_77 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_78 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_5_79 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_5_80 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_5_81 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_5_82 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_5_83 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_5_84 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_85 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_86 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_5_87 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_5_88 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_89 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_5_90 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_91 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_5_92 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_5_93 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_5_94 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_5_95 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_5_96 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_97 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_5_98 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_5_99 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_5_100 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_5_101 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_5_102 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_5_103 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_5_104 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_5_105 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_106 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_107 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_5_108 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_5_109 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_5_110 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_111 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_5_112 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_5_113 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_5_114 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_5_115 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_5_116 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_5_117 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_5_118 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_5_119 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_120 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_5_121 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_5_122 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_5_123 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_5_124 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_5_125 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_5_126 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_5_127 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_5_128 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_5_129 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_5_130 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_5_131 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_5_132 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_5_133 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_5_134 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_5_135 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_5_136 = 'b000001011;
logic signed [WIDTH-1:0] w_iz_5_137 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_5_138 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_5_139 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_140 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_141 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_5_142 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_5_143 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_5_144 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_5_145 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_5_146 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_147 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_148 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_149 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_5_150 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_5_151 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_152 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_5_153 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_5_154 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_5_155 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_5_156 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_5_157 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_5_158 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_5_159 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_5_160 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_161 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_5_162 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_5_163 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_5_164 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_165 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_5_166 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_5_167 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_168 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_5_169 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_5_170 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_5_171 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_5_172 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_5_173 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_5_174 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_5_175 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_5_176 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_5_177 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_5_178 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_5_179 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_180 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_5_181 = 'b111110010;
logic signed [WIDTH-1:0] w_iz_5_182 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_5_183 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_5_184 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_5_185 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_5_186 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_5_187 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_5_188 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_5_189 = 'b111110100;
logic signed [WIDTH-1:0] w_iz_5_190 = 'b111110001;
logic signed [WIDTH-1:0] w_iz_5_191 = 'b111110000;
logic signed [WIDTH-1:0] w_iz_5_192 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_5_193 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_5_194 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_5_195 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_5_196 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_5_197 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_5_198 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_5_199 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_5_200 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_5_201 = 'b111110100;
logic signed [WIDTH-1:0] w_iz_5_202 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_5_203 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_5_204 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_5_205 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_5_206 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_5_207 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_208 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_5_209 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_5_210 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_5_211 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_5_212 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_5_213 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_5_214 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_5_215 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_5_216 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_5_217 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_5_218 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_5_219 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_5_220 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_5_221 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_5_222 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_5_223 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_5_224 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_5_225 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_5_226 = 'b111110100;
logic signed [WIDTH-1:0] w_iz_5_227 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_5_228 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_5_229 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_230 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_5_231 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_5_232 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_5_233 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_5_234 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_5_235 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_5_236 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_5_237 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_5_238 = 'b000010010;
logic signed [WIDTH-1:0] w_iz_5_239 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_5_240 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_5_241 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_5_242 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_5_243 = 'b000001100;
logic signed [WIDTH-1:0] w_iz_5_244 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_5_245 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_5_246 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_5_247 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_5_248 = 'b000010010;
logic signed [WIDTH-1:0] w_iz_5_249 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_5_250 = 'b000010011;
logic signed [WIDTH-1:0] w_iz_5_251 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_5_252 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_5_253 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_5_254 = 'b000001100;
logic signed [WIDTH-1:0] w_iz_5_255 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_6_0 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_6_1 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_6_2 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_3 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_4 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_6_5 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_6 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_6_7 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_6_8 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_9 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_6_10 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_6_11 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_6_12 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_13 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_14 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_15 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_6_16 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_6_17 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_6_18 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_6_19 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_20 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_6_21 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_6_22 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_6_23 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_6_24 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_6_25 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_6_26 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_6_27 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_6_28 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_29 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_6_30 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_6_31 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_32 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_6_33 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_6_34 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_6_35 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_6_36 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_6_37 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_6_38 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_6_39 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_6_40 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_6_41 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_6_42 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_6_43 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_44 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_6_45 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_6_46 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_6_47 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_6_48 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_6_49 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_6_50 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_6_51 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_6_52 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_53 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_6_54 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_6_55 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_6_56 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_6_57 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_58 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_6_59 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_60 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_6_61 = 'b111110010;
logic signed [WIDTH-1:0] w_iz_6_62 = 'b111110000;
logic signed [WIDTH-1:0] w_iz_6_63 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_6_64 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_6_65 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_6_66 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_6_67 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_6_68 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_6_69 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_6_70 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_6_71 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_6_72 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_6_73 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_6_74 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_75 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_6_76 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_6_77 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_6_78 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_79 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_6_80 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_6_81 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_82 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_6_83 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_6_84 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_6_85 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_6_86 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_87 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_6_88 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_89 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_6_90 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_6_91 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_6_92 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_6_93 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_6_94 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_95 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_6_96 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_6_97 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_98 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_6_99 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_6_100 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_6_101 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_6_102 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_6_103 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_6_104 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_6_105 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_6_106 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_6_107 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_6_108 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_6_109 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_6_110 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_6_111 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_112 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_6_113 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_6_114 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_6_115 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_116 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_6_117 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_6_118 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_6_119 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_6_120 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_6_121 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_122 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_6_123 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_6_124 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_6_125 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_6_126 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_6_127 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_6_128 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_6_129 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_130 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_6_131 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_6_132 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_6_133 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_6_134 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_6_135 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_6_136 = 'b111110100;
logic signed [WIDTH-1:0] w_iz_6_137 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_138 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_6_139 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_6_140 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_6_141 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_6_142 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_6_143 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_6_144 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_145 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_6_146 = 'b111110100;
logic signed [WIDTH-1:0] w_iz_6_147 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_6_148 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_6_149 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_6_150 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_6_151 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_6_152 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_6_153 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_6_154 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_6_155 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_156 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_6_157 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_6_158 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_6_159 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_6_160 = 'b000001011;
logic signed [WIDTH-1:0] w_iz_6_161 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_6_162 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_6_163 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_6_164 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_6_165 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_6_166 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_6_167 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_6_168 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_169 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_6_170 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_6_171 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_6_172 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_6_173 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_6_174 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_175 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_176 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_6_177 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_6_178 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_6_179 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_6_180 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_6_181 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_6_182 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_6_183 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_6_184 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_6_185 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_6_186 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_6_187 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_6_188 = 'b000001111;
logic signed [WIDTH-1:0] w_iz_6_189 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_6_190 = 'b000010001;
logic signed [WIDTH-1:0] w_iz_6_191 = 'b000001101;
logic signed [WIDTH-1:0] w_iz_6_192 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_6_193 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_6_194 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_6_195 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_6_196 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_6_197 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_6_198 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_6_199 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_6_200 = 'b111110010;
logic signed [WIDTH-1:0] w_iz_6_201 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_6_202 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_6_203 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_6_204 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_6_205 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_6_206 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_207 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_208 = 'b000001011;
logic signed [WIDTH-1:0] w_iz_6_209 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_210 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_6_211 = 'b000001101;
logic signed [WIDTH-1:0] w_iz_6_212 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_213 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_6_214 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_6_215 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_6_216 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_6_217 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_218 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_6_219 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_6_220 = 'b000001101;
logic signed [WIDTH-1:0] w_iz_6_221 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_222 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_6_223 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_6_224 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_225 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_226 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_6_227 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_228 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_6_229 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_6_230 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_6_231 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_6_232 = 'b111110100;
logic signed [WIDTH-1:0] w_iz_6_233 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_6_234 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_6_235 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_6_236 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_6_237 = 'b000001100;
logic signed [WIDTH-1:0] w_iz_6_238 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_6_239 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_6_240 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_6_241 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_6_242 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_6_243 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_6_244 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_6_245 = 'b111110110;
logic signed [WIDTH-1:0] w_iz_6_246 = 'b000001100;
logic signed [WIDTH-1:0] w_iz_6_247 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_6_248 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_6_249 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_6_250 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_6_251 = 'b000001011;
logic signed [WIDTH-1:0] w_iz_6_252 = 'b000001011;
logic signed [WIDTH-1:0] w_iz_6_253 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_6_254 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_6_255 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_7_0 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_7_1 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_7_2 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_3 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_4 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_5 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_7_6 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_7 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_8 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_7_9 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_10 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_7_11 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_12 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_7_13 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_14 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_15 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_7_16 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_17 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_7_18 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_19 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_7_20 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_21 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_22 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_7_23 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_7_24 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_7_25 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_26 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_27 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_7_28 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_7_29 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_7_30 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_31 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_7_32 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_33 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_34 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_35 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_36 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_7_37 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_7_38 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_39 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_40 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_7_41 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_7_42 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_43 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_44 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_45 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_7_46 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_7_47 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_7_48 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_49 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_50 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_51 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_52 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_7_53 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_54 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_55 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_56 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_7_57 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_58 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_59 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_60 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_7_61 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_7_62 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_7_63 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_64 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_7_65 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_66 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_7_67 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_7_68 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_69 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_70 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_71 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_72 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_73 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_74 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_75 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_76 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_77 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_78 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_7_79 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_80 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_81 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_82 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_83 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_84 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_85 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_86 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_87 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_88 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_89 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_7_90 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_7_91 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_7_92 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_7_93 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_94 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_95 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_96 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_7_97 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_98 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_99 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_100 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_101 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_102 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_103 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_104 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_105 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_106 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_107 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_108 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_109 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_110 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_111 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_112 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_113 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_7_114 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_115 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_7_116 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_117 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_118 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_119 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_120 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_121 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_7_122 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_123 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_7_124 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_125 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_126 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_7_127 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_128 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_129 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_130 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_7_131 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_7_132 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_133 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_134 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_135 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_7_136 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_137 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_138 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_139 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_7_140 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_141 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_142 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_143 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_7_144 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_7_145 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_7_146 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_147 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_148 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_149 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_150 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_151 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_7_152 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_7_153 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_154 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_155 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_7_156 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_157 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_7_158 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_159 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_160 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_161 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_7_162 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_163 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_164 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_165 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_166 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_167 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_168 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_169 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_170 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_171 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_172 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_173 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_174 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_175 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_176 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_177 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_178 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_7_179 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_7_180 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_7_181 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_182 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_7_183 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_184 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_185 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_7_186 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_7_187 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_188 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_7_189 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_190 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_7_191 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_7_192 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_193 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_7_194 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_195 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_7_196 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_7_197 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_198 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_199 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_200 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_201 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_7_202 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_7_203 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_204 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_7_205 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_206 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_207 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_208 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_209 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_210 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_211 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_212 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_213 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_214 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_7_215 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_216 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_7_217 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_218 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_219 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_220 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_221 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_222 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_7_223 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_7_224 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_225 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_7_226 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_7_227 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_228 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_229 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_7_230 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_7_231 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_232 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_7_233 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_7_234 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_7_235 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_7_236 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_237 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_238 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_7_239 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_240 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_241 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_7_242 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_7_243 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_244 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_245 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_7_246 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_7_247 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_7_248 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_249 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_7_250 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_7_251 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_252 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_253 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_7_254 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_7_255 = 'b111111110;

logic signed [WIDTH-1:0] w_in_0_0 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_1 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_2 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_3 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_4 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_5 = 'b000000011;
logic signed [WIDTH-1:0] w_in_0_6 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_7 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_8 = 'b111111001;
logic signed [WIDTH-1:0] w_in_0_9 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_10 = 'b111111001;
logic signed [WIDTH-1:0] w_in_0_11 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_12 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_13 = 'b000000011;
logic signed [WIDTH-1:0] w_in_0_14 = 'b000000001;
logic signed [WIDTH-1:0] w_in_0_15 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_16 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_17 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_18 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_19 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_20 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_21 = 'b000000011;
logic signed [WIDTH-1:0] w_in_0_22 = 'b000001000;
logic signed [WIDTH-1:0] w_in_0_23 = 'b000000101;
logic signed [WIDTH-1:0] w_in_0_24 = 'b111111001;
logic signed [WIDTH-1:0] w_in_0_25 = 'b111111010;
logic signed [WIDTH-1:0] w_in_0_26 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_27 = 'b111111001;
logic signed [WIDTH-1:0] w_in_0_28 = 'b000000110;
logic signed [WIDTH-1:0] w_in_0_29 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_30 = 'b000000110;
logic signed [WIDTH-1:0] w_in_0_31 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_32 = 'b111111001;
logic signed [WIDTH-1:0] w_in_0_33 = 'b111111010;
logic signed [WIDTH-1:0] w_in_0_34 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_35 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_36 = 'b111111010;
logic signed [WIDTH-1:0] w_in_0_37 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_38 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_39 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_40 = 'b000000001;
logic signed [WIDTH-1:0] w_in_0_41 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_42 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_43 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_44 = 'b111111000;
logic signed [WIDTH-1:0] w_in_0_45 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_46 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_47 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_48 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_49 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_50 = 'b000000101;
logic signed [WIDTH-1:0] w_in_0_51 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_52 = 'b000000111;
logic signed [WIDTH-1:0] w_in_0_53 = 'b000000100;
logic signed [WIDTH-1:0] w_in_0_54 = 'b000001000;
logic signed [WIDTH-1:0] w_in_0_55 = 'b000000110;
logic signed [WIDTH-1:0] w_in_0_56 = 'b000000011;
logic signed [WIDTH-1:0] w_in_0_57 = 'b111111001;
logic signed [WIDTH-1:0] w_in_0_58 = 'b000000100;
logic signed [WIDTH-1:0] w_in_0_59 = 'b000001110;
logic signed [WIDTH-1:0] w_in_0_60 = 'b000001010;
logic signed [WIDTH-1:0] w_in_0_61 = 'b000001011;
logic signed [WIDTH-1:0] w_in_0_62 = 'b000001101;
logic signed [WIDTH-1:0] w_in_0_63 = 'b000001100;
logic signed [WIDTH-1:0] w_in_0_64 = 'b000000001;
logic signed [WIDTH-1:0] w_in_0_65 = 'b000000001;
logic signed [WIDTH-1:0] w_in_0_66 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_67 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_68 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_69 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_70 = 'b000000110;
logic signed [WIDTH-1:0] w_in_0_71 = 'b111111001;
logic signed [WIDTH-1:0] w_in_0_72 = 'b111111010;
logic signed [WIDTH-1:0] w_in_0_73 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_74 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_75 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_76 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_77 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_78 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_79 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_80 = 'b000000101;
logic signed [WIDTH-1:0] w_in_0_81 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_82 = 'b000000001;
logic signed [WIDTH-1:0] w_in_0_83 = 'b111111010;
logic signed [WIDTH-1:0] w_in_0_84 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_85 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_86 = 'b000000011;
logic signed [WIDTH-1:0] w_in_0_87 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_88 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_89 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_90 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_91 = 'b000000011;
logic signed [WIDTH-1:0] w_in_0_92 = 'b000000001;
logic signed [WIDTH-1:0] w_in_0_93 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_94 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_95 = 'b111111001;
logic signed [WIDTH-1:0] w_in_0_96 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_97 = 'b111111000;
logic signed [WIDTH-1:0] w_in_0_98 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_99 = 'b000000100;
logic signed [WIDTH-1:0] w_in_0_100 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_101 = 'b111111010;
logic signed [WIDTH-1:0] w_in_0_102 = 'b111110111;
logic signed [WIDTH-1:0] w_in_0_103 = 'b000000101;
logic signed [WIDTH-1:0] w_in_0_104 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_105 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_106 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_107 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_108 = 'b000000001;
logic signed [WIDTH-1:0] w_in_0_109 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_110 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_111 = 'b000000100;
logic signed [WIDTH-1:0] w_in_0_112 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_113 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_114 = 'b000000001;
logic signed [WIDTH-1:0] w_in_0_115 = 'b000000001;
logic signed [WIDTH-1:0] w_in_0_116 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_117 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_118 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_119 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_120 = 'b000000001;
logic signed [WIDTH-1:0] w_in_0_121 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_122 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_123 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_124 = 'b000000111;
logic signed [WIDTH-1:0] w_in_0_125 = 'b000000101;
logic signed [WIDTH-1:0] w_in_0_126 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_127 = 'b000000101;
logic signed [WIDTH-1:0] w_in_0_128 = 'b000000110;
logic signed [WIDTH-1:0] w_in_0_129 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_130 = 'b000001001;
logic signed [WIDTH-1:0] w_in_0_131 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_132 = 'b000000101;
logic signed [WIDTH-1:0] w_in_0_133 = 'b000000001;
logic signed [WIDTH-1:0] w_in_0_134 = 'b111111001;
logic signed [WIDTH-1:0] w_in_0_135 = 'b000001001;
logic signed [WIDTH-1:0] w_in_0_136 = 'b000001011;
logic signed [WIDTH-1:0] w_in_0_137 = 'b000000110;
logic signed [WIDTH-1:0] w_in_0_138 = 'b000001000;
logic signed [WIDTH-1:0] w_in_0_139 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_140 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_141 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_142 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_143 = 'b111111001;
logic signed [WIDTH-1:0] w_in_0_144 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_145 = 'b000000101;
logic signed [WIDTH-1:0] w_in_0_146 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_147 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_148 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_149 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_150 = 'b000001001;
logic signed [WIDTH-1:0] w_in_0_151 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_152 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_153 = 'b000000011;
logic signed [WIDTH-1:0] w_in_0_154 = 'b111111010;
logic signed [WIDTH-1:0] w_in_0_155 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_156 = 'b000000110;
logic signed [WIDTH-1:0] w_in_0_157 = 'b000000101;
logic signed [WIDTH-1:0] w_in_0_158 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_159 = 'b000000101;
logic signed [WIDTH-1:0] w_in_0_160 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_161 = 'b000000011;
logic signed [WIDTH-1:0] w_in_0_162 = 'b000000111;
logic signed [WIDTH-1:0] w_in_0_163 = 'b000001000;
logic signed [WIDTH-1:0] w_in_0_164 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_165 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_166 = 'b111111000;
logic signed [WIDTH-1:0] w_in_0_167 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_168 = 'b000000100;
logic signed [WIDTH-1:0] w_in_0_169 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_170 = 'b000001001;
logic signed [WIDTH-1:0] w_in_0_171 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_172 = 'b000000100;
logic signed [WIDTH-1:0] w_in_0_173 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_174 = 'b111111001;
logic signed [WIDTH-1:0] w_in_0_175 = 'b000001000;
logic signed [WIDTH-1:0] w_in_0_176 = 'b111111010;
logic signed [WIDTH-1:0] w_in_0_177 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_178 = 'b000000100;
logic signed [WIDTH-1:0] w_in_0_179 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_180 = 'b000000100;
logic signed [WIDTH-1:0] w_in_0_181 = 'b111110010;
logic signed [WIDTH-1:0] w_in_0_182 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_183 = 'b000000001;
logic signed [WIDTH-1:0] w_in_0_184 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_185 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_186 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_187 = 'b111111010;
logic signed [WIDTH-1:0] w_in_0_188 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_189 = 'b111110100;
logic signed [WIDTH-1:0] w_in_0_190 = 'b111110001;
logic signed [WIDTH-1:0] w_in_0_191 = 'b111110000;
logic signed [WIDTH-1:0] w_in_0_192 = 'b111110101;
logic signed [WIDTH-1:0] w_in_0_193 = 'b111110101;
logic signed [WIDTH-1:0] w_in_0_194 = 'b000000011;
logic signed [WIDTH-1:0] w_in_0_195 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_196 = 'b000000110;
logic signed [WIDTH-1:0] w_in_0_197 = 'b000001000;
logic signed [WIDTH-1:0] w_in_0_198 = 'b111111001;
logic signed [WIDTH-1:0] w_in_0_199 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_200 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_201 = 'b111110100;
logic signed [WIDTH-1:0] w_in_0_202 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_203 = 'b000000101;
logic signed [WIDTH-1:0] w_in_0_204 = 'b000000110;
logic signed [WIDTH-1:0] w_in_0_205 = 'b111111010;
logic signed [WIDTH-1:0] w_in_0_206 = 'b000000110;
logic signed [WIDTH-1:0] w_in_0_207 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_208 = 'b000000001;
logic signed [WIDTH-1:0] w_in_0_209 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_210 = 'b000000001;
logic signed [WIDTH-1:0] w_in_0_211 = 'b000000111;
logic signed [WIDTH-1:0] w_in_0_212 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_213 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_214 = 'b000001000;
logic signed [WIDTH-1:0] w_in_0_215 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_216 = 'b000000111;
logic signed [WIDTH-1:0] w_in_0_217 = 'b000000011;
logic signed [WIDTH-1:0] w_in_0_218 = 'b000000100;
logic signed [WIDTH-1:0] w_in_0_219 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_220 = 'b000000110;
logic signed [WIDTH-1:0] w_in_0_221 = 'b000001001;
logic signed [WIDTH-1:0] w_in_0_222 = 'b000000110;
logic signed [WIDTH-1:0] w_in_0_223 = 'b000000011;
logic signed [WIDTH-1:0] w_in_0_224 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_225 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_226 = 'b111110100;
logic signed [WIDTH-1:0] w_in_0_227 = 'b111111010;
logic signed [WIDTH-1:0] w_in_0_228 = 'b000001000;
logic signed [WIDTH-1:0] w_in_0_229 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_230 = 'b000000110;
logic signed [WIDTH-1:0] w_in_0_231 = 'b111110111;
logic signed [WIDTH-1:0] w_in_0_232 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_233 = 'b111111000;
logic signed [WIDTH-1:0] w_in_0_234 = 'b111110111;
logic signed [WIDTH-1:0] w_in_0_235 = 'b111110111;
logic signed [WIDTH-1:0] w_in_0_236 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_237 = 'b000000001;
logic signed [WIDTH-1:0] w_in_0_238 = 'b000010010;
logic signed [WIDTH-1:0] w_in_0_239 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_240 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_241 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_242 = 'b111111000;
logic signed [WIDTH-1:0] w_in_0_243 = 'b000001100;
logic signed [WIDTH-1:0] w_in_0_244 = 'b111110111;
logic signed [WIDTH-1:0] w_in_0_245 = 'b000000011;
logic signed [WIDTH-1:0] w_in_0_246 = 'b000001001;
logic signed [WIDTH-1:0] w_in_0_247 = 'b000000001;
logic signed [WIDTH-1:0] w_in_0_248 = 'b000010010;
logic signed [WIDTH-1:0] w_in_0_249 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_250 = 'b000010011;
logic signed [WIDTH-1:0] w_in_0_251 = 'b000000011;
logic signed [WIDTH-1:0] w_in_0_252 = 'b111111000;
logic signed [WIDTH-1:0] w_in_0_253 = 'b000001001;
logic signed [WIDTH-1:0] w_in_0_254 = 'b000001100;
logic signed [WIDTH-1:0] w_in_0_255 = 'b111111000;
logic signed [WIDTH-1:0] w_in_1_0 = 'b111111100;
logic signed [WIDTH-1:0] w_in_1_1 = 'b000000010;
logic signed [WIDTH-1:0] w_in_1_2 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_3 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_4 = 'b111111111;
logic signed [WIDTH-1:0] w_in_1_5 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_6 = 'b111111001;
logic signed [WIDTH-1:0] w_in_1_7 = 'b111111100;
logic signed [WIDTH-1:0] w_in_1_8 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_9 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_10 = 'b000000010;
logic signed [WIDTH-1:0] w_in_1_11 = 'b000000111;
logic signed [WIDTH-1:0] w_in_1_12 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_13 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_14 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_15 = 'b000000010;
logic signed [WIDTH-1:0] w_in_1_16 = 'b111111111;
logic signed [WIDTH-1:0] w_in_1_17 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_18 = 'b000001000;
logic signed [WIDTH-1:0] w_in_1_19 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_20 = 'b111111111;
logic signed [WIDTH-1:0] w_in_1_21 = 'b000000001;
logic signed [WIDTH-1:0] w_in_1_22 = 'b000000110;
logic signed [WIDTH-1:0] w_in_1_23 = 'b000000001;
logic signed [WIDTH-1:0] w_in_1_24 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_25 = 'b111111111;
logic signed [WIDTH-1:0] w_in_1_26 = 'b111111001;
logic signed [WIDTH-1:0] w_in_1_27 = 'b000000010;
logic signed [WIDTH-1:0] w_in_1_28 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_29 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_30 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_31 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_32 = 'b111111111;
logic signed [WIDTH-1:0] w_in_1_33 = 'b111111011;
logic signed [WIDTH-1:0] w_in_1_34 = 'b111111010;
logic signed [WIDTH-1:0] w_in_1_35 = 'b111111101;
logic signed [WIDTH-1:0] w_in_1_36 = 'b111111101;
logic signed [WIDTH-1:0] w_in_1_37 = 'b111110110;
logic signed [WIDTH-1:0] w_in_1_38 = 'b000000010;
logic signed [WIDTH-1:0] w_in_1_39 = 'b111111111;
logic signed [WIDTH-1:0] w_in_1_40 = 'b111111111;
logic signed [WIDTH-1:0] w_in_1_41 = 'b000000111;
logic signed [WIDTH-1:0] w_in_1_42 = 'b111111011;
logic signed [WIDTH-1:0] w_in_1_43 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_44 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_45 = 'b111111100;
logic signed [WIDTH-1:0] w_in_1_46 = 'b111111011;
logic signed [WIDTH-1:0] w_in_1_47 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_48 = 'b000000010;
logic signed [WIDTH-1:0] w_in_1_49 = 'b000001001;
logic signed [WIDTH-1:0] w_in_1_50 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_51 = 'b000000010;
logic signed [WIDTH-1:0] w_in_1_52 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_53 = 'b111111010;
logic signed [WIDTH-1:0] w_in_1_54 = 'b111111001;
logic signed [WIDTH-1:0] w_in_1_55 = 'b111111101;
logic signed [WIDTH-1:0] w_in_1_56 = 'b000000111;
logic signed [WIDTH-1:0] w_in_1_57 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_58 = 'b000001000;
logic signed [WIDTH-1:0] w_in_1_59 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_60 = 'b111110111;
logic signed [WIDTH-1:0] w_in_1_61 = 'b111110010;
logic signed [WIDTH-1:0] w_in_1_62 = 'b111110000;
logic signed [WIDTH-1:0] w_in_1_63 = 'b000000011;
logic signed [WIDTH-1:0] w_in_1_64 = 'b000000110;
logic signed [WIDTH-1:0] w_in_1_65 = 'b000000010;
logic signed [WIDTH-1:0] w_in_1_66 = 'b000000001;
logic signed [WIDTH-1:0] w_in_1_67 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_68 = 'b000000001;
logic signed [WIDTH-1:0] w_in_1_69 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_70 = 'b111111010;
logic signed [WIDTH-1:0] w_in_1_71 = 'b111111011;
logic signed [WIDTH-1:0] w_in_1_72 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_73 = 'b000001000;
logic signed [WIDTH-1:0] w_in_1_74 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_75 = 'b111111000;
logic signed [WIDTH-1:0] w_in_1_76 = 'b111111011;
logic signed [WIDTH-1:0] w_in_1_77 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_78 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_79 = 'b000000110;
logic signed [WIDTH-1:0] w_in_1_80 = 'b111111000;
logic signed [WIDTH-1:0] w_in_1_81 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_82 = 'b000001001;
logic signed [WIDTH-1:0] w_in_1_83 = 'b111111011;
logic signed [WIDTH-1:0] w_in_1_84 = 'b111111011;
logic signed [WIDTH-1:0] w_in_1_85 = 'b111111001;
logic signed [WIDTH-1:0] w_in_1_86 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_87 = 'b000001010;
logic signed [WIDTH-1:0] w_in_1_88 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_89 = 'b111111100;
logic signed [WIDTH-1:0] w_in_1_90 = 'b111111101;
logic signed [WIDTH-1:0] w_in_1_91 = 'b111111100;
logic signed [WIDTH-1:0] w_in_1_92 = 'b111111101;
logic signed [WIDTH-1:0] w_in_1_93 = 'b111111010;
logic signed [WIDTH-1:0] w_in_1_94 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_95 = 'b111111010;
logic signed [WIDTH-1:0] w_in_1_96 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_97 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_98 = 'b111111100;
logic signed [WIDTH-1:0] w_in_1_99 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_100 = 'b111110111;
logic signed [WIDTH-1:0] w_in_1_101 = 'b000000001;
logic signed [WIDTH-1:0] w_in_1_102 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_103 = 'b111111100;
logic signed [WIDTH-1:0] w_in_1_104 = 'b000000110;
logic signed [WIDTH-1:0] w_in_1_105 = 'b000000011;
logic signed [WIDTH-1:0] w_in_1_106 = 'b000000111;
logic signed [WIDTH-1:0] w_in_1_107 = 'b000000110;
logic signed [WIDTH-1:0] w_in_1_108 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_109 = 'b000000111;
logic signed [WIDTH-1:0] w_in_1_110 = 'b000000010;
logic signed [WIDTH-1:0] w_in_1_111 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_112 = 'b111111010;
logic signed [WIDTH-1:0] w_in_1_113 = 'b111111111;
logic signed [WIDTH-1:0] w_in_1_114 = 'b111111101;
logic signed [WIDTH-1:0] w_in_1_115 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_116 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_117 = 'b000000011;
logic signed [WIDTH-1:0] w_in_1_118 = 'b111111000;
logic signed [WIDTH-1:0] w_in_1_119 = 'b000001010;
logic signed [WIDTH-1:0] w_in_1_120 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_121 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_122 = 'b111111111;
logic signed [WIDTH-1:0] w_in_1_123 = 'b000000111;
logic signed [WIDTH-1:0] w_in_1_124 = 'b111110111;
logic signed [WIDTH-1:0] w_in_1_125 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_126 = 'b111111101;
logic signed [WIDTH-1:0] w_in_1_127 = 'b111111101;
logic signed [WIDTH-1:0] w_in_1_128 = 'b000000011;
logic signed [WIDTH-1:0] w_in_1_129 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_130 = 'b111111111;
logic signed [WIDTH-1:0] w_in_1_131 = 'b000000010;
logic signed [WIDTH-1:0] w_in_1_132 = 'b000000110;
logic signed [WIDTH-1:0] w_in_1_133 = 'b000000011;
logic signed [WIDTH-1:0] w_in_1_134 = 'b111110111;
logic signed [WIDTH-1:0] w_in_1_135 = 'b000000011;
logic signed [WIDTH-1:0] w_in_1_136 = 'b111110100;
logic signed [WIDTH-1:0] w_in_1_137 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_138 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_139 = 'b111111100;
logic signed [WIDTH-1:0] w_in_1_140 = 'b111111001;
logic signed [WIDTH-1:0] w_in_1_141 = 'b000000011;
logic signed [WIDTH-1:0] w_in_1_142 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_143 = 'b111110101;
logic signed [WIDTH-1:0] w_in_1_144 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_145 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_146 = 'b111110100;
logic signed [WIDTH-1:0] w_in_1_147 = 'b111111000;
logic signed [WIDTH-1:0] w_in_1_148 = 'b000000111;
logic signed [WIDTH-1:0] w_in_1_149 = 'b111111010;
logic signed [WIDTH-1:0] w_in_1_150 = 'b000000011;
logic signed [WIDTH-1:0] w_in_1_151 = 'b111111010;
logic signed [WIDTH-1:0] w_in_1_152 = 'b000000011;
logic signed [WIDTH-1:0] w_in_1_153 = 'b111111011;
logic signed [WIDTH-1:0] w_in_1_154 = 'b000001001;
logic signed [WIDTH-1:0] w_in_1_155 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_156 = 'b000000110;
logic signed [WIDTH-1:0] w_in_1_157 = 'b000001001;
logic signed [WIDTH-1:0] w_in_1_158 = 'b111111111;
logic signed [WIDTH-1:0] w_in_1_159 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_160 = 'b000001011;
logic signed [WIDTH-1:0] w_in_1_161 = 'b111111000;
logic signed [WIDTH-1:0] w_in_1_162 = 'b111111000;
logic signed [WIDTH-1:0] w_in_1_163 = 'b111111100;
logic signed [WIDTH-1:0] w_in_1_164 = 'b000001010;
logic signed [WIDTH-1:0] w_in_1_165 = 'b000001000;
logic signed [WIDTH-1:0] w_in_1_166 = 'b111111011;
logic signed [WIDTH-1:0] w_in_1_167 = 'b111110101;
logic signed [WIDTH-1:0] w_in_1_168 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_169 = 'b111111111;
logic signed [WIDTH-1:0] w_in_1_170 = 'b111111000;
logic signed [WIDTH-1:0] w_in_1_171 = 'b000000001;
logic signed [WIDTH-1:0] w_in_1_172 = 'b111111101;
logic signed [WIDTH-1:0] w_in_1_173 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_174 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_175 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_176 = 'b111111101;
logic signed [WIDTH-1:0] w_in_1_177 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_178 = 'b111111000;
logic signed [WIDTH-1:0] w_in_1_179 = 'b111111101;
logic signed [WIDTH-1:0] w_in_1_180 = 'b111111000;
logic signed [WIDTH-1:0] w_in_1_181 = 'b000000111;
logic signed [WIDTH-1:0] w_in_1_182 = 'b111111111;
logic signed [WIDTH-1:0] w_in_1_183 = 'b111111100;
logic signed [WIDTH-1:0] w_in_1_184 = 'b111111101;
logic signed [WIDTH-1:0] w_in_1_185 = 'b000000111;
logic signed [WIDTH-1:0] w_in_1_186 = 'b000001000;
logic signed [WIDTH-1:0] w_in_1_187 = 'b000001010;
logic signed [WIDTH-1:0] w_in_1_188 = 'b000001111;
logic signed [WIDTH-1:0] w_in_1_189 = 'b000001010;
logic signed [WIDTH-1:0] w_in_1_190 = 'b000010001;
logic signed [WIDTH-1:0] w_in_1_191 = 'b000001101;
logic signed [WIDTH-1:0] w_in_1_192 = 'b111110101;
logic signed [WIDTH-1:0] w_in_1_193 = 'b000001000;
logic signed [WIDTH-1:0] w_in_1_194 = 'b000000001;
logic signed [WIDTH-1:0] w_in_1_195 = 'b000001001;
logic signed [WIDTH-1:0] w_in_1_196 = 'b111110110;
logic signed [WIDTH-1:0] w_in_1_197 = 'b000000010;
logic signed [WIDTH-1:0] w_in_1_198 = 'b111110111;
logic signed [WIDTH-1:0] w_in_1_199 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_200 = 'b111110010;
logic signed [WIDTH-1:0] w_in_1_201 = 'b111110101;
logic signed [WIDTH-1:0] w_in_1_202 = 'b000001001;
logic signed [WIDTH-1:0] w_in_1_203 = 'b111110101;
logic signed [WIDTH-1:0] w_in_1_204 = 'b111110101;
logic signed [WIDTH-1:0] w_in_1_205 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_206 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_207 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_208 = 'b000001011;
logic signed [WIDTH-1:0] w_in_1_209 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_210 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_211 = 'b000001101;
logic signed [WIDTH-1:0] w_in_1_212 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_213 = 'b111111000;
logic signed [WIDTH-1:0] w_in_1_214 = 'b111111101;
logic signed [WIDTH-1:0] w_in_1_215 = 'b111111100;
logic signed [WIDTH-1:0] w_in_1_216 = 'b111110110;
logic signed [WIDTH-1:0] w_in_1_217 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_218 = 'b111111000;
logic signed [WIDTH-1:0] w_in_1_219 = 'b111110110;
logic signed [WIDTH-1:0] w_in_1_220 = 'b000001101;
logic signed [WIDTH-1:0] w_in_1_221 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_222 = 'b000000001;
logic signed [WIDTH-1:0] w_in_1_223 = 'b000000111;
logic signed [WIDTH-1:0] w_in_1_224 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_225 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_226 = 'b000000111;
logic signed [WIDTH-1:0] w_in_1_227 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_228 = 'b111110111;
logic signed [WIDTH-1:0] w_in_1_229 = 'b111110110;
logic signed [WIDTH-1:0] w_in_1_230 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_231 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_232 = 'b111110100;
logic signed [WIDTH-1:0] w_in_1_233 = 'b111110110;
logic signed [WIDTH-1:0] w_in_1_234 = 'b000001000;
logic signed [WIDTH-1:0] w_in_1_235 = 'b000000001;
logic signed [WIDTH-1:0] w_in_1_236 = 'b000000011;
logic signed [WIDTH-1:0] w_in_1_237 = 'b000001100;
logic signed [WIDTH-1:0] w_in_1_238 = 'b111111111;
logic signed [WIDTH-1:0] w_in_1_239 = 'b000001010;
logic signed [WIDTH-1:0] w_in_1_240 = 'b000000001;
logic signed [WIDTH-1:0] w_in_1_241 = 'b111111111;
logic signed [WIDTH-1:0] w_in_1_242 = 'b111111011;
logic signed [WIDTH-1:0] w_in_1_243 = 'b000000110;
logic signed [WIDTH-1:0] w_in_1_244 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_245 = 'b111110110;
logic signed [WIDTH-1:0] w_in_1_246 = 'b000001100;
logic signed [WIDTH-1:0] w_in_1_247 = 'b000000010;
logic signed [WIDTH-1:0] w_in_1_248 = 'b111111010;
logic signed [WIDTH-1:0] w_in_1_249 = 'b000000110;
logic signed [WIDTH-1:0] w_in_1_250 = 'b111111011;
logic signed [WIDTH-1:0] w_in_1_251 = 'b000001011;
logic signed [WIDTH-1:0] w_in_1_252 = 'b000001011;
logic signed [WIDTH-1:0] w_in_1_253 = 'b000000011;
logic signed [WIDTH-1:0] w_in_1_254 = 'b000000001;
logic signed [WIDTH-1:0] w_in_1_255 = 'b000001001;
logic signed [WIDTH-1:0] w_in_2_0 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_1 = 'b000000101;
logic signed [WIDTH-1:0] w_in_2_2 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_3 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_4 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_5 = 'b111111011;
logic signed [WIDTH-1:0] w_in_2_6 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_7 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_8 = 'b111111001;
logic signed [WIDTH-1:0] w_in_2_9 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_10 = 'b000001000;
logic signed [WIDTH-1:0] w_in_2_11 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_12 = 'b000000101;
logic signed [WIDTH-1:0] w_in_2_13 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_14 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_15 = 'b000000110;
logic signed [WIDTH-1:0] w_in_2_16 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_17 = 'b000000111;
logic signed [WIDTH-1:0] w_in_2_18 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_19 = 'b000000101;
logic signed [WIDTH-1:0] w_in_2_20 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_21 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_22 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_23 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_24 = 'b111111011;
logic signed [WIDTH-1:0] w_in_2_25 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_26 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_27 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_28 = 'b000000111;
logic signed [WIDTH-1:0] w_in_2_29 = 'b111111001;
logic signed [WIDTH-1:0] w_in_2_30 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_31 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_32 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_33 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_34 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_35 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_36 = 'b000001000;
logic signed [WIDTH-1:0] w_in_2_37 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_38 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_39 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_40 = 'b000000101;
logic signed [WIDTH-1:0] w_in_2_41 = 'b111111010;
logic signed [WIDTH-1:0] w_in_2_42 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_43 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_44 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_45 = 'b111111100;
logic signed [WIDTH-1:0] w_in_2_46 = 'b111111010;
logic signed [WIDTH-1:0] w_in_2_47 = 'b000000111;
logic signed [WIDTH-1:0] w_in_2_48 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_49 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_50 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_51 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_52 = 'b111111001;
logic signed [WIDTH-1:0] w_in_2_53 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_54 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_55 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_56 = 'b000000101;
logic signed [WIDTH-1:0] w_in_2_57 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_58 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_59 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_60 = 'b111111011;
logic signed [WIDTH-1:0] w_in_2_61 = 'b111111010;
logic signed [WIDTH-1:0] w_in_2_62 = 'b111111010;
logic signed [WIDTH-1:0] w_in_2_63 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_64 = 'b111111100;
logic signed [WIDTH-1:0] w_in_2_65 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_66 = 'b000000110;
logic signed [WIDTH-1:0] w_in_2_67 = 'b000000101;
logic signed [WIDTH-1:0] w_in_2_68 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_69 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_70 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_71 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_72 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_73 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_74 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_75 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_76 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_77 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_78 = 'b111111011;
logic signed [WIDTH-1:0] w_in_2_79 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_80 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_81 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_82 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_83 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_84 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_85 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_86 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_87 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_88 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_89 = 'b000000110;
logic signed [WIDTH-1:0] w_in_2_90 = 'b111111010;
logic signed [WIDTH-1:0] w_in_2_91 = 'b111111010;
logic signed [WIDTH-1:0] w_in_2_92 = 'b000000111;
logic signed [WIDTH-1:0] w_in_2_93 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_94 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_95 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_96 = 'b111111100;
logic signed [WIDTH-1:0] w_in_2_97 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_98 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_99 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_100 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_101 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_102 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_103 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_104 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_105 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_106 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_107 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_108 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_109 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_110 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_111 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_112 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_113 = 'b111111001;
logic signed [WIDTH-1:0] w_in_2_114 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_115 = 'b000000101;
logic signed [WIDTH-1:0] w_in_2_116 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_117 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_118 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_119 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_120 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_121 = 'b000000110;
logic signed [WIDTH-1:0] w_in_2_122 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_123 = 'b111111100;
logic signed [WIDTH-1:0] w_in_2_124 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_125 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_126 = 'b000000101;
logic signed [WIDTH-1:0] w_in_2_127 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_128 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_129 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_130 = 'b111111001;
logic signed [WIDTH-1:0] w_in_2_131 = 'b111111100;
logic signed [WIDTH-1:0] w_in_2_132 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_133 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_134 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_135 = 'b111111011;
logic signed [WIDTH-1:0] w_in_2_136 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_137 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_138 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_139 = 'b111111001;
logic signed [WIDTH-1:0] w_in_2_140 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_141 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_142 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_143 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_144 = 'b111111011;
logic signed [WIDTH-1:0] w_in_2_145 = 'b000000111;
logic signed [WIDTH-1:0] w_in_2_146 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_147 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_148 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_149 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_150 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_151 = 'b000000111;
logic signed [WIDTH-1:0] w_in_2_152 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_153 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_154 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_155 = 'b111111001;
logic signed [WIDTH-1:0] w_in_2_156 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_157 = 'b000001000;
logic signed [WIDTH-1:0] w_in_2_158 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_159 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_160 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_161 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_162 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_163 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_164 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_165 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_166 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_167 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_168 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_169 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_170 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_171 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_172 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_173 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_174 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_175 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_176 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_177 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_178 = 'b111111100;
logic signed [WIDTH-1:0] w_in_2_179 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_180 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_181 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_182 = 'b111111001;
logic signed [WIDTH-1:0] w_in_2_183 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_184 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_185 = 'b111111011;
logic signed [WIDTH-1:0] w_in_2_186 = 'b111111100;
logic signed [WIDTH-1:0] w_in_2_187 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_188 = 'b000000101;
logic signed [WIDTH-1:0] w_in_2_189 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_190 = 'b000000101;
logic signed [WIDTH-1:0] w_in_2_191 = 'b000001001;
logic signed [WIDTH-1:0] w_in_2_192 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_193 = 'b000001000;
logic signed [WIDTH-1:0] w_in_2_194 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_195 = 'b000000110;
logic signed [WIDTH-1:0] w_in_2_196 = 'b111111010;
logic signed [WIDTH-1:0] w_in_2_197 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_198 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_199 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_200 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_201 = 'b000000101;
logic signed [WIDTH-1:0] w_in_2_202 = 'b111111100;
logic signed [WIDTH-1:0] w_in_2_203 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_204 = 'b111111100;
logic signed [WIDTH-1:0] w_in_2_205 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_206 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_207 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_208 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_209 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_210 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_211 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_212 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_213 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_214 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_215 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_216 = 'b000000111;
logic signed [WIDTH-1:0] w_in_2_217 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_218 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_219 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_220 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_221 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_222 = 'b111111100;
logic signed [WIDTH-1:0] w_in_2_223 = 'b000001000;
logic signed [WIDTH-1:0] w_in_2_224 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_225 = 'b111111011;
logic signed [WIDTH-1:0] w_in_2_226 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_227 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_228 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_229 = 'b111111001;
logic signed [WIDTH-1:0] w_in_2_230 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_231 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_232 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_233 = 'b000000101;
logic signed [WIDTH-1:0] w_in_2_234 = 'b111111011;
logic signed [WIDTH-1:0] w_in_2_235 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_236 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_237 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_238 = 'b000000110;
logic signed [WIDTH-1:0] w_in_2_239 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_240 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_241 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_242 = 'b111111100;
logic signed [WIDTH-1:0] w_in_2_243 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_244 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_245 = 'b111111100;
logic signed [WIDTH-1:0] w_in_2_246 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_247 = 'b111111001;
logic signed [WIDTH-1:0] w_in_2_248 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_249 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_250 = 'b111111100;
logic signed [WIDTH-1:0] w_in_2_251 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_252 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_253 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_254 = 'b111111010;
logic signed [WIDTH-1:0] w_in_2_255 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_0 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_1 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_2 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_3 = 'b111111101;
logic signed [WIDTH-1:0] w_in_3_4 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_5 = 'b000000011;
logic signed [WIDTH-1:0] w_in_3_6 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_7 = 'b111111011;
logic signed [WIDTH-1:0] w_in_3_8 = 'b111111001;
logic signed [WIDTH-1:0] w_in_3_9 = 'b111111101;
logic signed [WIDTH-1:0] w_in_3_10 = 'b111111001;
logic signed [WIDTH-1:0] w_in_3_11 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_12 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_13 = 'b000000011;
logic signed [WIDTH-1:0] w_in_3_14 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_15 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_16 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_17 = 'b111111101;
logic signed [WIDTH-1:0] w_in_3_18 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_19 = 'b111111011;
logic signed [WIDTH-1:0] w_in_3_20 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_21 = 'b000000011;
logic signed [WIDTH-1:0] w_in_3_22 = 'b000001000;
logic signed [WIDTH-1:0] w_in_3_23 = 'b000000101;
logic signed [WIDTH-1:0] w_in_3_24 = 'b111111001;
logic signed [WIDTH-1:0] w_in_3_25 = 'b111111010;
logic signed [WIDTH-1:0] w_in_3_26 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_27 = 'b111111001;
logic signed [WIDTH-1:0] w_in_3_28 = 'b000000110;
logic signed [WIDTH-1:0] w_in_3_29 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_30 = 'b000000110;
logic signed [WIDTH-1:0] w_in_3_31 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_32 = 'b111111001;
logic signed [WIDTH-1:0] w_in_3_33 = 'b111111010;
logic signed [WIDTH-1:0] w_in_3_34 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_35 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_36 = 'b111111010;
logic signed [WIDTH-1:0] w_in_3_37 = 'b111111011;
logic signed [WIDTH-1:0] w_in_3_38 = 'b111111101;
logic signed [WIDTH-1:0] w_in_3_39 = 'b000000010;
logic signed [WIDTH-1:0] w_in_3_40 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_41 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_42 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_43 = 'b111111101;
logic signed [WIDTH-1:0] w_in_3_44 = 'b111111000;
logic signed [WIDTH-1:0] w_in_3_45 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_46 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_47 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_48 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_49 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_50 = 'b000000101;
logic signed [WIDTH-1:0] w_in_3_51 = 'b111111101;
logic signed [WIDTH-1:0] w_in_3_52 = 'b000000111;
logic signed [WIDTH-1:0] w_in_3_53 = 'b000000100;
logic signed [WIDTH-1:0] w_in_3_54 = 'b000001000;
logic signed [WIDTH-1:0] w_in_3_55 = 'b000000110;
logic signed [WIDTH-1:0] w_in_3_56 = 'b000000011;
logic signed [WIDTH-1:0] w_in_3_57 = 'b111111001;
logic signed [WIDTH-1:0] w_in_3_58 = 'b000000100;
logic signed [WIDTH-1:0] w_in_3_59 = 'b000001110;
logic signed [WIDTH-1:0] w_in_3_60 = 'b000001010;
logic signed [WIDTH-1:0] w_in_3_61 = 'b000001011;
logic signed [WIDTH-1:0] w_in_3_62 = 'b000001101;
logic signed [WIDTH-1:0] w_in_3_63 = 'b000001100;
logic signed [WIDTH-1:0] w_in_3_64 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_65 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_66 = 'b000000010;
logic signed [WIDTH-1:0] w_in_3_67 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_68 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_69 = 'b111111011;
logic signed [WIDTH-1:0] w_in_3_70 = 'b000000110;
logic signed [WIDTH-1:0] w_in_3_71 = 'b111111001;
logic signed [WIDTH-1:0] w_in_3_72 = 'b111111010;
logic signed [WIDTH-1:0] w_in_3_73 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_74 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_75 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_76 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_77 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_78 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_79 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_80 = 'b000000101;
logic signed [WIDTH-1:0] w_in_3_81 = 'b111111011;
logic signed [WIDTH-1:0] w_in_3_82 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_83 = 'b111111010;
logic signed [WIDTH-1:0] w_in_3_84 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_85 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_86 = 'b000000011;
logic signed [WIDTH-1:0] w_in_3_87 = 'b000000010;
logic signed [WIDTH-1:0] w_in_3_88 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_89 = 'b111111101;
logic signed [WIDTH-1:0] w_in_3_90 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_91 = 'b000000011;
logic signed [WIDTH-1:0] w_in_3_92 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_93 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_94 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_95 = 'b111111001;
logic signed [WIDTH-1:0] w_in_3_96 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_97 = 'b111111000;
logic signed [WIDTH-1:0] w_in_3_98 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_99 = 'b000000100;
logic signed [WIDTH-1:0] w_in_3_100 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_101 = 'b111111010;
logic signed [WIDTH-1:0] w_in_3_102 = 'b111110111;
logic signed [WIDTH-1:0] w_in_3_103 = 'b000000101;
logic signed [WIDTH-1:0] w_in_3_104 = 'b111111101;
logic signed [WIDTH-1:0] w_in_3_105 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_106 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_107 = 'b111111101;
logic signed [WIDTH-1:0] w_in_3_108 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_109 = 'b111111101;
logic signed [WIDTH-1:0] w_in_3_110 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_111 = 'b000000100;
logic signed [WIDTH-1:0] w_in_3_112 = 'b000000010;
logic signed [WIDTH-1:0] w_in_3_113 = 'b000000010;
logic signed [WIDTH-1:0] w_in_3_114 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_115 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_116 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_117 = 'b111111101;
logic signed [WIDTH-1:0] w_in_3_118 = 'b000000010;
logic signed [WIDTH-1:0] w_in_3_119 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_120 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_121 = 'b111111011;
logic signed [WIDTH-1:0] w_in_3_122 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_123 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_124 = 'b000000111;
logic signed [WIDTH-1:0] w_in_3_125 = 'b000000101;
logic signed [WIDTH-1:0] w_in_3_126 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_127 = 'b000000101;
logic signed [WIDTH-1:0] w_in_3_128 = 'b000000110;
logic signed [WIDTH-1:0] w_in_3_129 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_130 = 'b000001001;
logic signed [WIDTH-1:0] w_in_3_131 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_132 = 'b000000101;
logic signed [WIDTH-1:0] w_in_3_133 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_134 = 'b111111001;
logic signed [WIDTH-1:0] w_in_3_135 = 'b000001001;
logic signed [WIDTH-1:0] w_in_3_136 = 'b000001011;
logic signed [WIDTH-1:0] w_in_3_137 = 'b000000110;
logic signed [WIDTH-1:0] w_in_3_138 = 'b000001000;
logic signed [WIDTH-1:0] w_in_3_139 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_140 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_141 = 'b000000010;
logic signed [WIDTH-1:0] w_in_3_142 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_143 = 'b111111001;
logic signed [WIDTH-1:0] w_in_3_144 = 'b111111101;
logic signed [WIDTH-1:0] w_in_3_145 = 'b000000101;
logic signed [WIDTH-1:0] w_in_3_146 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_147 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_148 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_149 = 'b111111011;
logic signed [WIDTH-1:0] w_in_3_150 = 'b000001001;
logic signed [WIDTH-1:0] w_in_3_151 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_152 = 'b111111011;
logic signed [WIDTH-1:0] w_in_3_153 = 'b000000011;
logic signed [WIDTH-1:0] w_in_3_154 = 'b111111010;
logic signed [WIDTH-1:0] w_in_3_155 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_156 = 'b000000110;
logic signed [WIDTH-1:0] w_in_3_157 = 'b000000101;
logic signed [WIDTH-1:0] w_in_3_158 = 'b111111011;
logic signed [WIDTH-1:0] w_in_3_159 = 'b000000101;
logic signed [WIDTH-1:0] w_in_3_160 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_161 = 'b000000011;
logic signed [WIDTH-1:0] w_in_3_162 = 'b000000111;
logic signed [WIDTH-1:0] w_in_3_163 = 'b000001000;
logic signed [WIDTH-1:0] w_in_3_164 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_165 = 'b000000010;
logic signed [WIDTH-1:0] w_in_3_166 = 'b111111000;
logic signed [WIDTH-1:0] w_in_3_167 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_168 = 'b000000100;
logic signed [WIDTH-1:0] w_in_3_169 = 'b111111101;
logic signed [WIDTH-1:0] w_in_3_170 = 'b000001001;
logic signed [WIDTH-1:0] w_in_3_171 = 'b000000010;
logic signed [WIDTH-1:0] w_in_3_172 = 'b000000100;
logic signed [WIDTH-1:0] w_in_3_173 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_174 = 'b111111001;
logic signed [WIDTH-1:0] w_in_3_175 = 'b000001000;
logic signed [WIDTH-1:0] w_in_3_176 = 'b111111010;
logic signed [WIDTH-1:0] w_in_3_177 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_178 = 'b000000100;
logic signed [WIDTH-1:0] w_in_3_179 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_180 = 'b000000100;
logic signed [WIDTH-1:0] w_in_3_181 = 'b111110010;
logic signed [WIDTH-1:0] w_in_3_182 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_183 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_184 = 'b111111011;
logic signed [WIDTH-1:0] w_in_3_185 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_186 = 'b111111011;
logic signed [WIDTH-1:0] w_in_3_187 = 'b111111010;
logic signed [WIDTH-1:0] w_in_3_188 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_189 = 'b111110100;
logic signed [WIDTH-1:0] w_in_3_190 = 'b111110001;
logic signed [WIDTH-1:0] w_in_3_191 = 'b111110000;
logic signed [WIDTH-1:0] w_in_3_192 = 'b111110101;
logic signed [WIDTH-1:0] w_in_3_193 = 'b111110101;
logic signed [WIDTH-1:0] w_in_3_194 = 'b000000011;
logic signed [WIDTH-1:0] w_in_3_195 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_196 = 'b000000110;
logic signed [WIDTH-1:0] w_in_3_197 = 'b000001000;
logic signed [WIDTH-1:0] w_in_3_198 = 'b111111001;
logic signed [WIDTH-1:0] w_in_3_199 = 'b000000010;
logic signed [WIDTH-1:0] w_in_3_200 = 'b111111011;
logic signed [WIDTH-1:0] w_in_3_201 = 'b111110100;
logic signed [WIDTH-1:0] w_in_3_202 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_203 = 'b000000101;
logic signed [WIDTH-1:0] w_in_3_204 = 'b000000110;
logic signed [WIDTH-1:0] w_in_3_205 = 'b111111010;
logic signed [WIDTH-1:0] w_in_3_206 = 'b000000110;
logic signed [WIDTH-1:0] w_in_3_207 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_208 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_209 = 'b111111101;
logic signed [WIDTH-1:0] w_in_3_210 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_211 = 'b000000111;
logic signed [WIDTH-1:0] w_in_3_212 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_213 = 'b111111101;
logic signed [WIDTH-1:0] w_in_3_214 = 'b000001000;
logic signed [WIDTH-1:0] w_in_3_215 = 'b111111101;
logic signed [WIDTH-1:0] w_in_3_216 = 'b000000111;
logic signed [WIDTH-1:0] w_in_3_217 = 'b000000011;
logic signed [WIDTH-1:0] w_in_3_218 = 'b000000100;
logic signed [WIDTH-1:0] w_in_3_219 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_220 = 'b000000110;
logic signed [WIDTH-1:0] w_in_3_221 = 'b000001001;
logic signed [WIDTH-1:0] w_in_3_222 = 'b000000110;
logic signed [WIDTH-1:0] w_in_3_223 = 'b000000011;
logic signed [WIDTH-1:0] w_in_3_224 = 'b111111011;
logic signed [WIDTH-1:0] w_in_3_225 = 'b111111101;
logic signed [WIDTH-1:0] w_in_3_226 = 'b111110100;
logic signed [WIDTH-1:0] w_in_3_227 = 'b111111010;
logic signed [WIDTH-1:0] w_in_3_228 = 'b000001000;
logic signed [WIDTH-1:0] w_in_3_229 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_230 = 'b000000110;
logic signed [WIDTH-1:0] w_in_3_231 = 'b111110111;
logic signed [WIDTH-1:0] w_in_3_232 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_233 = 'b111111000;
logic signed [WIDTH-1:0] w_in_3_234 = 'b111110111;
logic signed [WIDTH-1:0] w_in_3_235 = 'b111110111;
logic signed [WIDTH-1:0] w_in_3_236 = 'b111111011;
logic signed [WIDTH-1:0] w_in_3_237 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_238 = 'b000010010;
logic signed [WIDTH-1:0] w_in_3_239 = 'b111111011;
logic signed [WIDTH-1:0] w_in_3_240 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_241 = 'b111111011;
logic signed [WIDTH-1:0] w_in_3_242 = 'b111111000;
logic signed [WIDTH-1:0] w_in_3_243 = 'b000001100;
logic signed [WIDTH-1:0] w_in_3_244 = 'b111110111;
logic signed [WIDTH-1:0] w_in_3_245 = 'b000000011;
logic signed [WIDTH-1:0] w_in_3_246 = 'b000001001;
logic signed [WIDTH-1:0] w_in_3_247 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_248 = 'b000010010;
logic signed [WIDTH-1:0] w_in_3_249 = 'b000000010;
logic signed [WIDTH-1:0] w_in_3_250 = 'b000010011;
logic signed [WIDTH-1:0] w_in_3_251 = 'b000000011;
logic signed [WIDTH-1:0] w_in_3_252 = 'b111111000;
logic signed [WIDTH-1:0] w_in_3_253 = 'b000001001;
logic signed [WIDTH-1:0] w_in_3_254 = 'b000001100;
logic signed [WIDTH-1:0] w_in_3_255 = 'b111111000;
logic signed [WIDTH-1:0] w_in_4_0 = 'b111111100;
logic signed [WIDTH-1:0] w_in_4_1 = 'b000000010;
logic signed [WIDTH-1:0] w_in_4_2 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_3 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_4 = 'b111111111;
logic signed [WIDTH-1:0] w_in_4_5 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_6 = 'b111111001;
logic signed [WIDTH-1:0] w_in_4_7 = 'b111111100;
logic signed [WIDTH-1:0] w_in_4_8 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_9 = 'b000000101;
logic signed [WIDTH-1:0] w_in_4_10 = 'b000000010;
logic signed [WIDTH-1:0] w_in_4_11 = 'b000000111;
logic signed [WIDTH-1:0] w_in_4_12 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_13 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_14 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_15 = 'b000000010;
logic signed [WIDTH-1:0] w_in_4_16 = 'b111111111;
logic signed [WIDTH-1:0] w_in_4_17 = 'b000000101;
logic signed [WIDTH-1:0] w_in_4_18 = 'b000001000;
logic signed [WIDTH-1:0] w_in_4_19 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_20 = 'b111111111;
logic signed [WIDTH-1:0] w_in_4_21 = 'b000000001;
logic signed [WIDTH-1:0] w_in_4_22 = 'b000000110;
logic signed [WIDTH-1:0] w_in_4_23 = 'b000000001;
logic signed [WIDTH-1:0] w_in_4_24 = 'b000000000;
logic signed [WIDTH-1:0] w_in_4_25 = 'b111111111;
logic signed [WIDTH-1:0] w_in_4_26 = 'b111111001;
logic signed [WIDTH-1:0] w_in_4_27 = 'b000000010;
logic signed [WIDTH-1:0] w_in_4_28 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_29 = 'b000000000;
logic signed [WIDTH-1:0] w_in_4_30 = 'b000000101;
logic signed [WIDTH-1:0] w_in_4_31 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_32 = 'b111111111;
logic signed [WIDTH-1:0] w_in_4_33 = 'b111111011;
logic signed [WIDTH-1:0] w_in_4_34 = 'b111111010;
logic signed [WIDTH-1:0] w_in_4_35 = 'b111111101;
logic signed [WIDTH-1:0] w_in_4_36 = 'b111111101;
logic signed [WIDTH-1:0] w_in_4_37 = 'b111110110;
logic signed [WIDTH-1:0] w_in_4_38 = 'b000000010;
logic signed [WIDTH-1:0] w_in_4_39 = 'b111111111;
logic signed [WIDTH-1:0] w_in_4_40 = 'b111111111;
logic signed [WIDTH-1:0] w_in_4_41 = 'b000000111;
logic signed [WIDTH-1:0] w_in_4_42 = 'b111111011;
logic signed [WIDTH-1:0] w_in_4_43 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_44 = 'b000000000;
logic signed [WIDTH-1:0] w_in_4_45 = 'b111111100;
logic signed [WIDTH-1:0] w_in_4_46 = 'b111111011;
logic signed [WIDTH-1:0] w_in_4_47 = 'b000000101;
logic signed [WIDTH-1:0] w_in_4_48 = 'b000000010;
logic signed [WIDTH-1:0] w_in_4_49 = 'b000001001;
logic signed [WIDTH-1:0] w_in_4_50 = 'b000000000;
logic signed [WIDTH-1:0] w_in_4_51 = 'b000000010;
logic signed [WIDTH-1:0] w_in_4_52 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_53 = 'b111111010;
logic signed [WIDTH-1:0] w_in_4_54 = 'b111111001;
logic signed [WIDTH-1:0] w_in_4_55 = 'b111111101;
logic signed [WIDTH-1:0] w_in_4_56 = 'b000000111;
logic signed [WIDTH-1:0] w_in_4_57 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_58 = 'b000001000;
logic signed [WIDTH-1:0] w_in_4_59 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_60 = 'b111110111;
logic signed [WIDTH-1:0] w_in_4_61 = 'b111110010;
logic signed [WIDTH-1:0] w_in_4_62 = 'b111110000;
logic signed [WIDTH-1:0] w_in_4_63 = 'b000000011;
logic signed [WIDTH-1:0] w_in_4_64 = 'b000000110;
logic signed [WIDTH-1:0] w_in_4_65 = 'b000000010;
logic signed [WIDTH-1:0] w_in_4_66 = 'b000000001;
logic signed [WIDTH-1:0] w_in_4_67 = 'b000000000;
logic signed [WIDTH-1:0] w_in_4_68 = 'b000000001;
logic signed [WIDTH-1:0] w_in_4_69 = 'b000000101;
logic signed [WIDTH-1:0] w_in_4_70 = 'b111111010;
logic signed [WIDTH-1:0] w_in_4_71 = 'b111111011;
logic signed [WIDTH-1:0] w_in_4_72 = 'b000000000;
logic signed [WIDTH-1:0] w_in_4_73 = 'b000001000;
logic signed [WIDTH-1:0] w_in_4_74 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_75 = 'b111111000;
logic signed [WIDTH-1:0] w_in_4_76 = 'b111111011;
logic signed [WIDTH-1:0] w_in_4_77 = 'b000000101;
logic signed [WIDTH-1:0] w_in_4_78 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_79 = 'b000000110;
logic signed [WIDTH-1:0] w_in_4_80 = 'b111111000;
logic signed [WIDTH-1:0] w_in_4_81 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_82 = 'b000001001;
logic signed [WIDTH-1:0] w_in_4_83 = 'b111111011;
logic signed [WIDTH-1:0] w_in_4_84 = 'b111111011;
logic signed [WIDTH-1:0] w_in_4_85 = 'b111111001;
logic signed [WIDTH-1:0] w_in_4_86 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_87 = 'b000001010;
logic signed [WIDTH-1:0] w_in_4_88 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_89 = 'b111111100;
logic signed [WIDTH-1:0] w_in_4_90 = 'b111111101;
logic signed [WIDTH-1:0] w_in_4_91 = 'b111111100;
logic signed [WIDTH-1:0] w_in_4_92 = 'b111111101;
logic signed [WIDTH-1:0] w_in_4_93 = 'b111111010;
logic signed [WIDTH-1:0] w_in_4_94 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_95 = 'b111111010;
logic signed [WIDTH-1:0] w_in_4_96 = 'b000000101;
logic signed [WIDTH-1:0] w_in_4_97 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_98 = 'b111111100;
logic signed [WIDTH-1:0] w_in_4_99 = 'b000000101;
logic signed [WIDTH-1:0] w_in_4_100 = 'b111110111;
logic signed [WIDTH-1:0] w_in_4_101 = 'b000000001;
logic signed [WIDTH-1:0] w_in_4_102 = 'b000000000;
logic signed [WIDTH-1:0] w_in_4_103 = 'b111111100;
logic signed [WIDTH-1:0] w_in_4_104 = 'b000000110;
logic signed [WIDTH-1:0] w_in_4_105 = 'b000000011;
logic signed [WIDTH-1:0] w_in_4_106 = 'b000000111;
logic signed [WIDTH-1:0] w_in_4_107 = 'b000000110;
logic signed [WIDTH-1:0] w_in_4_108 = 'b000000000;
logic signed [WIDTH-1:0] w_in_4_109 = 'b000000111;
logic signed [WIDTH-1:0] w_in_4_110 = 'b000000010;
logic signed [WIDTH-1:0] w_in_4_111 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_112 = 'b111111010;
logic signed [WIDTH-1:0] w_in_4_113 = 'b111111111;
logic signed [WIDTH-1:0] w_in_4_114 = 'b111111101;
logic signed [WIDTH-1:0] w_in_4_115 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_116 = 'b000000101;
logic signed [WIDTH-1:0] w_in_4_117 = 'b000000011;
logic signed [WIDTH-1:0] w_in_4_118 = 'b111111000;
logic signed [WIDTH-1:0] w_in_4_119 = 'b000001010;
logic signed [WIDTH-1:0] w_in_4_120 = 'b000000101;
logic signed [WIDTH-1:0] w_in_4_121 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_122 = 'b111111111;
logic signed [WIDTH-1:0] w_in_4_123 = 'b000000111;
logic signed [WIDTH-1:0] w_in_4_124 = 'b111110111;
logic signed [WIDTH-1:0] w_in_4_125 = 'b000000000;
logic signed [WIDTH-1:0] w_in_4_126 = 'b111111101;
logic signed [WIDTH-1:0] w_in_4_127 = 'b111111101;
logic signed [WIDTH-1:0] w_in_4_128 = 'b000000011;
logic signed [WIDTH-1:0] w_in_4_129 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_130 = 'b111111111;
logic signed [WIDTH-1:0] w_in_4_131 = 'b000000010;
logic signed [WIDTH-1:0] w_in_4_132 = 'b000000110;
logic signed [WIDTH-1:0] w_in_4_133 = 'b000000011;
logic signed [WIDTH-1:0] w_in_4_134 = 'b111110111;
logic signed [WIDTH-1:0] w_in_4_135 = 'b000000011;
logic signed [WIDTH-1:0] w_in_4_136 = 'b111110100;
logic signed [WIDTH-1:0] w_in_4_137 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_138 = 'b000000000;
logic signed [WIDTH-1:0] w_in_4_139 = 'b111111100;
logic signed [WIDTH-1:0] w_in_4_140 = 'b111111001;
logic signed [WIDTH-1:0] w_in_4_141 = 'b000000011;
logic signed [WIDTH-1:0] w_in_4_142 = 'b000000000;
logic signed [WIDTH-1:0] w_in_4_143 = 'b111110101;
logic signed [WIDTH-1:0] w_in_4_144 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_145 = 'b000000101;
logic signed [WIDTH-1:0] w_in_4_146 = 'b111110100;
logic signed [WIDTH-1:0] w_in_4_147 = 'b111111000;
logic signed [WIDTH-1:0] w_in_4_148 = 'b000000111;
logic signed [WIDTH-1:0] w_in_4_149 = 'b111111010;
logic signed [WIDTH-1:0] w_in_4_150 = 'b000000011;
logic signed [WIDTH-1:0] w_in_4_151 = 'b111111010;
logic signed [WIDTH-1:0] w_in_4_152 = 'b000000011;
logic signed [WIDTH-1:0] w_in_4_153 = 'b111111011;
logic signed [WIDTH-1:0] w_in_4_154 = 'b000001001;
logic signed [WIDTH-1:0] w_in_4_155 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_156 = 'b000000110;
logic signed [WIDTH-1:0] w_in_4_157 = 'b000001001;
logic signed [WIDTH-1:0] w_in_4_158 = 'b111111111;
logic signed [WIDTH-1:0] w_in_4_159 = 'b000000000;
logic signed [WIDTH-1:0] w_in_4_160 = 'b000001011;
logic signed [WIDTH-1:0] w_in_4_161 = 'b111111000;
logic signed [WIDTH-1:0] w_in_4_162 = 'b111111000;
logic signed [WIDTH-1:0] w_in_4_163 = 'b111111100;
logic signed [WIDTH-1:0] w_in_4_164 = 'b000001010;
logic signed [WIDTH-1:0] w_in_4_165 = 'b000001000;
logic signed [WIDTH-1:0] w_in_4_166 = 'b111111011;
logic signed [WIDTH-1:0] w_in_4_167 = 'b111110101;
logic signed [WIDTH-1:0] w_in_4_168 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_169 = 'b111111111;
logic signed [WIDTH-1:0] w_in_4_170 = 'b111111000;
logic signed [WIDTH-1:0] w_in_4_171 = 'b000000001;
logic signed [WIDTH-1:0] w_in_4_172 = 'b111111101;
logic signed [WIDTH-1:0] w_in_4_173 = 'b000000101;
logic signed [WIDTH-1:0] w_in_4_174 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_175 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_176 = 'b111111101;
logic signed [WIDTH-1:0] w_in_4_177 = 'b000000000;
logic signed [WIDTH-1:0] w_in_4_178 = 'b111111000;
logic signed [WIDTH-1:0] w_in_4_179 = 'b111111101;
logic signed [WIDTH-1:0] w_in_4_180 = 'b111111000;
logic signed [WIDTH-1:0] w_in_4_181 = 'b000000111;
logic signed [WIDTH-1:0] w_in_4_182 = 'b111111111;
logic signed [WIDTH-1:0] w_in_4_183 = 'b111111100;
logic signed [WIDTH-1:0] w_in_4_184 = 'b111111101;
logic signed [WIDTH-1:0] w_in_4_185 = 'b000000111;
logic signed [WIDTH-1:0] w_in_4_186 = 'b000001000;
logic signed [WIDTH-1:0] w_in_4_187 = 'b000001010;
logic signed [WIDTH-1:0] w_in_4_188 = 'b000001111;
logic signed [WIDTH-1:0] w_in_4_189 = 'b000001010;
logic signed [WIDTH-1:0] w_in_4_190 = 'b000010001;
logic signed [WIDTH-1:0] w_in_4_191 = 'b000001101;
logic signed [WIDTH-1:0] w_in_4_192 = 'b111110101;
logic signed [WIDTH-1:0] w_in_4_193 = 'b000001000;
logic signed [WIDTH-1:0] w_in_4_194 = 'b000000001;
logic signed [WIDTH-1:0] w_in_4_195 = 'b000001001;
logic signed [WIDTH-1:0] w_in_4_196 = 'b111110110;
logic signed [WIDTH-1:0] w_in_4_197 = 'b000000010;
logic signed [WIDTH-1:0] w_in_4_198 = 'b111110111;
logic signed [WIDTH-1:0] w_in_4_199 = 'b000000101;
logic signed [WIDTH-1:0] w_in_4_200 = 'b111110010;
logic signed [WIDTH-1:0] w_in_4_201 = 'b111110101;
logic signed [WIDTH-1:0] w_in_4_202 = 'b000001001;
logic signed [WIDTH-1:0] w_in_4_203 = 'b111110101;
logic signed [WIDTH-1:0] w_in_4_204 = 'b111110101;
logic signed [WIDTH-1:0] w_in_4_205 = 'b000000101;
logic signed [WIDTH-1:0] w_in_4_206 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_207 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_208 = 'b000001011;
logic signed [WIDTH-1:0] w_in_4_209 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_210 = 'b000000000;
logic signed [WIDTH-1:0] w_in_4_211 = 'b000001101;
logic signed [WIDTH-1:0] w_in_4_212 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_213 = 'b111111000;
logic signed [WIDTH-1:0] w_in_4_214 = 'b111111101;
logic signed [WIDTH-1:0] w_in_4_215 = 'b111111100;
logic signed [WIDTH-1:0] w_in_4_216 = 'b111110110;
logic signed [WIDTH-1:0] w_in_4_217 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_218 = 'b111111000;
logic signed [WIDTH-1:0] w_in_4_219 = 'b111110110;
logic signed [WIDTH-1:0] w_in_4_220 = 'b000001101;
logic signed [WIDTH-1:0] w_in_4_221 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_222 = 'b000000001;
logic signed [WIDTH-1:0] w_in_4_223 = 'b000000111;
logic signed [WIDTH-1:0] w_in_4_224 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_225 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_226 = 'b000000111;
logic signed [WIDTH-1:0] w_in_4_227 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_228 = 'b111110111;
logic signed [WIDTH-1:0] w_in_4_229 = 'b111110110;
logic signed [WIDTH-1:0] w_in_4_230 = 'b000000100;
logic signed [WIDTH-1:0] w_in_4_231 = 'b000000000;
logic signed [WIDTH-1:0] w_in_4_232 = 'b111110100;
logic signed [WIDTH-1:0] w_in_4_233 = 'b111110110;
logic signed [WIDTH-1:0] w_in_4_234 = 'b000001000;
logic signed [WIDTH-1:0] w_in_4_235 = 'b000000001;
logic signed [WIDTH-1:0] w_in_4_236 = 'b000000011;
logic signed [WIDTH-1:0] w_in_4_237 = 'b000001100;
logic signed [WIDTH-1:0] w_in_4_238 = 'b111111111;
logic signed [WIDTH-1:0] w_in_4_239 = 'b000001010;
logic signed [WIDTH-1:0] w_in_4_240 = 'b000000001;
logic signed [WIDTH-1:0] w_in_4_241 = 'b111111111;
logic signed [WIDTH-1:0] w_in_4_242 = 'b111111011;
logic signed [WIDTH-1:0] w_in_4_243 = 'b000000110;
logic signed [WIDTH-1:0] w_in_4_244 = 'b111111110;
logic signed [WIDTH-1:0] w_in_4_245 = 'b111110110;
logic signed [WIDTH-1:0] w_in_4_246 = 'b000001100;
logic signed [WIDTH-1:0] w_in_4_247 = 'b000000010;
logic signed [WIDTH-1:0] w_in_4_248 = 'b111111010;
logic signed [WIDTH-1:0] w_in_4_249 = 'b000000110;
logic signed [WIDTH-1:0] w_in_4_250 = 'b111111011;
logic signed [WIDTH-1:0] w_in_4_251 = 'b000001011;
logic signed [WIDTH-1:0] w_in_4_252 = 'b000001011;
logic signed [WIDTH-1:0] w_in_4_253 = 'b000000011;
logic signed [WIDTH-1:0] w_in_4_254 = 'b000000001;
logic signed [WIDTH-1:0] w_in_4_255 = 'b000001001;
logic signed [WIDTH-1:0] w_in_5_0 = 'b000000011;
logic signed [WIDTH-1:0] w_in_5_1 = 'b000000101;
logic signed [WIDTH-1:0] w_in_5_2 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_3 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_4 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_5 = 'b111111011;
logic signed [WIDTH-1:0] w_in_5_6 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_7 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_8 = 'b111111001;
logic signed [WIDTH-1:0] w_in_5_9 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_10 = 'b000001000;
logic signed [WIDTH-1:0] w_in_5_11 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_12 = 'b000000101;
logic signed [WIDTH-1:0] w_in_5_13 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_14 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_15 = 'b000000110;
logic signed [WIDTH-1:0] w_in_5_16 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_17 = 'b000000111;
logic signed [WIDTH-1:0] w_in_5_18 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_19 = 'b000000101;
logic signed [WIDTH-1:0] w_in_5_20 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_21 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_22 = 'b000000011;
logic signed [WIDTH-1:0] w_in_5_23 = 'b000000011;
logic signed [WIDTH-1:0] w_in_5_24 = 'b111111011;
logic signed [WIDTH-1:0] w_in_5_25 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_26 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_27 = 'b000000011;
logic signed [WIDTH-1:0] w_in_5_28 = 'b000000111;
logic signed [WIDTH-1:0] w_in_5_29 = 'b111111001;
logic signed [WIDTH-1:0] w_in_5_30 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_31 = 'b000000011;
logic signed [WIDTH-1:0] w_in_5_32 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_33 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_34 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_35 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_36 = 'b000001000;
logic signed [WIDTH-1:0] w_in_5_37 = 'b000000011;
logic signed [WIDTH-1:0] w_in_5_38 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_39 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_40 = 'b000000101;
logic signed [WIDTH-1:0] w_in_5_41 = 'b111111010;
logic signed [WIDTH-1:0] w_in_5_42 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_43 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_44 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_45 = 'b111111100;
logic signed [WIDTH-1:0] w_in_5_46 = 'b111111010;
logic signed [WIDTH-1:0] w_in_5_47 = 'b000000111;
logic signed [WIDTH-1:0] w_in_5_48 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_49 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_50 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_51 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_52 = 'b111111001;
logic signed [WIDTH-1:0] w_in_5_53 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_54 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_55 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_56 = 'b000000101;
logic signed [WIDTH-1:0] w_in_5_57 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_58 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_59 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_60 = 'b111111011;
logic signed [WIDTH-1:0] w_in_5_61 = 'b111111010;
logic signed [WIDTH-1:0] w_in_5_62 = 'b111111010;
logic signed [WIDTH-1:0] w_in_5_63 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_64 = 'b111111100;
logic signed [WIDTH-1:0] w_in_5_65 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_66 = 'b000000110;
logic signed [WIDTH-1:0] w_in_5_67 = 'b000000101;
logic signed [WIDTH-1:0] w_in_5_68 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_69 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_70 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_71 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_72 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_73 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_74 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_75 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_76 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_77 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_78 = 'b111111011;
logic signed [WIDTH-1:0] w_in_5_79 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_80 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_81 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_82 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_83 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_84 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_85 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_86 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_87 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_88 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_89 = 'b000000110;
logic signed [WIDTH-1:0] w_in_5_90 = 'b111111010;
logic signed [WIDTH-1:0] w_in_5_91 = 'b111111010;
logic signed [WIDTH-1:0] w_in_5_92 = 'b000000111;
logic signed [WIDTH-1:0] w_in_5_93 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_94 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_95 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_96 = 'b111111100;
logic signed [WIDTH-1:0] w_in_5_97 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_98 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_99 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_100 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_101 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_102 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_103 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_104 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_105 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_106 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_107 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_108 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_109 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_110 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_111 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_112 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_113 = 'b111111001;
logic signed [WIDTH-1:0] w_in_5_114 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_115 = 'b000000101;
logic signed [WIDTH-1:0] w_in_5_116 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_117 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_118 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_119 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_120 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_121 = 'b000000110;
logic signed [WIDTH-1:0] w_in_5_122 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_123 = 'b111111100;
logic signed [WIDTH-1:0] w_in_5_124 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_125 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_126 = 'b000000101;
logic signed [WIDTH-1:0] w_in_5_127 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_128 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_129 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_130 = 'b111111001;
logic signed [WIDTH-1:0] w_in_5_131 = 'b111111100;
logic signed [WIDTH-1:0] w_in_5_132 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_133 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_134 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_135 = 'b111111011;
logic signed [WIDTH-1:0] w_in_5_136 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_137 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_138 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_139 = 'b111111001;
logic signed [WIDTH-1:0] w_in_5_140 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_141 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_142 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_143 = 'b000000011;
logic signed [WIDTH-1:0] w_in_5_144 = 'b111111011;
logic signed [WIDTH-1:0] w_in_5_145 = 'b000000111;
logic signed [WIDTH-1:0] w_in_5_146 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_147 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_148 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_149 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_150 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_151 = 'b000000111;
logic signed [WIDTH-1:0] w_in_5_152 = 'b000000011;
logic signed [WIDTH-1:0] w_in_5_153 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_154 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_155 = 'b111111001;
logic signed [WIDTH-1:0] w_in_5_156 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_157 = 'b000001000;
logic signed [WIDTH-1:0] w_in_5_158 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_159 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_160 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_161 = 'b000000011;
logic signed [WIDTH-1:0] w_in_5_162 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_163 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_164 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_165 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_166 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_167 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_168 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_169 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_170 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_171 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_172 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_173 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_174 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_175 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_176 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_177 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_178 = 'b111111100;
logic signed [WIDTH-1:0] w_in_5_179 = 'b000000011;
logic signed [WIDTH-1:0] w_in_5_180 = 'b000000011;
logic signed [WIDTH-1:0] w_in_5_181 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_182 = 'b111111001;
logic signed [WIDTH-1:0] w_in_5_183 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_184 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_185 = 'b111111011;
logic signed [WIDTH-1:0] w_in_5_186 = 'b111111100;
logic signed [WIDTH-1:0] w_in_5_187 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_188 = 'b000000101;
logic signed [WIDTH-1:0] w_in_5_189 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_190 = 'b000000101;
logic signed [WIDTH-1:0] w_in_5_191 = 'b000001001;
logic signed [WIDTH-1:0] w_in_5_192 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_193 = 'b000001000;
logic signed [WIDTH-1:0] w_in_5_194 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_195 = 'b000000110;
logic signed [WIDTH-1:0] w_in_5_196 = 'b111111010;
logic signed [WIDTH-1:0] w_in_5_197 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_198 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_199 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_200 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_201 = 'b000000101;
logic signed [WIDTH-1:0] w_in_5_202 = 'b111111100;
logic signed [WIDTH-1:0] w_in_5_203 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_204 = 'b111111100;
logic signed [WIDTH-1:0] w_in_5_205 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_206 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_207 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_208 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_209 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_210 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_211 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_212 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_213 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_214 = 'b000000011;
logic signed [WIDTH-1:0] w_in_5_215 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_216 = 'b000000111;
logic signed [WIDTH-1:0] w_in_5_217 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_218 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_219 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_220 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_221 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_222 = 'b111111100;
logic signed [WIDTH-1:0] w_in_5_223 = 'b000001000;
logic signed [WIDTH-1:0] w_in_5_224 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_225 = 'b111111011;
logic signed [WIDTH-1:0] w_in_5_226 = 'b000000010;
logic signed [WIDTH-1:0] w_in_5_227 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_228 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_229 = 'b111111001;
logic signed [WIDTH-1:0] w_in_5_230 = 'b000000011;
logic signed [WIDTH-1:0] w_in_5_231 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_232 = 'b000000000;
logic signed [WIDTH-1:0] w_in_5_233 = 'b000000101;
logic signed [WIDTH-1:0] w_in_5_234 = 'b111111011;
logic signed [WIDTH-1:0] w_in_5_235 = 'b000000001;
logic signed [WIDTH-1:0] w_in_5_236 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_237 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_238 = 'b000000110;
logic signed [WIDTH-1:0] w_in_5_239 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_240 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_241 = 'b111111111;
logic signed [WIDTH-1:0] w_in_5_242 = 'b111111100;
logic signed [WIDTH-1:0] w_in_5_243 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_244 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_245 = 'b111111100;
logic signed [WIDTH-1:0] w_in_5_246 = 'b111111110;
logic signed [WIDTH-1:0] w_in_5_247 = 'b111111001;
logic signed [WIDTH-1:0] w_in_5_248 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_249 = 'b000000100;
logic signed [WIDTH-1:0] w_in_5_250 = 'b111111100;
logic signed [WIDTH-1:0] w_in_5_251 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_252 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_253 = 'b111111101;
logic signed [WIDTH-1:0] w_in_5_254 = 'b111111010;
logic signed [WIDTH-1:0] w_in_5_255 = 'b111111110;
logic signed [WIDTH-1:0] w_in_6_0 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_1 = 'b111111110;
logic signed [WIDTH-1:0] w_in_6_2 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_3 = 'b111111101;
logic signed [WIDTH-1:0] w_in_6_4 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_5 = 'b000000011;
logic signed [WIDTH-1:0] w_in_6_6 = 'b111111100;
logic signed [WIDTH-1:0] w_in_6_7 = 'b111111011;
logic signed [WIDTH-1:0] w_in_6_8 = 'b111111001;
logic signed [WIDTH-1:0] w_in_6_9 = 'b111111101;
logic signed [WIDTH-1:0] w_in_6_10 = 'b111111001;
logic signed [WIDTH-1:0] w_in_6_11 = 'b111111110;
logic signed [WIDTH-1:0] w_in_6_12 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_13 = 'b000000011;
logic signed [WIDTH-1:0] w_in_6_14 = 'b000000001;
logic signed [WIDTH-1:0] w_in_6_15 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_16 = 'b111111100;
logic signed [WIDTH-1:0] w_in_6_17 = 'b111111101;
logic signed [WIDTH-1:0] w_in_6_18 = 'b111111100;
logic signed [WIDTH-1:0] w_in_6_19 = 'b111111011;
logic signed [WIDTH-1:0] w_in_6_20 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_21 = 'b000000011;
logic signed [WIDTH-1:0] w_in_6_22 = 'b000001000;
logic signed [WIDTH-1:0] w_in_6_23 = 'b000000101;
logic signed [WIDTH-1:0] w_in_6_24 = 'b111111001;
logic signed [WIDTH-1:0] w_in_6_25 = 'b111111010;
logic signed [WIDTH-1:0] w_in_6_26 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_27 = 'b111111001;
logic signed [WIDTH-1:0] w_in_6_28 = 'b000000110;
logic signed [WIDTH-1:0] w_in_6_29 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_30 = 'b000000110;
logic signed [WIDTH-1:0] w_in_6_31 = 'b111111100;
logic signed [WIDTH-1:0] w_in_6_32 = 'b111111001;
logic signed [WIDTH-1:0] w_in_6_33 = 'b111111010;
logic signed [WIDTH-1:0] w_in_6_34 = 'b111111100;
logic signed [WIDTH-1:0] w_in_6_35 = 'b111111100;
logic signed [WIDTH-1:0] w_in_6_36 = 'b111111010;
logic signed [WIDTH-1:0] w_in_6_37 = 'b111111011;
logic signed [WIDTH-1:0] w_in_6_38 = 'b111111101;
logic signed [WIDTH-1:0] w_in_6_39 = 'b000000010;
logic signed [WIDTH-1:0] w_in_6_40 = 'b000000001;
logic signed [WIDTH-1:0] w_in_6_41 = 'b111111100;
logic signed [WIDTH-1:0] w_in_6_42 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_43 = 'b111111101;
logic signed [WIDTH-1:0] w_in_6_44 = 'b111111000;
logic signed [WIDTH-1:0] w_in_6_45 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_46 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_47 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_48 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_49 = 'b111111110;
logic signed [WIDTH-1:0] w_in_6_50 = 'b000000101;
logic signed [WIDTH-1:0] w_in_6_51 = 'b111111101;
logic signed [WIDTH-1:0] w_in_6_52 = 'b000000111;
logic signed [WIDTH-1:0] w_in_6_53 = 'b000000100;
logic signed [WIDTH-1:0] w_in_6_54 = 'b000001000;
logic signed [WIDTH-1:0] w_in_6_55 = 'b000000110;
logic signed [WIDTH-1:0] w_in_6_56 = 'b000000011;
logic signed [WIDTH-1:0] w_in_6_57 = 'b111111001;
logic signed [WIDTH-1:0] w_in_6_58 = 'b000000100;
logic signed [WIDTH-1:0] w_in_6_59 = 'b000001110;
logic signed [WIDTH-1:0] w_in_6_60 = 'b000001010;
logic signed [WIDTH-1:0] w_in_6_61 = 'b000001011;
logic signed [WIDTH-1:0] w_in_6_62 = 'b000001101;
logic signed [WIDTH-1:0] w_in_6_63 = 'b000001100;
logic signed [WIDTH-1:0] w_in_6_64 = 'b000000001;
logic signed [WIDTH-1:0] w_in_6_65 = 'b000000001;
logic signed [WIDTH-1:0] w_in_6_66 = 'b000000010;
logic signed [WIDTH-1:0] w_in_6_67 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_68 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_69 = 'b111111011;
logic signed [WIDTH-1:0] w_in_6_70 = 'b000000110;
logic signed [WIDTH-1:0] w_in_6_71 = 'b111111001;
logic signed [WIDTH-1:0] w_in_6_72 = 'b111111010;
logic signed [WIDTH-1:0] w_in_6_73 = 'b111111110;
logic signed [WIDTH-1:0] w_in_6_74 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_75 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_76 = 'b111111100;
logic signed [WIDTH-1:0] w_in_6_77 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_78 = 'b111111100;
logic signed [WIDTH-1:0] w_in_6_79 = 'b111111100;
logic signed [WIDTH-1:0] w_in_6_80 = 'b000000101;
logic signed [WIDTH-1:0] w_in_6_81 = 'b111111011;
logic signed [WIDTH-1:0] w_in_6_82 = 'b000000001;
logic signed [WIDTH-1:0] w_in_6_83 = 'b111111010;
logic signed [WIDTH-1:0] w_in_6_84 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_85 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_86 = 'b000000011;
logic signed [WIDTH-1:0] w_in_6_87 = 'b000000010;
logic signed [WIDTH-1:0] w_in_6_88 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_89 = 'b111111101;
logic signed [WIDTH-1:0] w_in_6_90 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_91 = 'b000000011;
logic signed [WIDTH-1:0] w_in_6_92 = 'b000000001;
logic signed [WIDTH-1:0] w_in_6_93 = 'b111111100;
logic signed [WIDTH-1:0] w_in_6_94 = 'b111111110;
logic signed [WIDTH-1:0] w_in_6_95 = 'b111111001;
logic signed [WIDTH-1:0] w_in_6_96 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_97 = 'b111111000;
logic signed [WIDTH-1:0] w_in_6_98 = 'b111111110;
logic signed [WIDTH-1:0] w_in_6_99 = 'b000000100;
logic signed [WIDTH-1:0] w_in_6_100 = 'b111111100;
logic signed [WIDTH-1:0] w_in_6_101 = 'b111111010;
logic signed [WIDTH-1:0] w_in_6_102 = 'b111110111;
logic signed [WIDTH-1:0] w_in_6_103 = 'b000000101;
logic signed [WIDTH-1:0] w_in_6_104 = 'b111111101;
logic signed [WIDTH-1:0] w_in_6_105 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_106 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_107 = 'b111111101;
logic signed [WIDTH-1:0] w_in_6_108 = 'b000000001;
logic signed [WIDTH-1:0] w_in_6_109 = 'b111111101;
logic signed [WIDTH-1:0] w_in_6_110 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_111 = 'b000000100;
logic signed [WIDTH-1:0] w_in_6_112 = 'b000000010;
logic signed [WIDTH-1:0] w_in_6_113 = 'b000000010;
logic signed [WIDTH-1:0] w_in_6_114 = 'b000000001;
logic signed [WIDTH-1:0] w_in_6_115 = 'b000000001;
logic signed [WIDTH-1:0] w_in_6_116 = 'b111111110;
logic signed [WIDTH-1:0] w_in_6_117 = 'b111111101;
logic signed [WIDTH-1:0] w_in_6_118 = 'b000000010;
logic signed [WIDTH-1:0] w_in_6_119 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_120 = 'b000000001;
logic signed [WIDTH-1:0] w_in_6_121 = 'b111111011;
logic signed [WIDTH-1:0] w_in_6_122 = 'b111111100;
logic signed [WIDTH-1:0] w_in_6_123 = 'b111111110;
logic signed [WIDTH-1:0] w_in_6_124 = 'b000000111;
logic signed [WIDTH-1:0] w_in_6_125 = 'b000000101;
logic signed [WIDTH-1:0] w_in_6_126 = 'b111111110;
logic signed [WIDTH-1:0] w_in_6_127 = 'b000000101;
logic signed [WIDTH-1:0] w_in_6_128 = 'b000000110;
logic signed [WIDTH-1:0] w_in_6_129 = 'b111111110;
logic signed [WIDTH-1:0] w_in_6_130 = 'b000001001;
logic signed [WIDTH-1:0] w_in_6_131 = 'b111111110;
logic signed [WIDTH-1:0] w_in_6_132 = 'b000000101;
logic signed [WIDTH-1:0] w_in_6_133 = 'b000000001;
logic signed [WIDTH-1:0] w_in_6_134 = 'b111111001;
logic signed [WIDTH-1:0] w_in_6_135 = 'b000001001;
logic signed [WIDTH-1:0] w_in_6_136 = 'b000001011;
logic signed [WIDTH-1:0] w_in_6_137 = 'b000000110;
logic signed [WIDTH-1:0] w_in_6_138 = 'b000001000;
logic signed [WIDTH-1:0] w_in_6_139 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_140 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_141 = 'b000000010;
logic signed [WIDTH-1:0] w_in_6_142 = 'b111111110;
logic signed [WIDTH-1:0] w_in_6_143 = 'b111111001;
logic signed [WIDTH-1:0] w_in_6_144 = 'b111111101;
logic signed [WIDTH-1:0] w_in_6_145 = 'b000000101;
logic signed [WIDTH-1:0] w_in_6_146 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_147 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_148 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_149 = 'b111111011;
logic signed [WIDTH-1:0] w_in_6_150 = 'b000001001;
logic signed [WIDTH-1:0] w_in_6_151 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_152 = 'b111111011;
logic signed [WIDTH-1:0] w_in_6_153 = 'b000000011;
logic signed [WIDTH-1:0] w_in_6_154 = 'b111111010;
logic signed [WIDTH-1:0] w_in_6_155 = 'b111111100;
logic signed [WIDTH-1:0] w_in_6_156 = 'b000000110;
logic signed [WIDTH-1:0] w_in_6_157 = 'b000000101;
logic signed [WIDTH-1:0] w_in_6_158 = 'b111111011;
logic signed [WIDTH-1:0] w_in_6_159 = 'b000000101;
logic signed [WIDTH-1:0] w_in_6_160 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_161 = 'b000000011;
logic signed [WIDTH-1:0] w_in_6_162 = 'b000000111;
logic signed [WIDTH-1:0] w_in_6_163 = 'b000001000;
logic signed [WIDTH-1:0] w_in_6_164 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_165 = 'b000000010;
logic signed [WIDTH-1:0] w_in_6_166 = 'b111111000;
logic signed [WIDTH-1:0] w_in_6_167 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_168 = 'b000000100;
logic signed [WIDTH-1:0] w_in_6_169 = 'b111111101;
logic signed [WIDTH-1:0] w_in_6_170 = 'b000001001;
logic signed [WIDTH-1:0] w_in_6_171 = 'b000000010;
logic signed [WIDTH-1:0] w_in_6_172 = 'b000000100;
logic signed [WIDTH-1:0] w_in_6_173 = 'b111111100;
logic signed [WIDTH-1:0] w_in_6_174 = 'b111111001;
logic signed [WIDTH-1:0] w_in_6_175 = 'b000001000;
logic signed [WIDTH-1:0] w_in_6_176 = 'b111111010;
logic signed [WIDTH-1:0] w_in_6_177 = 'b111111100;
logic signed [WIDTH-1:0] w_in_6_178 = 'b000000100;
logic signed [WIDTH-1:0] w_in_6_179 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_180 = 'b000000100;
logic signed [WIDTH-1:0] w_in_6_181 = 'b111110010;
logic signed [WIDTH-1:0] w_in_6_182 = 'b111111110;
logic signed [WIDTH-1:0] w_in_6_183 = 'b000000001;
logic signed [WIDTH-1:0] w_in_6_184 = 'b111111011;
logic signed [WIDTH-1:0] w_in_6_185 = 'b111111110;
logic signed [WIDTH-1:0] w_in_6_186 = 'b111111011;
logic signed [WIDTH-1:0] w_in_6_187 = 'b111111010;
logic signed [WIDTH-1:0] w_in_6_188 = 'b111111110;
logic signed [WIDTH-1:0] w_in_6_189 = 'b111110100;
logic signed [WIDTH-1:0] w_in_6_190 = 'b111110001;
logic signed [WIDTH-1:0] w_in_6_191 = 'b111110000;
logic signed [WIDTH-1:0] w_in_6_192 = 'b111110101;
logic signed [WIDTH-1:0] w_in_6_193 = 'b111110101;
logic signed [WIDTH-1:0] w_in_6_194 = 'b000000011;
logic signed [WIDTH-1:0] w_in_6_195 = 'b111111110;
logic signed [WIDTH-1:0] w_in_6_196 = 'b000000110;
logic signed [WIDTH-1:0] w_in_6_197 = 'b000001000;
logic signed [WIDTH-1:0] w_in_6_198 = 'b111111001;
logic signed [WIDTH-1:0] w_in_6_199 = 'b000000010;
logic signed [WIDTH-1:0] w_in_6_200 = 'b111111011;
logic signed [WIDTH-1:0] w_in_6_201 = 'b111110100;
logic signed [WIDTH-1:0] w_in_6_202 = 'b111111100;
logic signed [WIDTH-1:0] w_in_6_203 = 'b000000101;
logic signed [WIDTH-1:0] w_in_6_204 = 'b000000110;
logic signed [WIDTH-1:0] w_in_6_205 = 'b111111010;
logic signed [WIDTH-1:0] w_in_6_206 = 'b000000110;
logic signed [WIDTH-1:0] w_in_6_207 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_208 = 'b000000001;
logic signed [WIDTH-1:0] w_in_6_209 = 'b111111101;
logic signed [WIDTH-1:0] w_in_6_210 = 'b000000001;
logic signed [WIDTH-1:0] w_in_6_211 = 'b000000111;
logic signed [WIDTH-1:0] w_in_6_212 = 'b111111100;
logic signed [WIDTH-1:0] w_in_6_213 = 'b111111101;
logic signed [WIDTH-1:0] w_in_6_214 = 'b000001000;
logic signed [WIDTH-1:0] w_in_6_215 = 'b111111101;
logic signed [WIDTH-1:0] w_in_6_216 = 'b000000111;
logic signed [WIDTH-1:0] w_in_6_217 = 'b000000011;
logic signed [WIDTH-1:0] w_in_6_218 = 'b000000100;
logic signed [WIDTH-1:0] w_in_6_219 = 'b111111110;
logic signed [WIDTH-1:0] w_in_6_220 = 'b000000110;
logic signed [WIDTH-1:0] w_in_6_221 = 'b000001001;
logic signed [WIDTH-1:0] w_in_6_222 = 'b000000110;
logic signed [WIDTH-1:0] w_in_6_223 = 'b000000011;
logic signed [WIDTH-1:0] w_in_6_224 = 'b111111011;
logic signed [WIDTH-1:0] w_in_6_225 = 'b111111101;
logic signed [WIDTH-1:0] w_in_6_226 = 'b111110100;
logic signed [WIDTH-1:0] w_in_6_227 = 'b111111010;
logic signed [WIDTH-1:0] w_in_6_228 = 'b000001000;
logic signed [WIDTH-1:0] w_in_6_229 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_230 = 'b000000110;
logic signed [WIDTH-1:0] w_in_6_231 = 'b111110111;
logic signed [WIDTH-1:0] w_in_6_232 = 'b000000000;
logic signed [WIDTH-1:0] w_in_6_233 = 'b111111000;
logic signed [WIDTH-1:0] w_in_6_234 = 'b111110111;
logic signed [WIDTH-1:0] w_in_6_235 = 'b111110111;
logic signed [WIDTH-1:0] w_in_6_236 = 'b111111011;
logic signed [WIDTH-1:0] w_in_6_237 = 'b000000001;
logic signed [WIDTH-1:0] w_in_6_238 = 'b000010010;
logic signed [WIDTH-1:0] w_in_6_239 = 'b111111011;
logic signed [WIDTH-1:0] w_in_6_240 = 'b111111111;
logic signed [WIDTH-1:0] w_in_6_241 = 'b111111011;
logic signed [WIDTH-1:0] w_in_6_242 = 'b111111000;
logic signed [WIDTH-1:0] w_in_6_243 = 'b000001100;
logic signed [WIDTH-1:0] w_in_6_244 = 'b111110111;
logic signed [WIDTH-1:0] w_in_6_245 = 'b000000011;
logic signed [WIDTH-1:0] w_in_6_246 = 'b000001001;
logic signed [WIDTH-1:0] w_in_6_247 = 'b000000001;
logic signed [WIDTH-1:0] w_in_6_248 = 'b000010010;
logic signed [WIDTH-1:0] w_in_6_249 = 'b000000010;
logic signed [WIDTH-1:0] w_in_6_250 = 'b000010011;
logic signed [WIDTH-1:0] w_in_6_251 = 'b000000011;
logic signed [WIDTH-1:0] w_in_6_252 = 'b111111000;
logic signed [WIDTH-1:0] w_in_6_253 = 'b000001001;
logic signed [WIDTH-1:0] w_in_6_254 = 'b000001100;
logic signed [WIDTH-1:0] w_in_6_255 = 'b111111000;
logic signed [WIDTH-1:0] w_in_7_0 = 'b111111100;
logic signed [WIDTH-1:0] w_in_7_1 = 'b000000010;
logic signed [WIDTH-1:0] w_in_7_2 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_3 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_4 = 'b111111111;
logic signed [WIDTH-1:0] w_in_7_5 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_6 = 'b111111001;
logic signed [WIDTH-1:0] w_in_7_7 = 'b111111100;
logic signed [WIDTH-1:0] w_in_7_8 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_9 = 'b000000101;
logic signed [WIDTH-1:0] w_in_7_10 = 'b000000010;
logic signed [WIDTH-1:0] w_in_7_11 = 'b000000111;
logic signed [WIDTH-1:0] w_in_7_12 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_13 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_14 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_15 = 'b000000010;
logic signed [WIDTH-1:0] w_in_7_16 = 'b111111111;
logic signed [WIDTH-1:0] w_in_7_17 = 'b000000101;
logic signed [WIDTH-1:0] w_in_7_18 = 'b000001000;
logic signed [WIDTH-1:0] w_in_7_19 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_20 = 'b111111111;
logic signed [WIDTH-1:0] w_in_7_21 = 'b000000001;
logic signed [WIDTH-1:0] w_in_7_22 = 'b000000110;
logic signed [WIDTH-1:0] w_in_7_23 = 'b000000001;
logic signed [WIDTH-1:0] w_in_7_24 = 'b000000000;
logic signed [WIDTH-1:0] w_in_7_25 = 'b111111111;
logic signed [WIDTH-1:0] w_in_7_26 = 'b111111001;
logic signed [WIDTH-1:0] w_in_7_27 = 'b000000010;
logic signed [WIDTH-1:0] w_in_7_28 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_29 = 'b000000000;
logic signed [WIDTH-1:0] w_in_7_30 = 'b000000101;
logic signed [WIDTH-1:0] w_in_7_31 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_32 = 'b111111111;
logic signed [WIDTH-1:0] w_in_7_33 = 'b111111011;
logic signed [WIDTH-1:0] w_in_7_34 = 'b111111010;
logic signed [WIDTH-1:0] w_in_7_35 = 'b111111101;
logic signed [WIDTH-1:0] w_in_7_36 = 'b111111101;
logic signed [WIDTH-1:0] w_in_7_37 = 'b111110110;
logic signed [WIDTH-1:0] w_in_7_38 = 'b000000010;
logic signed [WIDTH-1:0] w_in_7_39 = 'b111111111;
logic signed [WIDTH-1:0] w_in_7_40 = 'b111111111;
logic signed [WIDTH-1:0] w_in_7_41 = 'b000000111;
logic signed [WIDTH-1:0] w_in_7_42 = 'b111111011;
logic signed [WIDTH-1:0] w_in_7_43 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_44 = 'b000000000;
logic signed [WIDTH-1:0] w_in_7_45 = 'b111111100;
logic signed [WIDTH-1:0] w_in_7_46 = 'b111111011;
logic signed [WIDTH-1:0] w_in_7_47 = 'b000000101;
logic signed [WIDTH-1:0] w_in_7_48 = 'b000000010;
logic signed [WIDTH-1:0] w_in_7_49 = 'b000001001;
logic signed [WIDTH-1:0] w_in_7_50 = 'b000000000;
logic signed [WIDTH-1:0] w_in_7_51 = 'b000000010;
logic signed [WIDTH-1:0] w_in_7_52 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_53 = 'b111111010;
logic signed [WIDTH-1:0] w_in_7_54 = 'b111111001;
logic signed [WIDTH-1:0] w_in_7_55 = 'b111111101;
logic signed [WIDTH-1:0] w_in_7_56 = 'b000000111;
logic signed [WIDTH-1:0] w_in_7_57 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_58 = 'b000001000;
logic signed [WIDTH-1:0] w_in_7_59 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_60 = 'b111110111;
logic signed [WIDTH-1:0] w_in_7_61 = 'b111110010;
logic signed [WIDTH-1:0] w_in_7_62 = 'b111110000;
logic signed [WIDTH-1:0] w_in_7_63 = 'b000000011;
logic signed [WIDTH-1:0] w_in_7_64 = 'b000000110;
logic signed [WIDTH-1:0] w_in_7_65 = 'b000000010;
logic signed [WIDTH-1:0] w_in_7_66 = 'b000000001;
logic signed [WIDTH-1:0] w_in_7_67 = 'b000000000;
logic signed [WIDTH-1:0] w_in_7_68 = 'b000000001;
logic signed [WIDTH-1:0] w_in_7_69 = 'b000000101;
logic signed [WIDTH-1:0] w_in_7_70 = 'b111111010;
logic signed [WIDTH-1:0] w_in_7_71 = 'b111111011;
logic signed [WIDTH-1:0] w_in_7_72 = 'b000000000;
logic signed [WIDTH-1:0] w_in_7_73 = 'b000001000;
logic signed [WIDTH-1:0] w_in_7_74 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_75 = 'b111111000;
logic signed [WIDTH-1:0] w_in_7_76 = 'b111111011;
logic signed [WIDTH-1:0] w_in_7_77 = 'b000000101;
logic signed [WIDTH-1:0] w_in_7_78 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_79 = 'b000000110;
logic signed [WIDTH-1:0] w_in_7_80 = 'b111111000;
logic signed [WIDTH-1:0] w_in_7_81 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_82 = 'b000001001;
logic signed [WIDTH-1:0] w_in_7_83 = 'b111111011;
logic signed [WIDTH-1:0] w_in_7_84 = 'b111111011;
logic signed [WIDTH-1:0] w_in_7_85 = 'b111111001;
logic signed [WIDTH-1:0] w_in_7_86 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_87 = 'b000001010;
logic signed [WIDTH-1:0] w_in_7_88 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_89 = 'b111111100;
logic signed [WIDTH-1:0] w_in_7_90 = 'b111111101;
logic signed [WIDTH-1:0] w_in_7_91 = 'b111111100;
logic signed [WIDTH-1:0] w_in_7_92 = 'b111111101;
logic signed [WIDTH-1:0] w_in_7_93 = 'b111111010;
logic signed [WIDTH-1:0] w_in_7_94 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_95 = 'b111111010;
logic signed [WIDTH-1:0] w_in_7_96 = 'b000000101;
logic signed [WIDTH-1:0] w_in_7_97 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_98 = 'b111111100;
logic signed [WIDTH-1:0] w_in_7_99 = 'b000000101;
logic signed [WIDTH-1:0] w_in_7_100 = 'b111110111;
logic signed [WIDTH-1:0] w_in_7_101 = 'b000000001;
logic signed [WIDTH-1:0] w_in_7_102 = 'b000000000;
logic signed [WIDTH-1:0] w_in_7_103 = 'b111111100;
logic signed [WIDTH-1:0] w_in_7_104 = 'b000000110;
logic signed [WIDTH-1:0] w_in_7_105 = 'b000000011;
logic signed [WIDTH-1:0] w_in_7_106 = 'b000000111;
logic signed [WIDTH-1:0] w_in_7_107 = 'b000000110;
logic signed [WIDTH-1:0] w_in_7_108 = 'b000000000;
logic signed [WIDTH-1:0] w_in_7_109 = 'b000000111;
logic signed [WIDTH-1:0] w_in_7_110 = 'b000000010;
logic signed [WIDTH-1:0] w_in_7_111 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_112 = 'b111111010;
logic signed [WIDTH-1:0] w_in_7_113 = 'b111111111;
logic signed [WIDTH-1:0] w_in_7_114 = 'b111111101;
logic signed [WIDTH-1:0] w_in_7_115 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_116 = 'b000000101;
logic signed [WIDTH-1:0] w_in_7_117 = 'b000000011;
logic signed [WIDTH-1:0] w_in_7_118 = 'b111111000;
logic signed [WIDTH-1:0] w_in_7_119 = 'b000001010;
logic signed [WIDTH-1:0] w_in_7_120 = 'b000000101;
logic signed [WIDTH-1:0] w_in_7_121 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_122 = 'b111111111;
logic signed [WIDTH-1:0] w_in_7_123 = 'b000000111;
logic signed [WIDTH-1:0] w_in_7_124 = 'b111110111;
logic signed [WIDTH-1:0] w_in_7_125 = 'b000000000;
logic signed [WIDTH-1:0] w_in_7_126 = 'b111111101;
logic signed [WIDTH-1:0] w_in_7_127 = 'b111111101;
logic signed [WIDTH-1:0] w_in_7_128 = 'b000000011;
logic signed [WIDTH-1:0] w_in_7_129 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_130 = 'b111111111;
logic signed [WIDTH-1:0] w_in_7_131 = 'b000000010;
logic signed [WIDTH-1:0] w_in_7_132 = 'b000000110;
logic signed [WIDTH-1:0] w_in_7_133 = 'b000000011;
logic signed [WIDTH-1:0] w_in_7_134 = 'b111110111;
logic signed [WIDTH-1:0] w_in_7_135 = 'b000000011;
logic signed [WIDTH-1:0] w_in_7_136 = 'b111110100;
logic signed [WIDTH-1:0] w_in_7_137 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_138 = 'b000000000;
logic signed [WIDTH-1:0] w_in_7_139 = 'b111111100;
logic signed [WIDTH-1:0] w_in_7_140 = 'b111111001;
logic signed [WIDTH-1:0] w_in_7_141 = 'b000000011;
logic signed [WIDTH-1:0] w_in_7_142 = 'b000000000;
logic signed [WIDTH-1:0] w_in_7_143 = 'b111110101;
logic signed [WIDTH-1:0] w_in_7_144 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_145 = 'b000000101;
logic signed [WIDTH-1:0] w_in_7_146 = 'b111110100;
logic signed [WIDTH-1:0] w_in_7_147 = 'b111111000;
logic signed [WIDTH-1:0] w_in_7_148 = 'b000000111;
logic signed [WIDTH-1:0] w_in_7_149 = 'b111111010;
logic signed [WIDTH-1:0] w_in_7_150 = 'b000000011;
logic signed [WIDTH-1:0] w_in_7_151 = 'b111111010;
logic signed [WIDTH-1:0] w_in_7_152 = 'b000000011;
logic signed [WIDTH-1:0] w_in_7_153 = 'b111111011;
logic signed [WIDTH-1:0] w_in_7_154 = 'b000001001;
logic signed [WIDTH-1:0] w_in_7_155 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_156 = 'b000000110;
logic signed [WIDTH-1:0] w_in_7_157 = 'b000001001;
logic signed [WIDTH-1:0] w_in_7_158 = 'b111111111;
logic signed [WIDTH-1:0] w_in_7_159 = 'b000000000;
logic signed [WIDTH-1:0] w_in_7_160 = 'b000001011;
logic signed [WIDTH-1:0] w_in_7_161 = 'b111111000;
logic signed [WIDTH-1:0] w_in_7_162 = 'b111111000;
logic signed [WIDTH-1:0] w_in_7_163 = 'b111111100;
logic signed [WIDTH-1:0] w_in_7_164 = 'b000001010;
logic signed [WIDTH-1:0] w_in_7_165 = 'b000001000;
logic signed [WIDTH-1:0] w_in_7_166 = 'b111111011;
logic signed [WIDTH-1:0] w_in_7_167 = 'b111110101;
logic signed [WIDTH-1:0] w_in_7_168 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_169 = 'b111111111;
logic signed [WIDTH-1:0] w_in_7_170 = 'b111111000;
logic signed [WIDTH-1:0] w_in_7_171 = 'b000000001;
logic signed [WIDTH-1:0] w_in_7_172 = 'b111111101;
logic signed [WIDTH-1:0] w_in_7_173 = 'b000000101;
logic signed [WIDTH-1:0] w_in_7_174 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_175 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_176 = 'b111111101;
logic signed [WIDTH-1:0] w_in_7_177 = 'b000000000;
logic signed [WIDTH-1:0] w_in_7_178 = 'b111111000;
logic signed [WIDTH-1:0] w_in_7_179 = 'b111111101;
logic signed [WIDTH-1:0] w_in_7_180 = 'b111111000;
logic signed [WIDTH-1:0] w_in_7_181 = 'b000000111;
logic signed [WIDTH-1:0] w_in_7_182 = 'b111111111;
logic signed [WIDTH-1:0] w_in_7_183 = 'b111111100;
logic signed [WIDTH-1:0] w_in_7_184 = 'b111111101;
logic signed [WIDTH-1:0] w_in_7_185 = 'b000000111;
logic signed [WIDTH-1:0] w_in_7_186 = 'b000001000;
logic signed [WIDTH-1:0] w_in_7_187 = 'b000001010;
logic signed [WIDTH-1:0] w_in_7_188 = 'b000001111;
logic signed [WIDTH-1:0] w_in_7_189 = 'b000001010;
logic signed [WIDTH-1:0] w_in_7_190 = 'b000010001;
logic signed [WIDTH-1:0] w_in_7_191 = 'b000001101;
logic signed [WIDTH-1:0] w_in_7_192 = 'b111110101;
logic signed [WIDTH-1:0] w_in_7_193 = 'b000001000;
logic signed [WIDTH-1:0] w_in_7_194 = 'b000000001;
logic signed [WIDTH-1:0] w_in_7_195 = 'b000001001;
logic signed [WIDTH-1:0] w_in_7_196 = 'b111110110;
logic signed [WIDTH-1:0] w_in_7_197 = 'b000000010;
logic signed [WIDTH-1:0] w_in_7_198 = 'b111110111;
logic signed [WIDTH-1:0] w_in_7_199 = 'b000000101;
logic signed [WIDTH-1:0] w_in_7_200 = 'b111110010;
logic signed [WIDTH-1:0] w_in_7_201 = 'b111110101;
logic signed [WIDTH-1:0] w_in_7_202 = 'b000001001;
logic signed [WIDTH-1:0] w_in_7_203 = 'b111110101;
logic signed [WIDTH-1:0] w_in_7_204 = 'b111110101;
logic signed [WIDTH-1:0] w_in_7_205 = 'b000000101;
logic signed [WIDTH-1:0] w_in_7_206 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_207 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_208 = 'b000001011;
logic signed [WIDTH-1:0] w_in_7_209 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_210 = 'b000000000;
logic signed [WIDTH-1:0] w_in_7_211 = 'b000001101;
logic signed [WIDTH-1:0] w_in_7_212 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_213 = 'b111111000;
logic signed [WIDTH-1:0] w_in_7_214 = 'b111111101;
logic signed [WIDTH-1:0] w_in_7_215 = 'b111111100;
logic signed [WIDTH-1:0] w_in_7_216 = 'b111110110;
logic signed [WIDTH-1:0] w_in_7_217 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_218 = 'b111111000;
logic signed [WIDTH-1:0] w_in_7_219 = 'b111110110;
logic signed [WIDTH-1:0] w_in_7_220 = 'b000001101;
logic signed [WIDTH-1:0] w_in_7_221 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_222 = 'b000000001;
logic signed [WIDTH-1:0] w_in_7_223 = 'b000000111;
logic signed [WIDTH-1:0] w_in_7_224 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_225 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_226 = 'b000000111;
logic signed [WIDTH-1:0] w_in_7_227 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_228 = 'b111110111;
logic signed [WIDTH-1:0] w_in_7_229 = 'b111110110;
logic signed [WIDTH-1:0] w_in_7_230 = 'b000000100;
logic signed [WIDTH-1:0] w_in_7_231 = 'b000000000;
logic signed [WIDTH-1:0] w_in_7_232 = 'b111110100;
logic signed [WIDTH-1:0] w_in_7_233 = 'b111110110;
logic signed [WIDTH-1:0] w_in_7_234 = 'b000001000;
logic signed [WIDTH-1:0] w_in_7_235 = 'b000000001;
logic signed [WIDTH-1:0] w_in_7_236 = 'b000000011;
logic signed [WIDTH-1:0] w_in_7_237 = 'b000001100;
logic signed [WIDTH-1:0] w_in_7_238 = 'b111111111;
logic signed [WIDTH-1:0] w_in_7_239 = 'b000001010;
logic signed [WIDTH-1:0] w_in_7_240 = 'b000000001;
logic signed [WIDTH-1:0] w_in_7_241 = 'b111111111;
logic signed [WIDTH-1:0] w_in_7_242 = 'b111111011;
logic signed [WIDTH-1:0] w_in_7_243 = 'b000000110;
logic signed [WIDTH-1:0] w_in_7_244 = 'b111111110;
logic signed [WIDTH-1:0] w_in_7_245 = 'b111110110;
logic signed [WIDTH-1:0] w_in_7_246 = 'b000001100;
logic signed [WIDTH-1:0] w_in_7_247 = 'b000000010;
logic signed [WIDTH-1:0] w_in_7_248 = 'b111111010;
logic signed [WIDTH-1:0] w_in_7_249 = 'b000000110;
logic signed [WIDTH-1:0] w_in_7_250 = 'b111111011;
logic signed [WIDTH-1:0] w_in_7_251 = 'b000001011;
logic signed [WIDTH-1:0] w_in_7_252 = 'b000001011;
logic signed [WIDTH-1:0] w_in_7_253 = 'b000000011;
logic signed [WIDTH-1:0] w_in_7_254 = 'b000000001;
logic signed [WIDTH-1:0] w_in_7_255 = 'b000001001;

// Recurrent weights (h×h for each gate)
logic signed [WIDTH-1:0] w_hr_0_0 = 'b000000000;
logic signed [WIDTH-1:0] w_hr_0_1 = 'b000000001;
logic signed [WIDTH-1:0] w_hr_0_2 = 'b000000010;
logic signed [WIDTH-1:0] w_hr_0_3 = 'b111111011;
logic signed [WIDTH-1:0] w_hr_0_4 = 'b000001001;
logic signed [WIDTH-1:0] w_hr_0_5 = 'b000001001;
logic signed [WIDTH-1:0] w_hr_0_6 = 'b000001001;
logic signed [WIDTH-1:0] w_hr_0_7 = 'b111110111;
logic signed [WIDTH-1:0] w_hr_1_0 = 'b000001000;
logic signed [WIDTH-1:0] w_hr_1_1 = 'b000001001;
logic signed [WIDTH-1:0] w_hr_1_2 = 'b111111100;
logic signed [WIDTH-1:0] w_hr_1_3 = 'b111111011;
logic signed [WIDTH-1:0] w_hr_1_4 = 'b000000100;
logic signed [WIDTH-1:0] w_hr_1_5 = 'b000000101;
logic signed [WIDTH-1:0] w_hr_1_6 = 'b000001011;
logic signed [WIDTH-1:0] w_hr_1_7 = 'b111111000;
logic signed [WIDTH-1:0] w_hr_2_0 = 'b000000111;
logic signed [WIDTH-1:0] w_hr_2_1 = 'b000000100;
logic signed [WIDTH-1:0] w_hr_2_2 = 'b111111101;
logic signed [WIDTH-1:0] w_hr_2_3 = 'b000000100;
logic signed [WIDTH-1:0] w_hr_2_4 = 'b000001101;
logic signed [WIDTH-1:0] w_hr_2_5 = 'b111110100;
logic signed [WIDTH-1:0] w_hr_2_6 = 'b000000000;
logic signed [WIDTH-1:0] w_hr_2_7 = 'b000001001;
logic signed [WIDTH-1:0] w_hr_3_0 = 'b000000111;
logic signed [WIDTH-1:0] w_hr_3_1 = 'b000000000;
logic signed [WIDTH-1:0] w_hr_3_2 = 'b111110000;
logic signed [WIDTH-1:0] w_hr_3_3 = 'b000001110;
logic signed [WIDTH-1:0] w_hr_3_4 = 'b000001100;
logic signed [WIDTH-1:0] w_hr_3_5 = 'b000000100;
logic signed [WIDTH-1:0] w_hr_3_6 = 'b111110111;
logic signed [WIDTH-1:0] w_hr_3_7 = 'b000010101;
logic signed [WIDTH-1:0] w_hr_4_0 = 'b111111111;
logic signed [WIDTH-1:0] w_hr_4_1 = 'b111111110;
logic signed [WIDTH-1:0] w_hr_4_2 = 'b000000101;
logic signed [WIDTH-1:0] w_hr_4_3 = 'b111111010;
logic signed [WIDTH-1:0] w_hr_4_4 = 'b111111010;
logic signed [WIDTH-1:0] w_hr_4_5 = 'b111111111;
logic signed [WIDTH-1:0] w_hr_4_6 = 'b000010111;
logic signed [WIDTH-1:0] w_hr_4_7 = 'b111110100;
logic signed [WIDTH-1:0] w_hr_5_0 = 'b111111111;
logic signed [WIDTH-1:0] w_hr_5_1 = 'b000001110;
logic signed [WIDTH-1:0] w_hr_5_2 = 'b000010100;
logic signed [WIDTH-1:0] w_hr_5_3 = 'b111110010;
logic signed [WIDTH-1:0] w_hr_5_4 = 'b111111011;
logic signed [WIDTH-1:0] w_hr_5_5 = 'b111110110;
logic signed [WIDTH-1:0] w_hr_5_6 = 'b111111001;
logic signed [WIDTH-1:0] w_hr_5_7 = 'b000001010;
logic signed [WIDTH-1:0] w_hr_6_0 = 'b000000000;
logic signed [WIDTH-1:0] w_hr_6_1 = 'b000000001;
logic signed [WIDTH-1:0] w_hr_6_2 = 'b000000010;
logic signed [WIDTH-1:0] w_hr_6_3 = 'b111111011;
logic signed [WIDTH-1:0] w_hr_6_4 = 'b000001001;
logic signed [WIDTH-1:0] w_hr_6_5 = 'b000001001;
logic signed [WIDTH-1:0] w_hr_6_6 = 'b000001001;
logic signed [WIDTH-1:0] w_hr_6_7 = 'b111110111;
logic signed [WIDTH-1:0] w_hr_7_0 = 'b000001000;
logic signed [WIDTH-1:0] w_hr_7_1 = 'b000001001;
logic signed [WIDTH-1:0] w_hr_7_2 = 'b111111100;
logic signed [WIDTH-1:0] w_hr_7_3 = 'b111111011;
logic signed [WIDTH-1:0] w_hr_7_4 = 'b000000100;
logic signed [WIDTH-1:0] w_hr_7_5 = 'b000000101;
logic signed [WIDTH-1:0] w_hr_7_6 = 'b000001011;
logic signed [WIDTH-1:0] w_hr_7_7 = 'b111111000;

logic signed [WIDTH-1:0] w_hz_0_0 = 'b000000111;
logic signed [WIDTH-1:0] w_hz_0_1 = 'b000000100;
logic signed [WIDTH-1:0] w_hz_0_2 = 'b111111101;
logic signed [WIDTH-1:0] w_hz_0_3 = 'b000000100;
logic signed [WIDTH-1:0] w_hz_0_4 = 'b000001101;
logic signed [WIDTH-1:0] w_hz_0_5 = 'b111110100;
logic signed [WIDTH-1:0] w_hz_0_6 = 'b000000000;
logic signed [WIDTH-1:0] w_hz_0_7 = 'b000001001;
logic signed [WIDTH-1:0] w_hz_1_0 = 'b000000111;
logic signed [WIDTH-1:0] w_hz_1_1 = 'b000000000;
logic signed [WIDTH-1:0] w_hz_1_2 = 'b111110000;
logic signed [WIDTH-1:0] w_hz_1_3 = 'b000001110;
logic signed [WIDTH-1:0] w_hz_1_4 = 'b000001100;
logic signed [WIDTH-1:0] w_hz_1_5 = 'b000000100;
logic signed [WIDTH-1:0] w_hz_1_6 = 'b111110111;
logic signed [WIDTH-1:0] w_hz_1_7 = 'b000010101;
logic signed [WIDTH-1:0] w_hz_2_0 = 'b111111111;
logic signed [WIDTH-1:0] w_hz_2_1 = 'b111111110;
logic signed [WIDTH-1:0] w_hz_2_2 = 'b000000101;
logic signed [WIDTH-1:0] w_hz_2_3 = 'b111111010;
logic signed [WIDTH-1:0] w_hz_2_4 = 'b111111010;
logic signed [WIDTH-1:0] w_hz_2_5 = 'b111111111;
logic signed [WIDTH-1:0] w_hz_2_6 = 'b000010111;
logic signed [WIDTH-1:0] w_hz_2_7 = 'b111110100;
logic signed [WIDTH-1:0] w_hz_3_0 = 'b111111111;
logic signed [WIDTH-1:0] w_hz_3_1 = 'b000001110;
logic signed [WIDTH-1:0] w_hz_3_2 = 'b000010100;
logic signed [WIDTH-1:0] w_hz_3_3 = 'b111110010;
logic signed [WIDTH-1:0] w_hz_3_4 = 'b111111011;
logic signed [WIDTH-1:0] w_hz_3_5 = 'b111110110;
logic signed [WIDTH-1:0] w_hz_3_6 = 'b111111001;
logic signed [WIDTH-1:0] w_hz_3_7 = 'b000001010;
logic signed [WIDTH-1:0] w_hz_4_0 = 'b000000000;
logic signed [WIDTH-1:0] w_hz_4_1 = 'b000000001;
logic signed [WIDTH-1:0] w_hz_4_2 = 'b000000010;
logic signed [WIDTH-1:0] w_hz_4_3 = 'b111111011;
logic signed [WIDTH-1:0] w_hz_4_4 = 'b000001001;
logic signed [WIDTH-1:0] w_hz_4_5 = 'b000001001;
logic signed [WIDTH-1:0] w_hz_4_6 = 'b000001001;
logic signed [WIDTH-1:0] w_hz_4_7 = 'b111110111;
logic signed [WIDTH-1:0] w_hz_5_0 = 'b000001000;
logic signed [WIDTH-1:0] w_hz_5_1 = 'b000001001;
logic signed [WIDTH-1:0] w_hz_5_2 = 'b111111100;
logic signed [WIDTH-1:0] w_hz_5_3 = 'b111111011;
logic signed [WIDTH-1:0] w_hz_5_4 = 'b000000100;
logic signed [WIDTH-1:0] w_hz_5_5 = 'b000000101;
logic signed [WIDTH-1:0] w_hz_5_6 = 'b000001011;
logic signed [WIDTH-1:0] w_hz_5_7 = 'b111111000;
logic signed [WIDTH-1:0] w_hz_6_0 = 'b000000111;
logic signed [WIDTH-1:0] w_hz_6_1 = 'b000000100;
logic signed [WIDTH-1:0] w_hz_6_2 = 'b111111101;
logic signed [WIDTH-1:0] w_hz_6_3 = 'b000000100;
logic signed [WIDTH-1:0] w_hz_6_4 = 'b000001101;
logic signed [WIDTH-1:0] w_hz_6_5 = 'b111110100;
logic signed [WIDTH-1:0] w_hz_6_6 = 'b000000000;
logic signed [WIDTH-1:0] w_hz_6_7 = 'b000001001;
logic signed [WIDTH-1:0] w_hz_7_0 = 'b000000111;
logic signed [WIDTH-1:0] w_hz_7_1 = 'b000000000;
logic signed [WIDTH-1:0] w_hz_7_2 = 'b111110000;
logic signed [WIDTH-1:0] w_hz_7_3 = 'b000001110;
logic signed [WIDTH-1:0] w_hz_7_4 = 'b000001100;
logic signed [WIDTH-1:0] w_hz_7_5 = 'b000000100;
logic signed [WIDTH-1:0] w_hz_7_6 = 'b111110111;
logic signed [WIDTH-1:0] w_hz_7_7 = 'b000010101;

logic signed [WIDTH-1:0] w_hn_0_0 = 'b111111111;
logic signed [WIDTH-1:0] w_hn_0_1 = 'b111111110;
logic signed [WIDTH-1:0] w_hn_0_2 = 'b000000101;
logic signed [WIDTH-1:0] w_hn_0_3 = 'b111111010;
logic signed [WIDTH-1:0] w_hn_0_4 = 'b111111010;
logic signed [WIDTH-1:0] w_hn_0_5 = 'b111111111;
logic signed [WIDTH-1:0] w_hn_0_6 = 'b000010111;
logic signed [WIDTH-1:0] w_hn_0_7 = 'b111110100;
logic signed [WIDTH-1:0] w_hn_1_0 = 'b111111111;
logic signed [WIDTH-1:0] w_hn_1_1 = 'b000001110;
logic signed [WIDTH-1:0] w_hn_1_2 = 'b000010100;
logic signed [WIDTH-1:0] w_hn_1_3 = 'b111110010;
logic signed [WIDTH-1:0] w_hn_1_4 = 'b111111011;
logic signed [WIDTH-1:0] w_hn_1_5 = 'b111110110;
logic signed [WIDTH-1:0] w_hn_1_6 = 'b111111001;
logic signed [WIDTH-1:0] w_hn_1_7 = 'b000001010;
logic signed [WIDTH-1:0] w_hn_2_0 = 'b000000000;
logic signed [WIDTH-1:0] w_hn_2_1 = 'b000000001;
logic signed [WIDTH-1:0] w_hn_2_2 = 'b000000010;
logic signed [WIDTH-1:0] w_hn_2_3 = 'b111111011;
logic signed [WIDTH-1:0] w_hn_2_4 = 'b000001001;
logic signed [WIDTH-1:0] w_hn_2_5 = 'b000001001;
logic signed [WIDTH-1:0] w_hn_2_6 = 'b000001001;
logic signed [WIDTH-1:0] w_hn_2_7 = 'b111110111;
logic signed [WIDTH-1:0] w_hn_3_0 = 'b000001000;
logic signed [WIDTH-1:0] w_hn_3_1 = 'b000001001;
logic signed [WIDTH-1:0] w_hn_3_2 = 'b111111100;
logic signed [WIDTH-1:0] w_hn_3_3 = 'b111111011;
logic signed [WIDTH-1:0] w_hn_3_4 = 'b000000100;
logic signed [WIDTH-1:0] w_hn_3_5 = 'b000000101;
logic signed [WIDTH-1:0] w_hn_3_6 = 'b000001011;
logic signed [WIDTH-1:0] w_hn_3_7 = 'b111111000;
logic signed [WIDTH-1:0] w_hn_4_0 = 'b000000111;
logic signed [WIDTH-1:0] w_hn_4_1 = 'b000000100;
logic signed [WIDTH-1:0] w_hn_4_2 = 'b111111101;
logic signed [WIDTH-1:0] w_hn_4_3 = 'b000000100;
logic signed [WIDTH-1:0] w_hn_4_4 = 'b000001101;
logic signed [WIDTH-1:0] w_hn_4_5 = 'b111110100;
logic signed [WIDTH-1:0] w_hn_4_6 = 'b000000000;
logic signed [WIDTH-1:0] w_hn_4_7 = 'b000001001;
logic signed [WIDTH-1:0] w_hn_5_0 = 'b000000111;
logic signed [WIDTH-1:0] w_hn_5_1 = 'b000000000;
logic signed [WIDTH-1:0] w_hn_5_2 = 'b111110000;
logic signed [WIDTH-1:0] w_hn_5_3 = 'b000001110;
logic signed [WIDTH-1:0] w_hn_5_4 = 'b000001100;
logic signed [WIDTH-1:0] w_hn_5_5 = 'b000000100;
logic signed [WIDTH-1:0] w_hn_5_6 = 'b111110111;
logic signed [WIDTH-1:0] w_hn_5_7 = 'b000010101;
logic signed [WIDTH-1:0] w_hn_6_0 = 'b111111111;
logic signed [WIDTH-1:0] w_hn_6_1 = 'b111111110;
logic signed [WIDTH-1:0] w_hn_6_2 = 'b000000101;
logic signed [WIDTH-1:0] w_hn_6_3 = 'b111111010;
logic signed [WIDTH-1:0] w_hn_6_4 = 'b111111010;
logic signed [WIDTH-1:0] w_hn_6_5 = 'b111111111;
logic signed [WIDTH-1:0] w_hn_6_6 = 'b000010111;
logic signed [WIDTH-1:0] w_hn_6_7 = 'b111110100;
logic signed [WIDTH-1:0] w_hn_7_0 = 'b111111111;
logic signed [WIDTH-1:0] w_hn_7_1 = 'b000001110;
logic signed [WIDTH-1:0] w_hn_7_2 = 'b000010100;
logic signed [WIDTH-1:0] w_hn_7_3 = 'b111110010;
logic signed [WIDTH-1:0] w_hn_7_4 = 'b111111011;
logic signed [WIDTH-1:0] w_hn_7_5 = 'b111110110;
logic signed [WIDTH-1:0] w_hn_7_6 = 'b111111001;
logic signed [WIDTH-1:0] w_hn_7_7 = 'b000001010;

// Biases (h for each gate type)
logic signed [WIDTH-1:0] b_ir_0 = 'b000000001;
logic signed [WIDTH-1:0] b_ir_1 = 'b000001000;
logic signed [WIDTH-1:0] b_ir_2 = 'b000001111;
logic signed [WIDTH-1:0] b_ir_3 = 'b000000101;
logic signed [WIDTH-1:0] b_ir_4 = 'b000000110;
logic signed [WIDTH-1:0] b_ir_5 = 'b000000100;
logic signed [WIDTH-1:0] b_ir_6 = 'b000010000;
logic signed [WIDTH-1:0] b_ir_7 = 'b000000000;

logic signed [WIDTH-1:0] b_iz_0 = 'b000001011;
logic signed [WIDTH-1:0] b_iz_1 = 'b000000010;
logic signed [WIDTH-1:0] b_iz_2 = 'b000001110;
logic signed [WIDTH-1:0] b_iz_3 = 'b000000010;
logic signed [WIDTH-1:0] b_iz_4 = 'b000000010;
logic signed [WIDTH-1:0] b_iz_5 = 'b000001010;
logic signed [WIDTH-1:0] b_iz_6 = 'b000000111;
logic signed [WIDTH-1:0] b_iz_7 = 'b000001101;

logic signed [WIDTH-1:0] b_in_0 = 'b000000111;
logic signed [WIDTH-1:0] b_in_1 = 'b000001001;
logic signed [WIDTH-1:0] b_in_2 = 'b000000101;
logic signed [WIDTH-1:0] b_in_3 = 'b000011010;
logic signed [WIDTH-1:0] b_in_4 = 'b000000011;
logic signed [WIDTH-1:0] b_in_5 = 'b000010011;
logic signed [WIDTH-1:0] b_in_6 = 'b000000111;
logic signed [WIDTH-1:0] b_in_7 = 'b111110001;

logic signed [WIDTH-1:0] b_hr_0 = 'b000000001;
logic signed [WIDTH-1:0] b_hr_1 = 'b000001000;
logic signed [WIDTH-1:0] b_hr_2 = 'b000001111;
logic signed [WIDTH-1:0] b_hr_3 = 'b000000101;
logic signed [WIDTH-1:0] b_hr_4 = 'b000000110;
logic signed [WIDTH-1:0] b_hr_5 = 'b000000100;
logic signed [WIDTH-1:0] b_hr_6 = 'b000010000;
logic signed [WIDTH-1:0] b_hr_7 = 'b000000000;

logic signed [WIDTH-1:0] b_hz_0 = 'b000001011;
logic signed [WIDTH-1:0] b_hz_1 = 'b000000010;
logic signed [WIDTH-1:0] b_hz_2 = 'b000001110;
logic signed [WIDTH-1:0] b_hz_3 = 'b000000010;
logic signed [WIDTH-1:0] b_hz_4 = 'b000000010;
logic signed [WIDTH-1:0] b_hz_5 = 'b000001010;
logic signed [WIDTH-1:0] b_hz_6 = 'b000000111;
logic signed [WIDTH-1:0] b_hz_7 = 'b000001101;

logic signed [WIDTH-1:0] b_hn_0 = 'b000000111;
logic signed [WIDTH-1:0] b_hn_1 = 'b000001001;
logic signed [WIDTH-1:0] b_hn_2 = 'b000000101;
logic signed [WIDTH-1:0] b_hn_3 = 'b000011010;
logic signed [WIDTH-1:0] b_hn_4 = 'b000000011;
logic signed [WIDTH-1:0] b_hn_5 = 'b000010011;
logic signed [WIDTH-1:0] b_hn_6 = 'b000000111;
logic signed [WIDTH-1:0] b_hn_7 = 'b111110001;

// Outputs (h=8)
logic signed [WIDTH-1:0]  y_0 = 0;
logic signed [WIDTH-1:0]  y_1 = 0;
logic signed [WIDTH-1:0]  y_2 = 0;
logic signed [WIDTH-1:0]  y_3 = 0;
logic signed [WIDTH-1:0]  y_4 = 0;
logic signed [WIDTH-1:0]  y_5 = 0;
logic signed [WIDTH-1:0]  y_6 = 0;
logic signed [WIDTH-1:0]  y_7 = 0;

gru #(
        .INT_WIDTH(INT_WIDTH),
        .FRAC_WIDTH(FRAC_WIDTH)
    ) gru_inst (
        .clk(clk),
        .reset(reset),
        // Input features (d=64)
        	
.x_0(x_0), .x_1(x_1), .x_2(x_2), .x_3(x_3), .x_4(x_4), .x_5(x_5), .x_6(x_6), .x_7(x_7), .x_8(x_8), .x_9(x_9), .x_10(x_10), .x_11(x_11), .x_12(x_12), .x_13(x_13), .x_14(x_14), .x_15(x_15), .x_16(x_16), .x_17(x_17), .x_18(x_18), .x_19(x_19), .x_20(x_20), .x_21(x_21), .x_22(x_22), .x_23(x_23), .x_24(x_24), .x_25(x_25), .x_26(x_26), .x_27(x_27), .x_28(x_28), .x_29(x_29), .x_30(x_30), .x_31(x_31), .x_32(x_32), .x_33(x_33), .x_34(x_34), .x_35(x_35), .x_36(x_36), .x_37(x_37), .x_38(x_38), .x_39(x_39), .x_40(x_40), .x_41(x_41), .x_42(x_42), .x_43(x_43), .x_44(x_44), .x_45(x_45), .x_46(x_46), .x_47(x_47), .x_48(x_48), .x_49(x_49), .x_50(x_50), .x_51(x_51), .x_52(x_52), .x_53(x_53), .x_54(x_54), .x_55(x_55), .x_56(x_56), .x_57(x_57), .x_58(x_58), .x_59(x_59), .x_60(x_60), .x_61(x_61), .x_62(x_62), .x_63(x_63), .x_64(x_64), .x_65(x_65), .x_66(x_66), .x_67(x_67), .x_68(x_68), .x_69(x_69), .x_70(x_70), .x_71(x_71), .x_72(x_72), .x_73(x_73), .x_74(x_74), .x_75(x_75), .x_76(x_76), .x_77(x_77), .x_78(x_78), .x_79(x_79), .x_80(x_80), .x_81(x_81), .x_82(x_82), .x_83(x_83), .x_84(x_84), .x_85(x_85), .x_86(x_86), .x_87(x_87), .x_88(x_88), .x_89(x_89), .x_90(x_90), .x_91(x_91), .x_92(x_92), .x_93(x_93), .x_94(x_94), .x_95(x_95), .x_96(x_96), .x_97(x_97), .x_98(x_98), .x_99(x_99), .x_100(x_100), .x_101(x_101), .x_102(x_102), .x_103(x_103), .x_104(x_104), .x_105(x_105), .x_106(x_106), .x_107(x_107), .x_108(x_108), .x_109(x_109), .x_110(x_110), .x_111(x_111), .x_112(x_112), .x_113(x_113), .x_114(x_114), .x_115(x_115), .x_116(x_116), .x_117(x_117), .x_118(x_118), .x_119(x_119), .x_120(x_120), .x_121(x_121), .x_122(x_122), .x_123(x_123), .x_124(x_124), .x_125(x_125), .x_126(x_126), .x_127(x_127), .x_128(x_128), .x_129(x_129), .x_130(x_130), .x_131(x_131), .x_132(x_132), .x_133(x_133), .x_134(x_134), .x_135(x_135), .x_136(x_136), .x_137(x_137), .x_138(x_138), .x_139(x_139), .x_140(x_140), .x_141(x_141), .x_142(x_142), .x_143(x_143), .x_144(x_144), .x_145(x_145), .x_146(x_146), .x_147(x_147), .x_148(x_148), .x_149(x_149), .x_150(x_150), .x_151(x_151), .x_152(x_152), .x_153(x_153), .x_154(x_154), .x_155(x_155), .x_156(x_156), .x_157(x_157), .x_158(x_158), .x_159(x_159), .x_160(x_160), .x_161(x_161), .x_162(x_162), .x_163(x_163), .x_164(x_164), .x_165(x_165), .x_166(x_166), .x_167(x_167), .x_168(x_168), .x_169(x_169), .x_170(x_170), .x_171(x_171), .x_172(x_172), .x_173(x_173), .x_174(x_174), .x_175(x_175), .x_176(x_176), .x_177(x_177), .x_178(x_178), .x_179(x_179), .x_180(x_180), .x_181(x_181), .x_182(x_182), .x_183(x_183), .x_184(x_184), .x_185(x_185), .x_186(x_186), .x_187(x_187), .x_188(x_188), .x_189(x_189), .x_190(x_190), .x_191(x_191), .x_192(x_192), .x_193(x_193), .x_194(x_194), .x_195(x_195), .x_196(x_196), .x_197(x_197), .x_198(x_198), .x_199(x_199), .x_200(x_200), .x_201(x_201), .x_202(x_202), .x_203(x_203), .x_204(x_204), .x_205(x_205), .x_206(x_206), .x_207(x_207), .x_208(x_208), .x_209(x_209), .x_210(x_210), .x_211(x_211), .x_212(x_212), .x_213(x_213), .x_214(x_214), .x_215(x_215), .x_216(x_216), .x_217(x_217), .x_218(x_218), .x_219(x_219), .x_220(x_220), .x_221(x_221), .x_222(x_222), .x_223(x_223), .x_224(x_224), .x_225(x_225), .x_226(x_226), .x_227(x_227), .x_228(x_228), .x_229(x_229), .x_230(x_230), .x_231(x_231), .x_232(x_232), .x_233(x_233), .x_234(x_234), .x_235(x_235), .x_236(x_236), .x_237(x_237), .x_238(x_238), .x_239(x_239), .x_240(x_240), .x_241(x_241), .x_242(x_242), .x_243(x_243), .x_244(x_244), .x_245(x_245), .x_246(x_246), .x_247(x_247), .x_248(x_248), .x_249(x_249), .x_250(x_250), .x_251(x_251), .x_252(x_252), .x_253(x_253), .x_254(x_254), .x_255(x_255), 	
.h_0(h_0), .h_1(h_1), .h_2(h_2), .h_3(h_3), .h_4(h_4), .h_5(h_5), .h_6(h_6), .h_7(h_7), 	
.w_ir_0_0(w_ir_0_0), .w_ir_0_1(w_ir_0_1), .w_ir_0_2(w_ir_0_2), .w_ir_0_3(w_ir_0_3), .w_ir_0_4(w_ir_0_4), .w_ir_0_5(w_ir_0_5), .w_ir_0_6(w_ir_0_6), .w_ir_0_7(w_ir_0_7), .w_ir_0_8(w_ir_0_8), .w_ir_0_9(w_ir_0_9), .w_ir_0_10(w_ir_0_10), .w_ir_0_11(w_ir_0_11), .w_ir_0_12(w_ir_0_12), .w_ir_0_13(w_ir_0_13), .w_ir_0_14(w_ir_0_14), .w_ir_0_15(w_ir_0_15), .w_ir_0_16(w_ir_0_16), .w_ir_0_17(w_ir_0_17), .w_ir_0_18(w_ir_0_18), .w_ir_0_19(w_ir_0_19), .w_ir_0_20(w_ir_0_20), .w_ir_0_21(w_ir_0_21), .w_ir_0_22(w_ir_0_22), .w_ir_0_23(w_ir_0_23), .w_ir_0_24(w_ir_0_24), .w_ir_0_25(w_ir_0_25), .w_ir_0_26(w_ir_0_26), .w_ir_0_27(w_ir_0_27), .w_ir_0_28(w_ir_0_28), .w_ir_0_29(w_ir_0_29), .w_ir_0_30(w_ir_0_30), .w_ir_0_31(w_ir_0_31), .w_ir_0_32(w_ir_0_32), .w_ir_0_33(w_ir_0_33), .w_ir_0_34(w_ir_0_34), .w_ir_0_35(w_ir_0_35), .w_ir_0_36(w_ir_0_36), .w_ir_0_37(w_ir_0_37), .w_ir_0_38(w_ir_0_38), .w_ir_0_39(w_ir_0_39), .w_ir_0_40(w_ir_0_40), .w_ir_0_41(w_ir_0_41), .w_ir_0_42(w_ir_0_42), .w_ir_0_43(w_ir_0_43), .w_ir_0_44(w_ir_0_44), .w_ir_0_45(w_ir_0_45), .w_ir_0_46(w_ir_0_46), .w_ir_0_47(w_ir_0_47), .w_ir_0_48(w_ir_0_48), .w_ir_0_49(w_ir_0_49), .w_ir_0_50(w_ir_0_50), .w_ir_0_51(w_ir_0_51), .w_ir_0_52(w_ir_0_52), .w_ir_0_53(w_ir_0_53), .w_ir_0_54(w_ir_0_54), .w_ir_0_55(w_ir_0_55), .w_ir_0_56(w_ir_0_56), .w_ir_0_57(w_ir_0_57), .w_ir_0_58(w_ir_0_58), .w_ir_0_59(w_ir_0_59), .w_ir_0_60(w_ir_0_60), .w_ir_0_61(w_ir_0_61), .w_ir_0_62(w_ir_0_62), .w_ir_0_63(w_ir_0_63), .w_ir_0_64(w_ir_0_64), .w_ir_0_65(w_ir_0_65), .w_ir_0_66(w_ir_0_66), .w_ir_0_67(w_ir_0_67), .w_ir_0_68(w_ir_0_68), .w_ir_0_69(w_ir_0_69), .w_ir_0_70(w_ir_0_70), .w_ir_0_71(w_ir_0_71), .w_ir_0_72(w_ir_0_72), .w_ir_0_73(w_ir_0_73), .w_ir_0_74(w_ir_0_74), .w_ir_0_75(w_ir_0_75), .w_ir_0_76(w_ir_0_76), .w_ir_0_77(w_ir_0_77), .w_ir_0_78(w_ir_0_78), .w_ir_0_79(w_ir_0_79), .w_ir_0_80(w_ir_0_80), .w_ir_0_81(w_ir_0_81), .w_ir_0_82(w_ir_0_82), .w_ir_0_83(w_ir_0_83), .w_ir_0_84(w_ir_0_84), .w_ir_0_85(w_ir_0_85), .w_ir_0_86(w_ir_0_86), .w_ir_0_87(w_ir_0_87), .w_ir_0_88(w_ir_0_88), .w_ir_0_89(w_ir_0_89), .w_ir_0_90(w_ir_0_90), .w_ir_0_91(w_ir_0_91), .w_ir_0_92(w_ir_0_92), .w_ir_0_93(w_ir_0_93), .w_ir_0_94(w_ir_0_94), .w_ir_0_95(w_ir_0_95), .w_ir_0_96(w_ir_0_96), .w_ir_0_97(w_ir_0_97), .w_ir_0_98(w_ir_0_98), .w_ir_0_99(w_ir_0_99), .w_ir_0_100(w_ir_0_100), .w_ir_0_101(w_ir_0_101), .w_ir_0_102(w_ir_0_102), .w_ir_0_103(w_ir_0_103), .w_ir_0_104(w_ir_0_104), .w_ir_0_105(w_ir_0_105), .w_ir_0_106(w_ir_0_106), .w_ir_0_107(w_ir_0_107), .w_ir_0_108(w_ir_0_108), .w_ir_0_109(w_ir_0_109), .w_ir_0_110(w_ir_0_110), .w_ir_0_111(w_ir_0_111), .w_ir_0_112(w_ir_0_112), .w_ir_0_113(w_ir_0_113), .w_ir_0_114(w_ir_0_114), .w_ir_0_115(w_ir_0_115), .w_ir_0_116(w_ir_0_116), .w_ir_0_117(w_ir_0_117), .w_ir_0_118(w_ir_0_118), .w_ir_0_119(w_ir_0_119), .w_ir_0_120(w_ir_0_120), .w_ir_0_121(w_ir_0_121), .w_ir_0_122(w_ir_0_122), .w_ir_0_123(w_ir_0_123), .w_ir_0_124(w_ir_0_124), .w_ir_0_125(w_ir_0_125), .w_ir_0_126(w_ir_0_126), .w_ir_0_127(w_ir_0_127), .w_ir_0_128(w_ir_0_128), .w_ir_0_129(w_ir_0_129), .w_ir_0_130(w_ir_0_130), .w_ir_0_131(w_ir_0_131), .w_ir_0_132(w_ir_0_132), .w_ir_0_133(w_ir_0_133), .w_ir_0_134(w_ir_0_134), .w_ir_0_135(w_ir_0_135), .w_ir_0_136(w_ir_0_136), .w_ir_0_137(w_ir_0_137), .w_ir_0_138(w_ir_0_138), .w_ir_0_139(w_ir_0_139), .w_ir_0_140(w_ir_0_140), .w_ir_0_141(w_ir_0_141), .w_ir_0_142(w_ir_0_142), .w_ir_0_143(w_ir_0_143), .w_ir_0_144(w_ir_0_144), .w_ir_0_145(w_ir_0_145), .w_ir_0_146(w_ir_0_146), .w_ir_0_147(w_ir_0_147), .w_ir_0_148(w_ir_0_148), .w_ir_0_149(w_ir_0_149), .w_ir_0_150(w_ir_0_150), .w_ir_0_151(w_ir_0_151), .w_ir_0_152(w_ir_0_152), .w_ir_0_153(w_ir_0_153), .w_ir_0_154(w_ir_0_154), .w_ir_0_155(w_ir_0_155), .w_ir_0_156(w_ir_0_156), .w_ir_0_157(w_ir_0_157), .w_ir_0_158(w_ir_0_158), .w_ir_0_159(w_ir_0_159), .w_ir_0_160(w_ir_0_160), .w_ir_0_161(w_ir_0_161), .w_ir_0_162(w_ir_0_162), .w_ir_0_163(w_ir_0_163), .w_ir_0_164(w_ir_0_164), .w_ir_0_165(w_ir_0_165), .w_ir_0_166(w_ir_0_166), .w_ir_0_167(w_ir_0_167), .w_ir_0_168(w_ir_0_168), .w_ir_0_169(w_ir_0_169), .w_ir_0_170(w_ir_0_170), .w_ir_0_171(w_ir_0_171), .w_ir_0_172(w_ir_0_172), .w_ir_0_173(w_ir_0_173), .w_ir_0_174(w_ir_0_174), .w_ir_0_175(w_ir_0_175), .w_ir_0_176(w_ir_0_176), .w_ir_0_177(w_ir_0_177), .w_ir_0_178(w_ir_0_178), .w_ir_0_179(w_ir_0_179), .w_ir_0_180(w_ir_0_180), .w_ir_0_181(w_ir_0_181), .w_ir_0_182(w_ir_0_182), .w_ir_0_183(w_ir_0_183), .w_ir_0_184(w_ir_0_184), .w_ir_0_185(w_ir_0_185), .w_ir_0_186(w_ir_0_186), .w_ir_0_187(w_ir_0_187), .w_ir_0_188(w_ir_0_188), .w_ir_0_189(w_ir_0_189), .w_ir_0_190(w_ir_0_190), .w_ir_0_191(w_ir_0_191), .w_ir_0_192(w_ir_0_192), .w_ir_0_193(w_ir_0_193), .w_ir_0_194(w_ir_0_194), .w_ir_0_195(w_ir_0_195), .w_ir_0_196(w_ir_0_196), .w_ir_0_197(w_ir_0_197), .w_ir_0_198(w_ir_0_198), .w_ir_0_199(w_ir_0_199), .w_ir_0_200(w_ir_0_200), .w_ir_0_201(w_ir_0_201), .w_ir_0_202(w_ir_0_202), .w_ir_0_203(w_ir_0_203), .w_ir_0_204(w_ir_0_204), .w_ir_0_205(w_ir_0_205), .w_ir_0_206(w_ir_0_206), .w_ir_0_207(w_ir_0_207), .w_ir_0_208(w_ir_0_208), .w_ir_0_209(w_ir_0_209), .w_ir_0_210(w_ir_0_210), .w_ir_0_211(w_ir_0_211), .w_ir_0_212(w_ir_0_212), .w_ir_0_213(w_ir_0_213), .w_ir_0_214(w_ir_0_214), .w_ir_0_215(w_ir_0_215), .w_ir_0_216(w_ir_0_216), .w_ir_0_217(w_ir_0_217), .w_ir_0_218(w_ir_0_218), .w_ir_0_219(w_ir_0_219), .w_ir_0_220(w_ir_0_220), .w_ir_0_221(w_ir_0_221), .w_ir_0_222(w_ir_0_222), .w_ir_0_223(w_ir_0_223), .w_ir_0_224(w_ir_0_224), .w_ir_0_225(w_ir_0_225), .w_ir_0_226(w_ir_0_226), .w_ir_0_227(w_ir_0_227), .w_ir_0_228(w_ir_0_228), .w_ir_0_229(w_ir_0_229), .w_ir_0_230(w_ir_0_230), .w_ir_0_231(w_ir_0_231), .w_ir_0_232(w_ir_0_232), .w_ir_0_233(w_ir_0_233), .w_ir_0_234(w_ir_0_234), .w_ir_0_235(w_ir_0_235), .w_ir_0_236(w_ir_0_236), .w_ir_0_237(w_ir_0_237), .w_ir_0_238(w_ir_0_238), .w_ir_0_239(w_ir_0_239), .w_ir_0_240(w_ir_0_240), .w_ir_0_241(w_ir_0_241), .w_ir_0_242(w_ir_0_242), .w_ir_0_243(w_ir_0_243), .w_ir_0_244(w_ir_0_244), .w_ir_0_245(w_ir_0_245), .w_ir_0_246(w_ir_0_246), .w_ir_0_247(w_ir_0_247), .w_ir_0_248(w_ir_0_248), .w_ir_0_249(w_ir_0_249), .w_ir_0_250(w_ir_0_250), .w_ir_0_251(w_ir_0_251), .w_ir_0_252(w_ir_0_252), .w_ir_0_253(w_ir_0_253), .w_ir_0_254(w_ir_0_254), .w_ir_0_255(w_ir_0_255), .w_ir_1_0(w_ir_1_0), .w_ir_1_1(w_ir_1_1), .w_ir_1_2(w_ir_1_2), .w_ir_1_3(w_ir_1_3), .w_ir_1_4(w_ir_1_4), .w_ir_1_5(w_ir_1_5), .w_ir_1_6(w_ir_1_6), .w_ir_1_7(w_ir_1_7), .w_ir_1_8(w_ir_1_8), .w_ir_1_9(w_ir_1_9), .w_ir_1_10(w_ir_1_10), .w_ir_1_11(w_ir_1_11), .w_ir_1_12(w_ir_1_12), .w_ir_1_13(w_ir_1_13), .w_ir_1_14(w_ir_1_14), .w_ir_1_15(w_ir_1_15), .w_ir_1_16(w_ir_1_16), .w_ir_1_17(w_ir_1_17), .w_ir_1_18(w_ir_1_18), .w_ir_1_19(w_ir_1_19), .w_ir_1_20(w_ir_1_20), .w_ir_1_21(w_ir_1_21), .w_ir_1_22(w_ir_1_22), .w_ir_1_23(w_ir_1_23), .w_ir_1_24(w_ir_1_24), .w_ir_1_25(w_ir_1_25), .w_ir_1_26(w_ir_1_26), .w_ir_1_27(w_ir_1_27), .w_ir_1_28(w_ir_1_28), .w_ir_1_29(w_ir_1_29), .w_ir_1_30(w_ir_1_30), .w_ir_1_31(w_ir_1_31), .w_ir_1_32(w_ir_1_32), .w_ir_1_33(w_ir_1_33), .w_ir_1_34(w_ir_1_34), .w_ir_1_35(w_ir_1_35), .w_ir_1_36(w_ir_1_36), .w_ir_1_37(w_ir_1_37), .w_ir_1_38(w_ir_1_38), .w_ir_1_39(w_ir_1_39), .w_ir_1_40(w_ir_1_40), .w_ir_1_41(w_ir_1_41), .w_ir_1_42(w_ir_1_42), .w_ir_1_43(w_ir_1_43), .w_ir_1_44(w_ir_1_44), .w_ir_1_45(w_ir_1_45), .w_ir_1_46(w_ir_1_46), .w_ir_1_47(w_ir_1_47), .w_ir_1_48(w_ir_1_48), .w_ir_1_49(w_ir_1_49), .w_ir_1_50(w_ir_1_50), .w_ir_1_51(w_ir_1_51), .w_ir_1_52(w_ir_1_52), .w_ir_1_53(w_ir_1_53), .w_ir_1_54(w_ir_1_54), .w_ir_1_55(w_ir_1_55), .w_ir_1_56(w_ir_1_56), .w_ir_1_57(w_ir_1_57), .w_ir_1_58(w_ir_1_58), .w_ir_1_59(w_ir_1_59), .w_ir_1_60(w_ir_1_60), .w_ir_1_61(w_ir_1_61), .w_ir_1_62(w_ir_1_62), .w_ir_1_63(w_ir_1_63), .w_ir_1_64(w_ir_1_64), .w_ir_1_65(w_ir_1_65), .w_ir_1_66(w_ir_1_66), .w_ir_1_67(w_ir_1_67), .w_ir_1_68(w_ir_1_68), .w_ir_1_69(w_ir_1_69), .w_ir_1_70(w_ir_1_70), .w_ir_1_71(w_ir_1_71), .w_ir_1_72(w_ir_1_72), .w_ir_1_73(w_ir_1_73), .w_ir_1_74(w_ir_1_74), .w_ir_1_75(w_ir_1_75), .w_ir_1_76(w_ir_1_76), .w_ir_1_77(w_ir_1_77), .w_ir_1_78(w_ir_1_78), .w_ir_1_79(w_ir_1_79), .w_ir_1_80(w_ir_1_80), .w_ir_1_81(w_ir_1_81), .w_ir_1_82(w_ir_1_82), .w_ir_1_83(w_ir_1_83), .w_ir_1_84(w_ir_1_84), .w_ir_1_85(w_ir_1_85), .w_ir_1_86(w_ir_1_86), .w_ir_1_87(w_ir_1_87), .w_ir_1_88(w_ir_1_88), .w_ir_1_89(w_ir_1_89), .w_ir_1_90(w_ir_1_90), .w_ir_1_91(w_ir_1_91), .w_ir_1_92(w_ir_1_92), .w_ir_1_93(w_ir_1_93), .w_ir_1_94(w_ir_1_94), .w_ir_1_95(w_ir_1_95), .w_ir_1_96(w_ir_1_96), .w_ir_1_97(w_ir_1_97), .w_ir_1_98(w_ir_1_98), .w_ir_1_99(w_ir_1_99), .w_ir_1_100(w_ir_1_100), .w_ir_1_101(w_ir_1_101), .w_ir_1_102(w_ir_1_102), .w_ir_1_103(w_ir_1_103), .w_ir_1_104(w_ir_1_104), .w_ir_1_105(w_ir_1_105), .w_ir_1_106(w_ir_1_106), .w_ir_1_107(w_ir_1_107), .w_ir_1_108(w_ir_1_108), .w_ir_1_109(w_ir_1_109), .w_ir_1_110(w_ir_1_110), .w_ir_1_111(w_ir_1_111), .w_ir_1_112(w_ir_1_112), .w_ir_1_113(w_ir_1_113), .w_ir_1_114(w_ir_1_114), .w_ir_1_115(w_ir_1_115), .w_ir_1_116(w_ir_1_116), .w_ir_1_117(w_ir_1_117), .w_ir_1_118(w_ir_1_118), .w_ir_1_119(w_ir_1_119), .w_ir_1_120(w_ir_1_120), .w_ir_1_121(w_ir_1_121), .w_ir_1_122(w_ir_1_122), .w_ir_1_123(w_ir_1_123), .w_ir_1_124(w_ir_1_124), .w_ir_1_125(w_ir_1_125), .w_ir_1_126(w_ir_1_126), .w_ir_1_127(w_ir_1_127), .w_ir_1_128(w_ir_1_128), .w_ir_1_129(w_ir_1_129), .w_ir_1_130(w_ir_1_130), .w_ir_1_131(w_ir_1_131), .w_ir_1_132(w_ir_1_132), .w_ir_1_133(w_ir_1_133), .w_ir_1_134(w_ir_1_134), .w_ir_1_135(w_ir_1_135), .w_ir_1_136(w_ir_1_136), .w_ir_1_137(w_ir_1_137), .w_ir_1_138(w_ir_1_138), .w_ir_1_139(w_ir_1_139), .w_ir_1_140(w_ir_1_140), .w_ir_1_141(w_ir_1_141), .w_ir_1_142(w_ir_1_142), .w_ir_1_143(w_ir_1_143), .w_ir_1_144(w_ir_1_144), .w_ir_1_145(w_ir_1_145), .w_ir_1_146(w_ir_1_146), .w_ir_1_147(w_ir_1_147), .w_ir_1_148(w_ir_1_148), .w_ir_1_149(w_ir_1_149), .w_ir_1_150(w_ir_1_150), .w_ir_1_151(w_ir_1_151), .w_ir_1_152(w_ir_1_152), .w_ir_1_153(w_ir_1_153), .w_ir_1_154(w_ir_1_154), .w_ir_1_155(w_ir_1_155), .w_ir_1_156(w_ir_1_156), .w_ir_1_157(w_ir_1_157), .w_ir_1_158(w_ir_1_158), .w_ir_1_159(w_ir_1_159), .w_ir_1_160(w_ir_1_160), .w_ir_1_161(w_ir_1_161), .w_ir_1_162(w_ir_1_162), .w_ir_1_163(w_ir_1_163), .w_ir_1_164(w_ir_1_164), .w_ir_1_165(w_ir_1_165), .w_ir_1_166(w_ir_1_166), .w_ir_1_167(w_ir_1_167), .w_ir_1_168(w_ir_1_168), .w_ir_1_169(w_ir_1_169), .w_ir_1_170(w_ir_1_170), .w_ir_1_171(w_ir_1_171), .w_ir_1_172(w_ir_1_172), .w_ir_1_173(w_ir_1_173), .w_ir_1_174(w_ir_1_174), .w_ir_1_175(w_ir_1_175), .w_ir_1_176(w_ir_1_176), .w_ir_1_177(w_ir_1_177), .w_ir_1_178(w_ir_1_178), .w_ir_1_179(w_ir_1_179), .w_ir_1_180(w_ir_1_180), .w_ir_1_181(w_ir_1_181), .w_ir_1_182(w_ir_1_182), .w_ir_1_183(w_ir_1_183), .w_ir_1_184(w_ir_1_184), .w_ir_1_185(w_ir_1_185), .w_ir_1_186(w_ir_1_186), .w_ir_1_187(w_ir_1_187), .w_ir_1_188(w_ir_1_188), .w_ir_1_189(w_ir_1_189), .w_ir_1_190(w_ir_1_190), .w_ir_1_191(w_ir_1_191), .w_ir_1_192(w_ir_1_192), .w_ir_1_193(w_ir_1_193), .w_ir_1_194(w_ir_1_194), .w_ir_1_195(w_ir_1_195), .w_ir_1_196(w_ir_1_196), .w_ir_1_197(w_ir_1_197), .w_ir_1_198(w_ir_1_198), .w_ir_1_199(w_ir_1_199), .w_ir_1_200(w_ir_1_200), .w_ir_1_201(w_ir_1_201), .w_ir_1_202(w_ir_1_202), .w_ir_1_203(w_ir_1_203), .w_ir_1_204(w_ir_1_204), .w_ir_1_205(w_ir_1_205), .w_ir_1_206(w_ir_1_206), .w_ir_1_207(w_ir_1_207), .w_ir_1_208(w_ir_1_208), .w_ir_1_209(w_ir_1_209), .w_ir_1_210(w_ir_1_210), .w_ir_1_211(w_ir_1_211), .w_ir_1_212(w_ir_1_212), .w_ir_1_213(w_ir_1_213), .w_ir_1_214(w_ir_1_214), .w_ir_1_215(w_ir_1_215), .w_ir_1_216(w_ir_1_216), .w_ir_1_217(w_ir_1_217), .w_ir_1_218(w_ir_1_218), .w_ir_1_219(w_ir_1_219), .w_ir_1_220(w_ir_1_220), .w_ir_1_221(w_ir_1_221), .w_ir_1_222(w_ir_1_222), .w_ir_1_223(w_ir_1_223), .w_ir_1_224(w_ir_1_224), .w_ir_1_225(w_ir_1_225), .w_ir_1_226(w_ir_1_226), .w_ir_1_227(w_ir_1_227), .w_ir_1_228(w_ir_1_228), .w_ir_1_229(w_ir_1_229), .w_ir_1_230(w_ir_1_230), .w_ir_1_231(w_ir_1_231), .w_ir_1_232(w_ir_1_232), .w_ir_1_233(w_ir_1_233), .w_ir_1_234(w_ir_1_234), .w_ir_1_235(w_ir_1_235), .w_ir_1_236(w_ir_1_236), .w_ir_1_237(w_ir_1_237), .w_ir_1_238(w_ir_1_238), .w_ir_1_239(w_ir_1_239), .w_ir_1_240(w_ir_1_240), .w_ir_1_241(w_ir_1_241), .w_ir_1_242(w_ir_1_242), .w_ir_1_243(w_ir_1_243), .w_ir_1_244(w_ir_1_244), .w_ir_1_245(w_ir_1_245), .w_ir_1_246(w_ir_1_246), .w_ir_1_247(w_ir_1_247), .w_ir_1_248(w_ir_1_248), .w_ir_1_249(w_ir_1_249), .w_ir_1_250(w_ir_1_250), .w_ir_1_251(w_ir_1_251), .w_ir_1_252(w_ir_1_252), .w_ir_1_253(w_ir_1_253), .w_ir_1_254(w_ir_1_254), .w_ir_1_255(w_ir_1_255), .w_ir_2_0(w_ir_2_0), .w_ir_2_1(w_ir_2_1), .w_ir_2_2(w_ir_2_2), .w_ir_2_3(w_ir_2_3), .w_ir_2_4(w_ir_2_4), .w_ir_2_5(w_ir_2_5), .w_ir_2_6(w_ir_2_6), .w_ir_2_7(w_ir_2_7), .w_ir_2_8(w_ir_2_8), .w_ir_2_9(w_ir_2_9), .w_ir_2_10(w_ir_2_10), .w_ir_2_11(w_ir_2_11), .w_ir_2_12(w_ir_2_12), .w_ir_2_13(w_ir_2_13), .w_ir_2_14(w_ir_2_14), .w_ir_2_15(w_ir_2_15), .w_ir_2_16(w_ir_2_16), .w_ir_2_17(w_ir_2_17), .w_ir_2_18(w_ir_2_18), .w_ir_2_19(w_ir_2_19), .w_ir_2_20(w_ir_2_20), .w_ir_2_21(w_ir_2_21), .w_ir_2_22(w_ir_2_22), .w_ir_2_23(w_ir_2_23), .w_ir_2_24(w_ir_2_24), .w_ir_2_25(w_ir_2_25), .w_ir_2_26(w_ir_2_26), .w_ir_2_27(w_ir_2_27), .w_ir_2_28(w_ir_2_28), .w_ir_2_29(w_ir_2_29), .w_ir_2_30(w_ir_2_30), .w_ir_2_31(w_ir_2_31), .w_ir_2_32(w_ir_2_32), .w_ir_2_33(w_ir_2_33), .w_ir_2_34(w_ir_2_34), .w_ir_2_35(w_ir_2_35), .w_ir_2_36(w_ir_2_36), .w_ir_2_37(w_ir_2_37), .w_ir_2_38(w_ir_2_38), .w_ir_2_39(w_ir_2_39), .w_ir_2_40(w_ir_2_40), .w_ir_2_41(w_ir_2_41), .w_ir_2_42(w_ir_2_42), .w_ir_2_43(w_ir_2_43), .w_ir_2_44(w_ir_2_44), .w_ir_2_45(w_ir_2_45), .w_ir_2_46(w_ir_2_46), .w_ir_2_47(w_ir_2_47), .w_ir_2_48(w_ir_2_48), .w_ir_2_49(w_ir_2_49), .w_ir_2_50(w_ir_2_50), .w_ir_2_51(w_ir_2_51), .w_ir_2_52(w_ir_2_52), .w_ir_2_53(w_ir_2_53), .w_ir_2_54(w_ir_2_54), .w_ir_2_55(w_ir_2_55), .w_ir_2_56(w_ir_2_56), .w_ir_2_57(w_ir_2_57), .w_ir_2_58(w_ir_2_58), .w_ir_2_59(w_ir_2_59), .w_ir_2_60(w_ir_2_60), .w_ir_2_61(w_ir_2_61), .w_ir_2_62(w_ir_2_62), .w_ir_2_63(w_ir_2_63), .w_ir_2_64(w_ir_2_64), .w_ir_2_65(w_ir_2_65), .w_ir_2_66(w_ir_2_66), .w_ir_2_67(w_ir_2_67), .w_ir_2_68(w_ir_2_68), .w_ir_2_69(w_ir_2_69), .w_ir_2_70(w_ir_2_70), .w_ir_2_71(w_ir_2_71), .w_ir_2_72(w_ir_2_72), .w_ir_2_73(w_ir_2_73), .w_ir_2_74(w_ir_2_74), .w_ir_2_75(w_ir_2_75), .w_ir_2_76(w_ir_2_76), .w_ir_2_77(w_ir_2_77), .w_ir_2_78(w_ir_2_78), .w_ir_2_79(w_ir_2_79), .w_ir_2_80(w_ir_2_80), .w_ir_2_81(w_ir_2_81), .w_ir_2_82(w_ir_2_82), .w_ir_2_83(w_ir_2_83), .w_ir_2_84(w_ir_2_84), .w_ir_2_85(w_ir_2_85), .w_ir_2_86(w_ir_2_86), .w_ir_2_87(w_ir_2_87), .w_ir_2_88(w_ir_2_88), .w_ir_2_89(w_ir_2_89), .w_ir_2_90(w_ir_2_90), .w_ir_2_91(w_ir_2_91), .w_ir_2_92(w_ir_2_92), .w_ir_2_93(w_ir_2_93), .w_ir_2_94(w_ir_2_94), .w_ir_2_95(w_ir_2_95), .w_ir_2_96(w_ir_2_96), .w_ir_2_97(w_ir_2_97), .w_ir_2_98(w_ir_2_98), .w_ir_2_99(w_ir_2_99), .w_ir_2_100(w_ir_2_100), .w_ir_2_101(w_ir_2_101), .w_ir_2_102(w_ir_2_102), .w_ir_2_103(w_ir_2_103), .w_ir_2_104(w_ir_2_104), .w_ir_2_105(w_ir_2_105), .w_ir_2_106(w_ir_2_106), .w_ir_2_107(w_ir_2_107), .w_ir_2_108(w_ir_2_108), .w_ir_2_109(w_ir_2_109), .w_ir_2_110(w_ir_2_110), .w_ir_2_111(w_ir_2_111), .w_ir_2_112(w_ir_2_112), .w_ir_2_113(w_ir_2_113), .w_ir_2_114(w_ir_2_114), .w_ir_2_115(w_ir_2_115), .w_ir_2_116(w_ir_2_116), .w_ir_2_117(w_ir_2_117), .w_ir_2_118(w_ir_2_118), .w_ir_2_119(w_ir_2_119), .w_ir_2_120(w_ir_2_120), .w_ir_2_121(w_ir_2_121), .w_ir_2_122(w_ir_2_122), .w_ir_2_123(w_ir_2_123), .w_ir_2_124(w_ir_2_124), .w_ir_2_125(w_ir_2_125), .w_ir_2_126(w_ir_2_126), .w_ir_2_127(w_ir_2_127), .w_ir_2_128(w_ir_2_128), .w_ir_2_129(w_ir_2_129), .w_ir_2_130(w_ir_2_130), .w_ir_2_131(w_ir_2_131), .w_ir_2_132(w_ir_2_132), .w_ir_2_133(w_ir_2_133), .w_ir_2_134(w_ir_2_134), .w_ir_2_135(w_ir_2_135), .w_ir_2_136(w_ir_2_136), .w_ir_2_137(w_ir_2_137), .w_ir_2_138(w_ir_2_138), .w_ir_2_139(w_ir_2_139), .w_ir_2_140(w_ir_2_140), .w_ir_2_141(w_ir_2_141), .w_ir_2_142(w_ir_2_142), .w_ir_2_143(w_ir_2_143), .w_ir_2_144(w_ir_2_144), .w_ir_2_145(w_ir_2_145), .w_ir_2_146(w_ir_2_146), .w_ir_2_147(w_ir_2_147), .w_ir_2_148(w_ir_2_148), .w_ir_2_149(w_ir_2_149), .w_ir_2_150(w_ir_2_150), .w_ir_2_151(w_ir_2_151), .w_ir_2_152(w_ir_2_152), .w_ir_2_153(w_ir_2_153), .w_ir_2_154(w_ir_2_154), .w_ir_2_155(w_ir_2_155), .w_ir_2_156(w_ir_2_156), .w_ir_2_157(w_ir_2_157), .w_ir_2_158(w_ir_2_158), .w_ir_2_159(w_ir_2_159), .w_ir_2_160(w_ir_2_160), .w_ir_2_161(w_ir_2_161), .w_ir_2_162(w_ir_2_162), .w_ir_2_163(w_ir_2_163), .w_ir_2_164(w_ir_2_164), .w_ir_2_165(w_ir_2_165), .w_ir_2_166(w_ir_2_166), .w_ir_2_167(w_ir_2_167), .w_ir_2_168(w_ir_2_168), .w_ir_2_169(w_ir_2_169), .w_ir_2_170(w_ir_2_170), .w_ir_2_171(w_ir_2_171), .w_ir_2_172(w_ir_2_172), .w_ir_2_173(w_ir_2_173), .w_ir_2_174(w_ir_2_174), .w_ir_2_175(w_ir_2_175), .w_ir_2_176(w_ir_2_176), .w_ir_2_177(w_ir_2_177), .w_ir_2_178(w_ir_2_178), .w_ir_2_179(w_ir_2_179), .w_ir_2_180(w_ir_2_180), .w_ir_2_181(w_ir_2_181), .w_ir_2_182(w_ir_2_182), .w_ir_2_183(w_ir_2_183), .w_ir_2_184(w_ir_2_184), .w_ir_2_185(w_ir_2_185), .w_ir_2_186(w_ir_2_186), .w_ir_2_187(w_ir_2_187), .w_ir_2_188(w_ir_2_188), .w_ir_2_189(w_ir_2_189), .w_ir_2_190(w_ir_2_190), .w_ir_2_191(w_ir_2_191), .w_ir_2_192(w_ir_2_192), .w_ir_2_193(w_ir_2_193), .w_ir_2_194(w_ir_2_194), .w_ir_2_195(w_ir_2_195), .w_ir_2_196(w_ir_2_196), .w_ir_2_197(w_ir_2_197), .w_ir_2_198(w_ir_2_198), .w_ir_2_199(w_ir_2_199), .w_ir_2_200(w_ir_2_200), .w_ir_2_201(w_ir_2_201), .w_ir_2_202(w_ir_2_202), .w_ir_2_203(w_ir_2_203), .w_ir_2_204(w_ir_2_204), .w_ir_2_205(w_ir_2_205), .w_ir_2_206(w_ir_2_206), .w_ir_2_207(w_ir_2_207), .w_ir_2_208(w_ir_2_208), .w_ir_2_209(w_ir_2_209), .w_ir_2_210(w_ir_2_210), .w_ir_2_211(w_ir_2_211), .w_ir_2_212(w_ir_2_212), .w_ir_2_213(w_ir_2_213), .w_ir_2_214(w_ir_2_214), .w_ir_2_215(w_ir_2_215), .w_ir_2_216(w_ir_2_216), .w_ir_2_217(w_ir_2_217), .w_ir_2_218(w_ir_2_218), .w_ir_2_219(w_ir_2_219), .w_ir_2_220(w_ir_2_220), .w_ir_2_221(w_ir_2_221), .w_ir_2_222(w_ir_2_222), .w_ir_2_223(w_ir_2_223), .w_ir_2_224(w_ir_2_224), .w_ir_2_225(w_ir_2_225), .w_ir_2_226(w_ir_2_226), .w_ir_2_227(w_ir_2_227), .w_ir_2_228(w_ir_2_228), .w_ir_2_229(w_ir_2_229), .w_ir_2_230(w_ir_2_230), .w_ir_2_231(w_ir_2_231), .w_ir_2_232(w_ir_2_232), .w_ir_2_233(w_ir_2_233), .w_ir_2_234(w_ir_2_234), .w_ir_2_235(w_ir_2_235), .w_ir_2_236(w_ir_2_236), .w_ir_2_237(w_ir_2_237), .w_ir_2_238(w_ir_2_238), .w_ir_2_239(w_ir_2_239), .w_ir_2_240(w_ir_2_240), .w_ir_2_241(w_ir_2_241), .w_ir_2_242(w_ir_2_242), .w_ir_2_243(w_ir_2_243), .w_ir_2_244(w_ir_2_244), .w_ir_2_245(w_ir_2_245), .w_ir_2_246(w_ir_2_246), .w_ir_2_247(w_ir_2_247), .w_ir_2_248(w_ir_2_248), .w_ir_2_249(w_ir_2_249), .w_ir_2_250(w_ir_2_250), .w_ir_2_251(w_ir_2_251), .w_ir_2_252(w_ir_2_252), .w_ir_2_253(w_ir_2_253), .w_ir_2_254(w_ir_2_254), .w_ir_2_255(w_ir_2_255), .w_ir_3_0(w_ir_3_0), .w_ir_3_1(w_ir_3_1), .w_ir_3_2(w_ir_3_2), .w_ir_3_3(w_ir_3_3), .w_ir_3_4(w_ir_3_4), .w_ir_3_5(w_ir_3_5), .w_ir_3_6(w_ir_3_6), .w_ir_3_7(w_ir_3_7), .w_ir_3_8(w_ir_3_8), .w_ir_3_9(w_ir_3_9), .w_ir_3_10(w_ir_3_10), .w_ir_3_11(w_ir_3_11), .w_ir_3_12(w_ir_3_12), .w_ir_3_13(w_ir_3_13), .w_ir_3_14(w_ir_3_14), .w_ir_3_15(w_ir_3_15), .w_ir_3_16(w_ir_3_16), .w_ir_3_17(w_ir_3_17), .w_ir_3_18(w_ir_3_18), .w_ir_3_19(w_ir_3_19), .w_ir_3_20(w_ir_3_20), .w_ir_3_21(w_ir_3_21), .w_ir_3_22(w_ir_3_22), .w_ir_3_23(w_ir_3_23), .w_ir_3_24(w_ir_3_24), .w_ir_3_25(w_ir_3_25), .w_ir_3_26(w_ir_3_26), .w_ir_3_27(w_ir_3_27), .w_ir_3_28(w_ir_3_28), .w_ir_3_29(w_ir_3_29), .w_ir_3_30(w_ir_3_30), .w_ir_3_31(w_ir_3_31), .w_ir_3_32(w_ir_3_32), .w_ir_3_33(w_ir_3_33), .w_ir_3_34(w_ir_3_34), .w_ir_3_35(w_ir_3_35), .w_ir_3_36(w_ir_3_36), .w_ir_3_37(w_ir_3_37), .w_ir_3_38(w_ir_3_38), .w_ir_3_39(w_ir_3_39), .w_ir_3_40(w_ir_3_40), .w_ir_3_41(w_ir_3_41), .w_ir_3_42(w_ir_3_42), .w_ir_3_43(w_ir_3_43), .w_ir_3_44(w_ir_3_44), .w_ir_3_45(w_ir_3_45), .w_ir_3_46(w_ir_3_46), .w_ir_3_47(w_ir_3_47), .w_ir_3_48(w_ir_3_48), .w_ir_3_49(w_ir_3_49), .w_ir_3_50(w_ir_3_50), .w_ir_3_51(w_ir_3_51), .w_ir_3_52(w_ir_3_52), .w_ir_3_53(w_ir_3_53), .w_ir_3_54(w_ir_3_54), .w_ir_3_55(w_ir_3_55), .w_ir_3_56(w_ir_3_56), .w_ir_3_57(w_ir_3_57), .w_ir_3_58(w_ir_3_58), .w_ir_3_59(w_ir_3_59), .w_ir_3_60(w_ir_3_60), .w_ir_3_61(w_ir_3_61), .w_ir_3_62(w_ir_3_62), .w_ir_3_63(w_ir_3_63), .w_ir_3_64(w_ir_3_64), .w_ir_3_65(w_ir_3_65), .w_ir_3_66(w_ir_3_66), .w_ir_3_67(w_ir_3_67), .w_ir_3_68(w_ir_3_68), .w_ir_3_69(w_ir_3_69), .w_ir_3_70(w_ir_3_70), .w_ir_3_71(w_ir_3_71), .w_ir_3_72(w_ir_3_72), .w_ir_3_73(w_ir_3_73), .w_ir_3_74(w_ir_3_74), .w_ir_3_75(w_ir_3_75), .w_ir_3_76(w_ir_3_76), .w_ir_3_77(w_ir_3_77), .w_ir_3_78(w_ir_3_78), .w_ir_3_79(w_ir_3_79), .w_ir_3_80(w_ir_3_80), .w_ir_3_81(w_ir_3_81), .w_ir_3_82(w_ir_3_82), .w_ir_3_83(w_ir_3_83), .w_ir_3_84(w_ir_3_84), .w_ir_3_85(w_ir_3_85), .w_ir_3_86(w_ir_3_86), .w_ir_3_87(w_ir_3_87), .w_ir_3_88(w_ir_3_88), .w_ir_3_89(w_ir_3_89), .w_ir_3_90(w_ir_3_90), .w_ir_3_91(w_ir_3_91), .w_ir_3_92(w_ir_3_92), .w_ir_3_93(w_ir_3_93), .w_ir_3_94(w_ir_3_94), .w_ir_3_95(w_ir_3_95), .w_ir_3_96(w_ir_3_96), .w_ir_3_97(w_ir_3_97), .w_ir_3_98(w_ir_3_98), .w_ir_3_99(w_ir_3_99), .w_ir_3_100(w_ir_3_100), .w_ir_3_101(w_ir_3_101), .w_ir_3_102(w_ir_3_102), .w_ir_3_103(w_ir_3_103), .w_ir_3_104(w_ir_3_104), .w_ir_3_105(w_ir_3_105), .w_ir_3_106(w_ir_3_106), .w_ir_3_107(w_ir_3_107), .w_ir_3_108(w_ir_3_108), .w_ir_3_109(w_ir_3_109), .w_ir_3_110(w_ir_3_110), .w_ir_3_111(w_ir_3_111), .w_ir_3_112(w_ir_3_112), .w_ir_3_113(w_ir_3_113), .w_ir_3_114(w_ir_3_114), .w_ir_3_115(w_ir_3_115), .w_ir_3_116(w_ir_3_116), .w_ir_3_117(w_ir_3_117), .w_ir_3_118(w_ir_3_118), .w_ir_3_119(w_ir_3_119), .w_ir_3_120(w_ir_3_120), .w_ir_3_121(w_ir_3_121), .w_ir_3_122(w_ir_3_122), .w_ir_3_123(w_ir_3_123), .w_ir_3_124(w_ir_3_124), .w_ir_3_125(w_ir_3_125), .w_ir_3_126(w_ir_3_126), .w_ir_3_127(w_ir_3_127), .w_ir_3_128(w_ir_3_128), .w_ir_3_129(w_ir_3_129), .w_ir_3_130(w_ir_3_130), .w_ir_3_131(w_ir_3_131), .w_ir_3_132(w_ir_3_132), .w_ir_3_133(w_ir_3_133), .w_ir_3_134(w_ir_3_134), .w_ir_3_135(w_ir_3_135), .w_ir_3_136(w_ir_3_136), .w_ir_3_137(w_ir_3_137), .w_ir_3_138(w_ir_3_138), .w_ir_3_139(w_ir_3_139), .w_ir_3_140(w_ir_3_140), .w_ir_3_141(w_ir_3_141), .w_ir_3_142(w_ir_3_142), .w_ir_3_143(w_ir_3_143), .w_ir_3_144(w_ir_3_144), .w_ir_3_145(w_ir_3_145), .w_ir_3_146(w_ir_3_146), .w_ir_3_147(w_ir_3_147), .w_ir_3_148(w_ir_3_148), .w_ir_3_149(w_ir_3_149), .w_ir_3_150(w_ir_3_150), .w_ir_3_151(w_ir_3_151), .w_ir_3_152(w_ir_3_152), .w_ir_3_153(w_ir_3_153), .w_ir_3_154(w_ir_3_154), .w_ir_3_155(w_ir_3_155), .w_ir_3_156(w_ir_3_156), .w_ir_3_157(w_ir_3_157), .w_ir_3_158(w_ir_3_158), .w_ir_3_159(w_ir_3_159), .w_ir_3_160(w_ir_3_160), .w_ir_3_161(w_ir_3_161), .w_ir_3_162(w_ir_3_162), .w_ir_3_163(w_ir_3_163), .w_ir_3_164(w_ir_3_164), .w_ir_3_165(w_ir_3_165), .w_ir_3_166(w_ir_3_166), .w_ir_3_167(w_ir_3_167), .w_ir_3_168(w_ir_3_168), .w_ir_3_169(w_ir_3_169), .w_ir_3_170(w_ir_3_170), .w_ir_3_171(w_ir_3_171), .w_ir_3_172(w_ir_3_172), .w_ir_3_173(w_ir_3_173), .w_ir_3_174(w_ir_3_174), .w_ir_3_175(w_ir_3_175), .w_ir_3_176(w_ir_3_176), .w_ir_3_177(w_ir_3_177), .w_ir_3_178(w_ir_3_178), .w_ir_3_179(w_ir_3_179), .w_ir_3_180(w_ir_3_180), .w_ir_3_181(w_ir_3_181), .w_ir_3_182(w_ir_3_182), .w_ir_3_183(w_ir_3_183), .w_ir_3_184(w_ir_3_184), .w_ir_3_185(w_ir_3_185), .w_ir_3_186(w_ir_3_186), .w_ir_3_187(w_ir_3_187), .w_ir_3_188(w_ir_3_188), .w_ir_3_189(w_ir_3_189), .w_ir_3_190(w_ir_3_190), .w_ir_3_191(w_ir_3_191), .w_ir_3_192(w_ir_3_192), .w_ir_3_193(w_ir_3_193), .w_ir_3_194(w_ir_3_194), .w_ir_3_195(w_ir_3_195), .w_ir_3_196(w_ir_3_196), .w_ir_3_197(w_ir_3_197), .w_ir_3_198(w_ir_3_198), .w_ir_3_199(w_ir_3_199), .w_ir_3_200(w_ir_3_200), .w_ir_3_201(w_ir_3_201), .w_ir_3_202(w_ir_3_202), .w_ir_3_203(w_ir_3_203), .w_ir_3_204(w_ir_3_204), .w_ir_3_205(w_ir_3_205), .w_ir_3_206(w_ir_3_206), .w_ir_3_207(w_ir_3_207), .w_ir_3_208(w_ir_3_208), .w_ir_3_209(w_ir_3_209), .w_ir_3_210(w_ir_3_210), .w_ir_3_211(w_ir_3_211), .w_ir_3_212(w_ir_3_212), .w_ir_3_213(w_ir_3_213), .w_ir_3_214(w_ir_3_214), .w_ir_3_215(w_ir_3_215), .w_ir_3_216(w_ir_3_216), .w_ir_3_217(w_ir_3_217), .w_ir_3_218(w_ir_3_218), .w_ir_3_219(w_ir_3_219), .w_ir_3_220(w_ir_3_220), .w_ir_3_221(w_ir_3_221), .w_ir_3_222(w_ir_3_222), .w_ir_3_223(w_ir_3_223), .w_ir_3_224(w_ir_3_224), .w_ir_3_225(w_ir_3_225), .w_ir_3_226(w_ir_3_226), .w_ir_3_227(w_ir_3_227), .w_ir_3_228(w_ir_3_228), .w_ir_3_229(w_ir_3_229), .w_ir_3_230(w_ir_3_230), .w_ir_3_231(w_ir_3_231), .w_ir_3_232(w_ir_3_232), .w_ir_3_233(w_ir_3_233), .w_ir_3_234(w_ir_3_234), .w_ir_3_235(w_ir_3_235), .w_ir_3_236(w_ir_3_236), .w_ir_3_237(w_ir_3_237), .w_ir_3_238(w_ir_3_238), .w_ir_3_239(w_ir_3_239), .w_ir_3_240(w_ir_3_240), .w_ir_3_241(w_ir_3_241), .w_ir_3_242(w_ir_3_242), .w_ir_3_243(w_ir_3_243), .w_ir_3_244(w_ir_3_244), .w_ir_3_245(w_ir_3_245), .w_ir_3_246(w_ir_3_246), .w_ir_3_247(w_ir_3_247), .w_ir_3_248(w_ir_3_248), .w_ir_3_249(w_ir_3_249), .w_ir_3_250(w_ir_3_250), .w_ir_3_251(w_ir_3_251), .w_ir_3_252(w_ir_3_252), .w_ir_3_253(w_ir_3_253), .w_ir_3_254(w_ir_3_254), .w_ir_3_255(w_ir_3_255), .w_ir_4_0(w_ir_4_0), .w_ir_4_1(w_ir_4_1), .w_ir_4_2(w_ir_4_2), .w_ir_4_3(w_ir_4_3), .w_ir_4_4(w_ir_4_4), .w_ir_4_5(w_ir_4_5), .w_ir_4_6(w_ir_4_6), .w_ir_4_7(w_ir_4_7), .w_ir_4_8(w_ir_4_8), .w_ir_4_9(w_ir_4_9), .w_ir_4_10(w_ir_4_10), .w_ir_4_11(w_ir_4_11), .w_ir_4_12(w_ir_4_12), .w_ir_4_13(w_ir_4_13), .w_ir_4_14(w_ir_4_14), .w_ir_4_15(w_ir_4_15), .w_ir_4_16(w_ir_4_16), .w_ir_4_17(w_ir_4_17), .w_ir_4_18(w_ir_4_18), .w_ir_4_19(w_ir_4_19), .w_ir_4_20(w_ir_4_20), .w_ir_4_21(w_ir_4_21), .w_ir_4_22(w_ir_4_22), .w_ir_4_23(w_ir_4_23), .w_ir_4_24(w_ir_4_24), .w_ir_4_25(w_ir_4_25), .w_ir_4_26(w_ir_4_26), .w_ir_4_27(w_ir_4_27), .w_ir_4_28(w_ir_4_28), .w_ir_4_29(w_ir_4_29), .w_ir_4_30(w_ir_4_30), .w_ir_4_31(w_ir_4_31), .w_ir_4_32(w_ir_4_32), .w_ir_4_33(w_ir_4_33), .w_ir_4_34(w_ir_4_34), .w_ir_4_35(w_ir_4_35), .w_ir_4_36(w_ir_4_36), .w_ir_4_37(w_ir_4_37), .w_ir_4_38(w_ir_4_38), .w_ir_4_39(w_ir_4_39), .w_ir_4_40(w_ir_4_40), .w_ir_4_41(w_ir_4_41), .w_ir_4_42(w_ir_4_42), .w_ir_4_43(w_ir_4_43), .w_ir_4_44(w_ir_4_44), .w_ir_4_45(w_ir_4_45), .w_ir_4_46(w_ir_4_46), .w_ir_4_47(w_ir_4_47), .w_ir_4_48(w_ir_4_48), .w_ir_4_49(w_ir_4_49), .w_ir_4_50(w_ir_4_50), .w_ir_4_51(w_ir_4_51), .w_ir_4_52(w_ir_4_52), .w_ir_4_53(w_ir_4_53), .w_ir_4_54(w_ir_4_54), .w_ir_4_55(w_ir_4_55), .w_ir_4_56(w_ir_4_56), .w_ir_4_57(w_ir_4_57), .w_ir_4_58(w_ir_4_58), .w_ir_4_59(w_ir_4_59), .w_ir_4_60(w_ir_4_60), .w_ir_4_61(w_ir_4_61), .w_ir_4_62(w_ir_4_62), .w_ir_4_63(w_ir_4_63), .w_ir_4_64(w_ir_4_64), .w_ir_4_65(w_ir_4_65), .w_ir_4_66(w_ir_4_66), .w_ir_4_67(w_ir_4_67), .w_ir_4_68(w_ir_4_68), .w_ir_4_69(w_ir_4_69), .w_ir_4_70(w_ir_4_70), .w_ir_4_71(w_ir_4_71), .w_ir_4_72(w_ir_4_72), .w_ir_4_73(w_ir_4_73), .w_ir_4_74(w_ir_4_74), .w_ir_4_75(w_ir_4_75), .w_ir_4_76(w_ir_4_76), .w_ir_4_77(w_ir_4_77), .w_ir_4_78(w_ir_4_78), .w_ir_4_79(w_ir_4_79), .w_ir_4_80(w_ir_4_80), .w_ir_4_81(w_ir_4_81), .w_ir_4_82(w_ir_4_82), .w_ir_4_83(w_ir_4_83), .w_ir_4_84(w_ir_4_84), .w_ir_4_85(w_ir_4_85), .w_ir_4_86(w_ir_4_86), .w_ir_4_87(w_ir_4_87), .w_ir_4_88(w_ir_4_88), .w_ir_4_89(w_ir_4_89), .w_ir_4_90(w_ir_4_90), .w_ir_4_91(w_ir_4_91), .w_ir_4_92(w_ir_4_92), .w_ir_4_93(w_ir_4_93), .w_ir_4_94(w_ir_4_94), .w_ir_4_95(w_ir_4_95), .w_ir_4_96(w_ir_4_96), .w_ir_4_97(w_ir_4_97), .w_ir_4_98(w_ir_4_98), .w_ir_4_99(w_ir_4_99), .w_ir_4_100(w_ir_4_100), .w_ir_4_101(w_ir_4_101), .w_ir_4_102(w_ir_4_102), .w_ir_4_103(w_ir_4_103), .w_ir_4_104(w_ir_4_104), .w_ir_4_105(w_ir_4_105), .w_ir_4_106(w_ir_4_106), .w_ir_4_107(w_ir_4_107), .w_ir_4_108(w_ir_4_108), .w_ir_4_109(w_ir_4_109), .w_ir_4_110(w_ir_4_110), .w_ir_4_111(w_ir_4_111), .w_ir_4_112(w_ir_4_112), .w_ir_4_113(w_ir_4_113), .w_ir_4_114(w_ir_4_114), .w_ir_4_115(w_ir_4_115), .w_ir_4_116(w_ir_4_116), .w_ir_4_117(w_ir_4_117), .w_ir_4_118(w_ir_4_118), .w_ir_4_119(w_ir_4_119), .w_ir_4_120(w_ir_4_120), .w_ir_4_121(w_ir_4_121), .w_ir_4_122(w_ir_4_122), .w_ir_4_123(w_ir_4_123), .w_ir_4_124(w_ir_4_124), .w_ir_4_125(w_ir_4_125), .w_ir_4_126(w_ir_4_126), .w_ir_4_127(w_ir_4_127), .w_ir_4_128(w_ir_4_128), .w_ir_4_129(w_ir_4_129), .w_ir_4_130(w_ir_4_130), .w_ir_4_131(w_ir_4_131), .w_ir_4_132(w_ir_4_132), .w_ir_4_133(w_ir_4_133), .w_ir_4_134(w_ir_4_134), .w_ir_4_135(w_ir_4_135), .w_ir_4_136(w_ir_4_136), .w_ir_4_137(w_ir_4_137), .w_ir_4_138(w_ir_4_138), .w_ir_4_139(w_ir_4_139), .w_ir_4_140(w_ir_4_140), .w_ir_4_141(w_ir_4_141), .w_ir_4_142(w_ir_4_142), .w_ir_4_143(w_ir_4_143), .w_ir_4_144(w_ir_4_144), .w_ir_4_145(w_ir_4_145), .w_ir_4_146(w_ir_4_146), .w_ir_4_147(w_ir_4_147), .w_ir_4_148(w_ir_4_148), .w_ir_4_149(w_ir_4_149), .w_ir_4_150(w_ir_4_150), .w_ir_4_151(w_ir_4_151), .w_ir_4_152(w_ir_4_152), .w_ir_4_153(w_ir_4_153), .w_ir_4_154(w_ir_4_154), .w_ir_4_155(w_ir_4_155), .w_ir_4_156(w_ir_4_156), .w_ir_4_157(w_ir_4_157), .w_ir_4_158(w_ir_4_158), .w_ir_4_159(w_ir_4_159), .w_ir_4_160(w_ir_4_160), .w_ir_4_161(w_ir_4_161), .w_ir_4_162(w_ir_4_162), .w_ir_4_163(w_ir_4_163), .w_ir_4_164(w_ir_4_164), .w_ir_4_165(w_ir_4_165), .w_ir_4_166(w_ir_4_166), .w_ir_4_167(w_ir_4_167), .w_ir_4_168(w_ir_4_168), .w_ir_4_169(w_ir_4_169), .w_ir_4_170(w_ir_4_170), .w_ir_4_171(w_ir_4_171), .w_ir_4_172(w_ir_4_172), .w_ir_4_173(w_ir_4_173), .w_ir_4_174(w_ir_4_174), .w_ir_4_175(w_ir_4_175), .w_ir_4_176(w_ir_4_176), .w_ir_4_177(w_ir_4_177), .w_ir_4_178(w_ir_4_178), .w_ir_4_179(w_ir_4_179), .w_ir_4_180(w_ir_4_180), .w_ir_4_181(w_ir_4_181), .w_ir_4_182(w_ir_4_182), .w_ir_4_183(w_ir_4_183), .w_ir_4_184(w_ir_4_184), .w_ir_4_185(w_ir_4_185), .w_ir_4_186(w_ir_4_186), .w_ir_4_187(w_ir_4_187), .w_ir_4_188(w_ir_4_188), .w_ir_4_189(w_ir_4_189), .w_ir_4_190(w_ir_4_190), .w_ir_4_191(w_ir_4_191), .w_ir_4_192(w_ir_4_192), .w_ir_4_193(w_ir_4_193), .w_ir_4_194(w_ir_4_194), .w_ir_4_195(w_ir_4_195), .w_ir_4_196(w_ir_4_196), .w_ir_4_197(w_ir_4_197), .w_ir_4_198(w_ir_4_198), .w_ir_4_199(w_ir_4_199), .w_ir_4_200(w_ir_4_200), .w_ir_4_201(w_ir_4_201), .w_ir_4_202(w_ir_4_202), .w_ir_4_203(w_ir_4_203), .w_ir_4_204(w_ir_4_204), .w_ir_4_205(w_ir_4_205), .w_ir_4_206(w_ir_4_206), .w_ir_4_207(w_ir_4_207), .w_ir_4_208(w_ir_4_208), .w_ir_4_209(w_ir_4_209), .w_ir_4_210(w_ir_4_210), .w_ir_4_211(w_ir_4_211), .w_ir_4_212(w_ir_4_212), .w_ir_4_213(w_ir_4_213), .w_ir_4_214(w_ir_4_214), .w_ir_4_215(w_ir_4_215), .w_ir_4_216(w_ir_4_216), .w_ir_4_217(w_ir_4_217), .w_ir_4_218(w_ir_4_218), .w_ir_4_219(w_ir_4_219), .w_ir_4_220(w_ir_4_220), .w_ir_4_221(w_ir_4_221), .w_ir_4_222(w_ir_4_222), .w_ir_4_223(w_ir_4_223), .w_ir_4_224(w_ir_4_224), .w_ir_4_225(w_ir_4_225), .w_ir_4_226(w_ir_4_226), .w_ir_4_227(w_ir_4_227), .w_ir_4_228(w_ir_4_228), .w_ir_4_229(w_ir_4_229), .w_ir_4_230(w_ir_4_230), .w_ir_4_231(w_ir_4_231), .w_ir_4_232(w_ir_4_232), .w_ir_4_233(w_ir_4_233), .w_ir_4_234(w_ir_4_234), .w_ir_4_235(w_ir_4_235), .w_ir_4_236(w_ir_4_236), .w_ir_4_237(w_ir_4_237), .w_ir_4_238(w_ir_4_238), .w_ir_4_239(w_ir_4_239), .w_ir_4_240(w_ir_4_240), .w_ir_4_241(w_ir_4_241), .w_ir_4_242(w_ir_4_242), .w_ir_4_243(w_ir_4_243), .w_ir_4_244(w_ir_4_244), .w_ir_4_245(w_ir_4_245), .w_ir_4_246(w_ir_4_246), .w_ir_4_247(w_ir_4_247), .w_ir_4_248(w_ir_4_248), .w_ir_4_249(w_ir_4_249), .w_ir_4_250(w_ir_4_250), .w_ir_4_251(w_ir_4_251), .w_ir_4_252(w_ir_4_252), .w_ir_4_253(w_ir_4_253), .w_ir_4_254(w_ir_4_254), .w_ir_4_255(w_ir_4_255), .w_ir_5_0(w_ir_5_0), .w_ir_5_1(w_ir_5_1), .w_ir_5_2(w_ir_5_2), .w_ir_5_3(w_ir_5_3), .w_ir_5_4(w_ir_5_4), .w_ir_5_5(w_ir_5_5), .w_ir_5_6(w_ir_5_6), .w_ir_5_7(w_ir_5_7), .w_ir_5_8(w_ir_5_8), .w_ir_5_9(w_ir_5_9), .w_ir_5_10(w_ir_5_10), .w_ir_5_11(w_ir_5_11), .w_ir_5_12(w_ir_5_12), .w_ir_5_13(w_ir_5_13), .w_ir_5_14(w_ir_5_14), .w_ir_5_15(w_ir_5_15), .w_ir_5_16(w_ir_5_16), .w_ir_5_17(w_ir_5_17), .w_ir_5_18(w_ir_5_18), .w_ir_5_19(w_ir_5_19), .w_ir_5_20(w_ir_5_20), .w_ir_5_21(w_ir_5_21), .w_ir_5_22(w_ir_5_22), .w_ir_5_23(w_ir_5_23), .w_ir_5_24(w_ir_5_24), .w_ir_5_25(w_ir_5_25), .w_ir_5_26(w_ir_5_26), .w_ir_5_27(w_ir_5_27), .w_ir_5_28(w_ir_5_28), .w_ir_5_29(w_ir_5_29), .w_ir_5_30(w_ir_5_30), .w_ir_5_31(w_ir_5_31), .w_ir_5_32(w_ir_5_32), .w_ir_5_33(w_ir_5_33), .w_ir_5_34(w_ir_5_34), .w_ir_5_35(w_ir_5_35), .w_ir_5_36(w_ir_5_36), .w_ir_5_37(w_ir_5_37), .w_ir_5_38(w_ir_5_38), .w_ir_5_39(w_ir_5_39), .w_ir_5_40(w_ir_5_40), .w_ir_5_41(w_ir_5_41), .w_ir_5_42(w_ir_5_42), .w_ir_5_43(w_ir_5_43), .w_ir_5_44(w_ir_5_44), .w_ir_5_45(w_ir_5_45), .w_ir_5_46(w_ir_5_46), .w_ir_5_47(w_ir_5_47), .w_ir_5_48(w_ir_5_48), .w_ir_5_49(w_ir_5_49), .w_ir_5_50(w_ir_5_50), .w_ir_5_51(w_ir_5_51), .w_ir_5_52(w_ir_5_52), .w_ir_5_53(w_ir_5_53), .w_ir_5_54(w_ir_5_54), .w_ir_5_55(w_ir_5_55), .w_ir_5_56(w_ir_5_56), .w_ir_5_57(w_ir_5_57), .w_ir_5_58(w_ir_5_58), .w_ir_5_59(w_ir_5_59), .w_ir_5_60(w_ir_5_60), .w_ir_5_61(w_ir_5_61), .w_ir_5_62(w_ir_5_62), .w_ir_5_63(w_ir_5_63), .w_ir_5_64(w_ir_5_64), .w_ir_5_65(w_ir_5_65), .w_ir_5_66(w_ir_5_66), .w_ir_5_67(w_ir_5_67), .w_ir_5_68(w_ir_5_68), .w_ir_5_69(w_ir_5_69), .w_ir_5_70(w_ir_5_70), .w_ir_5_71(w_ir_5_71), .w_ir_5_72(w_ir_5_72), .w_ir_5_73(w_ir_5_73), .w_ir_5_74(w_ir_5_74), .w_ir_5_75(w_ir_5_75), .w_ir_5_76(w_ir_5_76), .w_ir_5_77(w_ir_5_77), .w_ir_5_78(w_ir_5_78), .w_ir_5_79(w_ir_5_79), .w_ir_5_80(w_ir_5_80), .w_ir_5_81(w_ir_5_81), .w_ir_5_82(w_ir_5_82), .w_ir_5_83(w_ir_5_83), .w_ir_5_84(w_ir_5_84), .w_ir_5_85(w_ir_5_85), .w_ir_5_86(w_ir_5_86), .w_ir_5_87(w_ir_5_87), .w_ir_5_88(w_ir_5_88), .w_ir_5_89(w_ir_5_89), .w_ir_5_90(w_ir_5_90), .w_ir_5_91(w_ir_5_91), .w_ir_5_92(w_ir_5_92), .w_ir_5_93(w_ir_5_93), .w_ir_5_94(w_ir_5_94), .w_ir_5_95(w_ir_5_95), .w_ir_5_96(w_ir_5_96), .w_ir_5_97(w_ir_5_97), .w_ir_5_98(w_ir_5_98), .w_ir_5_99(w_ir_5_99), .w_ir_5_100(w_ir_5_100), .w_ir_5_101(w_ir_5_101), .w_ir_5_102(w_ir_5_102), .w_ir_5_103(w_ir_5_103), .w_ir_5_104(w_ir_5_104), .w_ir_5_105(w_ir_5_105), .w_ir_5_106(w_ir_5_106), .w_ir_5_107(w_ir_5_107), .w_ir_5_108(w_ir_5_108), .w_ir_5_109(w_ir_5_109), .w_ir_5_110(w_ir_5_110), .w_ir_5_111(w_ir_5_111), .w_ir_5_112(w_ir_5_112), .w_ir_5_113(w_ir_5_113), .w_ir_5_114(w_ir_5_114), .w_ir_5_115(w_ir_5_115), .w_ir_5_116(w_ir_5_116), .w_ir_5_117(w_ir_5_117), .w_ir_5_118(w_ir_5_118), .w_ir_5_119(w_ir_5_119), .w_ir_5_120(w_ir_5_120), .w_ir_5_121(w_ir_5_121), .w_ir_5_122(w_ir_5_122), .w_ir_5_123(w_ir_5_123), .w_ir_5_124(w_ir_5_124), .w_ir_5_125(w_ir_5_125), .w_ir_5_126(w_ir_5_126), .w_ir_5_127(w_ir_5_127), .w_ir_5_128(w_ir_5_128), .w_ir_5_129(w_ir_5_129), .w_ir_5_130(w_ir_5_130), .w_ir_5_131(w_ir_5_131), .w_ir_5_132(w_ir_5_132), .w_ir_5_133(w_ir_5_133), .w_ir_5_134(w_ir_5_134), .w_ir_5_135(w_ir_5_135), .w_ir_5_136(w_ir_5_136), .w_ir_5_137(w_ir_5_137), .w_ir_5_138(w_ir_5_138), .w_ir_5_139(w_ir_5_139), .w_ir_5_140(w_ir_5_140), .w_ir_5_141(w_ir_5_141), .w_ir_5_142(w_ir_5_142), .w_ir_5_143(w_ir_5_143), .w_ir_5_144(w_ir_5_144), .w_ir_5_145(w_ir_5_145), .w_ir_5_146(w_ir_5_146), .w_ir_5_147(w_ir_5_147), .w_ir_5_148(w_ir_5_148), .w_ir_5_149(w_ir_5_149), .w_ir_5_150(w_ir_5_150), .w_ir_5_151(w_ir_5_151), .w_ir_5_152(w_ir_5_152), .w_ir_5_153(w_ir_5_153), .w_ir_5_154(w_ir_5_154), .w_ir_5_155(w_ir_5_155), .w_ir_5_156(w_ir_5_156), .w_ir_5_157(w_ir_5_157), .w_ir_5_158(w_ir_5_158), .w_ir_5_159(w_ir_5_159), .w_ir_5_160(w_ir_5_160), .w_ir_5_161(w_ir_5_161), .w_ir_5_162(w_ir_5_162), .w_ir_5_163(w_ir_5_163), .w_ir_5_164(w_ir_5_164), .w_ir_5_165(w_ir_5_165), .w_ir_5_166(w_ir_5_166), .w_ir_5_167(w_ir_5_167), .w_ir_5_168(w_ir_5_168), .w_ir_5_169(w_ir_5_169), .w_ir_5_170(w_ir_5_170), .w_ir_5_171(w_ir_5_171), .w_ir_5_172(w_ir_5_172), .w_ir_5_173(w_ir_5_173), .w_ir_5_174(w_ir_5_174), .w_ir_5_175(w_ir_5_175), .w_ir_5_176(w_ir_5_176), .w_ir_5_177(w_ir_5_177), .w_ir_5_178(w_ir_5_178), .w_ir_5_179(w_ir_5_179), .w_ir_5_180(w_ir_5_180), .w_ir_5_181(w_ir_5_181), .w_ir_5_182(w_ir_5_182), .w_ir_5_183(w_ir_5_183), .w_ir_5_184(w_ir_5_184), .w_ir_5_185(w_ir_5_185), .w_ir_5_186(w_ir_5_186), .w_ir_5_187(w_ir_5_187), .w_ir_5_188(w_ir_5_188), .w_ir_5_189(w_ir_5_189), .w_ir_5_190(w_ir_5_190), .w_ir_5_191(w_ir_5_191), .w_ir_5_192(w_ir_5_192), .w_ir_5_193(w_ir_5_193), .w_ir_5_194(w_ir_5_194), .w_ir_5_195(w_ir_5_195), .w_ir_5_196(w_ir_5_196), .w_ir_5_197(w_ir_5_197), .w_ir_5_198(w_ir_5_198), .w_ir_5_199(w_ir_5_199), .w_ir_5_200(w_ir_5_200), .w_ir_5_201(w_ir_5_201), .w_ir_5_202(w_ir_5_202), .w_ir_5_203(w_ir_5_203), .w_ir_5_204(w_ir_5_204), .w_ir_5_205(w_ir_5_205), .w_ir_5_206(w_ir_5_206), .w_ir_5_207(w_ir_5_207), .w_ir_5_208(w_ir_5_208), .w_ir_5_209(w_ir_5_209), .w_ir_5_210(w_ir_5_210), .w_ir_5_211(w_ir_5_211), .w_ir_5_212(w_ir_5_212), .w_ir_5_213(w_ir_5_213), .w_ir_5_214(w_ir_5_214), .w_ir_5_215(w_ir_5_215), .w_ir_5_216(w_ir_5_216), .w_ir_5_217(w_ir_5_217), .w_ir_5_218(w_ir_5_218), .w_ir_5_219(w_ir_5_219), .w_ir_5_220(w_ir_5_220), .w_ir_5_221(w_ir_5_221), .w_ir_5_222(w_ir_5_222), .w_ir_5_223(w_ir_5_223), .w_ir_5_224(w_ir_5_224), .w_ir_5_225(w_ir_5_225), .w_ir_5_226(w_ir_5_226), .w_ir_5_227(w_ir_5_227), .w_ir_5_228(w_ir_5_228), .w_ir_5_229(w_ir_5_229), .w_ir_5_230(w_ir_5_230), .w_ir_5_231(w_ir_5_231), .w_ir_5_232(w_ir_5_232), .w_ir_5_233(w_ir_5_233), .w_ir_5_234(w_ir_5_234), .w_ir_5_235(w_ir_5_235), .w_ir_5_236(w_ir_5_236), .w_ir_5_237(w_ir_5_237), .w_ir_5_238(w_ir_5_238), .w_ir_5_239(w_ir_5_239), .w_ir_5_240(w_ir_5_240), .w_ir_5_241(w_ir_5_241), .w_ir_5_242(w_ir_5_242), .w_ir_5_243(w_ir_5_243), .w_ir_5_244(w_ir_5_244), .w_ir_5_245(w_ir_5_245), .w_ir_5_246(w_ir_5_246), .w_ir_5_247(w_ir_5_247), .w_ir_5_248(w_ir_5_248), .w_ir_5_249(w_ir_5_249), .w_ir_5_250(w_ir_5_250), .w_ir_5_251(w_ir_5_251), .w_ir_5_252(w_ir_5_252), .w_ir_5_253(w_ir_5_253), .w_ir_5_254(w_ir_5_254), .w_ir_5_255(w_ir_5_255), .w_ir_6_0(w_ir_6_0), .w_ir_6_1(w_ir_6_1), .w_ir_6_2(w_ir_6_2), .w_ir_6_3(w_ir_6_3), .w_ir_6_4(w_ir_6_4), .w_ir_6_5(w_ir_6_5), .w_ir_6_6(w_ir_6_6), .w_ir_6_7(w_ir_6_7), .w_ir_6_8(w_ir_6_8), .w_ir_6_9(w_ir_6_9), .w_ir_6_10(w_ir_6_10), .w_ir_6_11(w_ir_6_11), .w_ir_6_12(w_ir_6_12), .w_ir_6_13(w_ir_6_13), .w_ir_6_14(w_ir_6_14), .w_ir_6_15(w_ir_6_15), .w_ir_6_16(w_ir_6_16), .w_ir_6_17(w_ir_6_17), .w_ir_6_18(w_ir_6_18), .w_ir_6_19(w_ir_6_19), .w_ir_6_20(w_ir_6_20), .w_ir_6_21(w_ir_6_21), .w_ir_6_22(w_ir_6_22), .w_ir_6_23(w_ir_6_23), .w_ir_6_24(w_ir_6_24), .w_ir_6_25(w_ir_6_25), .w_ir_6_26(w_ir_6_26), .w_ir_6_27(w_ir_6_27), .w_ir_6_28(w_ir_6_28), .w_ir_6_29(w_ir_6_29), .w_ir_6_30(w_ir_6_30), .w_ir_6_31(w_ir_6_31), .w_ir_6_32(w_ir_6_32), .w_ir_6_33(w_ir_6_33), .w_ir_6_34(w_ir_6_34), .w_ir_6_35(w_ir_6_35), .w_ir_6_36(w_ir_6_36), .w_ir_6_37(w_ir_6_37), .w_ir_6_38(w_ir_6_38), .w_ir_6_39(w_ir_6_39), .w_ir_6_40(w_ir_6_40), .w_ir_6_41(w_ir_6_41), .w_ir_6_42(w_ir_6_42), .w_ir_6_43(w_ir_6_43), .w_ir_6_44(w_ir_6_44), .w_ir_6_45(w_ir_6_45), .w_ir_6_46(w_ir_6_46), .w_ir_6_47(w_ir_6_47), .w_ir_6_48(w_ir_6_48), .w_ir_6_49(w_ir_6_49), .w_ir_6_50(w_ir_6_50), .w_ir_6_51(w_ir_6_51), .w_ir_6_52(w_ir_6_52), .w_ir_6_53(w_ir_6_53), .w_ir_6_54(w_ir_6_54), .w_ir_6_55(w_ir_6_55), .w_ir_6_56(w_ir_6_56), .w_ir_6_57(w_ir_6_57), .w_ir_6_58(w_ir_6_58), .w_ir_6_59(w_ir_6_59), .w_ir_6_60(w_ir_6_60), .w_ir_6_61(w_ir_6_61), .w_ir_6_62(w_ir_6_62), .w_ir_6_63(w_ir_6_63), .w_ir_6_64(w_ir_6_64), .w_ir_6_65(w_ir_6_65), .w_ir_6_66(w_ir_6_66), .w_ir_6_67(w_ir_6_67), .w_ir_6_68(w_ir_6_68), .w_ir_6_69(w_ir_6_69), .w_ir_6_70(w_ir_6_70), .w_ir_6_71(w_ir_6_71), .w_ir_6_72(w_ir_6_72), .w_ir_6_73(w_ir_6_73), .w_ir_6_74(w_ir_6_74), .w_ir_6_75(w_ir_6_75), .w_ir_6_76(w_ir_6_76), .w_ir_6_77(w_ir_6_77), .w_ir_6_78(w_ir_6_78), .w_ir_6_79(w_ir_6_79), .w_ir_6_80(w_ir_6_80), .w_ir_6_81(w_ir_6_81), .w_ir_6_82(w_ir_6_82), .w_ir_6_83(w_ir_6_83), .w_ir_6_84(w_ir_6_84), .w_ir_6_85(w_ir_6_85), .w_ir_6_86(w_ir_6_86), .w_ir_6_87(w_ir_6_87), .w_ir_6_88(w_ir_6_88), .w_ir_6_89(w_ir_6_89), .w_ir_6_90(w_ir_6_90), .w_ir_6_91(w_ir_6_91), .w_ir_6_92(w_ir_6_92), .w_ir_6_93(w_ir_6_93), .w_ir_6_94(w_ir_6_94), .w_ir_6_95(w_ir_6_95), .w_ir_6_96(w_ir_6_96), .w_ir_6_97(w_ir_6_97), .w_ir_6_98(w_ir_6_98), .w_ir_6_99(w_ir_6_99), .w_ir_6_100(w_ir_6_100), .w_ir_6_101(w_ir_6_101), .w_ir_6_102(w_ir_6_102), .w_ir_6_103(w_ir_6_103), .w_ir_6_104(w_ir_6_104), .w_ir_6_105(w_ir_6_105), .w_ir_6_106(w_ir_6_106), .w_ir_6_107(w_ir_6_107), .w_ir_6_108(w_ir_6_108), .w_ir_6_109(w_ir_6_109), .w_ir_6_110(w_ir_6_110), .w_ir_6_111(w_ir_6_111), .w_ir_6_112(w_ir_6_112), .w_ir_6_113(w_ir_6_113), .w_ir_6_114(w_ir_6_114), .w_ir_6_115(w_ir_6_115), .w_ir_6_116(w_ir_6_116), .w_ir_6_117(w_ir_6_117), .w_ir_6_118(w_ir_6_118), .w_ir_6_119(w_ir_6_119), .w_ir_6_120(w_ir_6_120), .w_ir_6_121(w_ir_6_121), .w_ir_6_122(w_ir_6_122), .w_ir_6_123(w_ir_6_123), .w_ir_6_124(w_ir_6_124), .w_ir_6_125(w_ir_6_125), .w_ir_6_126(w_ir_6_126), .w_ir_6_127(w_ir_6_127), .w_ir_6_128(w_ir_6_128), .w_ir_6_129(w_ir_6_129), .w_ir_6_130(w_ir_6_130), .w_ir_6_131(w_ir_6_131), .w_ir_6_132(w_ir_6_132), .w_ir_6_133(w_ir_6_133), .w_ir_6_134(w_ir_6_134), .w_ir_6_135(w_ir_6_135), .w_ir_6_136(w_ir_6_136), .w_ir_6_137(w_ir_6_137), .w_ir_6_138(w_ir_6_138), .w_ir_6_139(w_ir_6_139), .w_ir_6_140(w_ir_6_140), .w_ir_6_141(w_ir_6_141), .w_ir_6_142(w_ir_6_142), .w_ir_6_143(w_ir_6_143), .w_ir_6_144(w_ir_6_144), .w_ir_6_145(w_ir_6_145), .w_ir_6_146(w_ir_6_146), .w_ir_6_147(w_ir_6_147), .w_ir_6_148(w_ir_6_148), .w_ir_6_149(w_ir_6_149), .w_ir_6_150(w_ir_6_150), .w_ir_6_151(w_ir_6_151), .w_ir_6_152(w_ir_6_152), .w_ir_6_153(w_ir_6_153), .w_ir_6_154(w_ir_6_154), .w_ir_6_155(w_ir_6_155), .w_ir_6_156(w_ir_6_156), .w_ir_6_157(w_ir_6_157), .w_ir_6_158(w_ir_6_158), .w_ir_6_159(w_ir_6_159), .w_ir_6_160(w_ir_6_160), .w_ir_6_161(w_ir_6_161), .w_ir_6_162(w_ir_6_162), .w_ir_6_163(w_ir_6_163), .w_ir_6_164(w_ir_6_164), .w_ir_6_165(w_ir_6_165), .w_ir_6_166(w_ir_6_166), .w_ir_6_167(w_ir_6_167), .w_ir_6_168(w_ir_6_168), .w_ir_6_169(w_ir_6_169), .w_ir_6_170(w_ir_6_170), .w_ir_6_171(w_ir_6_171), .w_ir_6_172(w_ir_6_172), .w_ir_6_173(w_ir_6_173), .w_ir_6_174(w_ir_6_174), .w_ir_6_175(w_ir_6_175), .w_ir_6_176(w_ir_6_176), .w_ir_6_177(w_ir_6_177), .w_ir_6_178(w_ir_6_178), .w_ir_6_179(w_ir_6_179), .w_ir_6_180(w_ir_6_180), .w_ir_6_181(w_ir_6_181), .w_ir_6_182(w_ir_6_182), .w_ir_6_183(w_ir_6_183), .w_ir_6_184(w_ir_6_184), .w_ir_6_185(w_ir_6_185), .w_ir_6_186(w_ir_6_186), .w_ir_6_187(w_ir_6_187), .w_ir_6_188(w_ir_6_188), .w_ir_6_189(w_ir_6_189), .w_ir_6_190(w_ir_6_190), .w_ir_6_191(w_ir_6_191), .w_ir_6_192(w_ir_6_192), .w_ir_6_193(w_ir_6_193), .w_ir_6_194(w_ir_6_194), .w_ir_6_195(w_ir_6_195), .w_ir_6_196(w_ir_6_196), .w_ir_6_197(w_ir_6_197), .w_ir_6_198(w_ir_6_198), .w_ir_6_199(w_ir_6_199), .w_ir_6_200(w_ir_6_200), .w_ir_6_201(w_ir_6_201), .w_ir_6_202(w_ir_6_202), .w_ir_6_203(w_ir_6_203), .w_ir_6_204(w_ir_6_204), .w_ir_6_205(w_ir_6_205), .w_ir_6_206(w_ir_6_206), .w_ir_6_207(w_ir_6_207), .w_ir_6_208(w_ir_6_208), .w_ir_6_209(w_ir_6_209), .w_ir_6_210(w_ir_6_210), .w_ir_6_211(w_ir_6_211), .w_ir_6_212(w_ir_6_212), .w_ir_6_213(w_ir_6_213), .w_ir_6_214(w_ir_6_214), .w_ir_6_215(w_ir_6_215), .w_ir_6_216(w_ir_6_216), .w_ir_6_217(w_ir_6_217), .w_ir_6_218(w_ir_6_218), .w_ir_6_219(w_ir_6_219), .w_ir_6_220(w_ir_6_220), .w_ir_6_221(w_ir_6_221), .w_ir_6_222(w_ir_6_222), .w_ir_6_223(w_ir_6_223), .w_ir_6_224(w_ir_6_224), .w_ir_6_225(w_ir_6_225), .w_ir_6_226(w_ir_6_226), .w_ir_6_227(w_ir_6_227), .w_ir_6_228(w_ir_6_228), .w_ir_6_229(w_ir_6_229), .w_ir_6_230(w_ir_6_230), .w_ir_6_231(w_ir_6_231), .w_ir_6_232(w_ir_6_232), .w_ir_6_233(w_ir_6_233), .w_ir_6_234(w_ir_6_234), .w_ir_6_235(w_ir_6_235), .w_ir_6_236(w_ir_6_236), .w_ir_6_237(w_ir_6_237), .w_ir_6_238(w_ir_6_238), .w_ir_6_239(w_ir_6_239), .w_ir_6_240(w_ir_6_240), .w_ir_6_241(w_ir_6_241), .w_ir_6_242(w_ir_6_242), .w_ir_6_243(w_ir_6_243), .w_ir_6_244(w_ir_6_244), .w_ir_6_245(w_ir_6_245), .w_ir_6_246(w_ir_6_246), .w_ir_6_247(w_ir_6_247), .w_ir_6_248(w_ir_6_248), .w_ir_6_249(w_ir_6_249), .w_ir_6_250(w_ir_6_250), .w_ir_6_251(w_ir_6_251), .w_ir_6_252(w_ir_6_252), .w_ir_6_253(w_ir_6_253), .w_ir_6_254(w_ir_6_254), .w_ir_6_255(w_ir_6_255), .w_ir_7_0(w_ir_7_0), .w_ir_7_1(w_ir_7_1), .w_ir_7_2(w_ir_7_2), .w_ir_7_3(w_ir_7_3), .w_ir_7_4(w_ir_7_4), .w_ir_7_5(w_ir_7_5), .w_ir_7_6(w_ir_7_6), .w_ir_7_7(w_ir_7_7), .w_ir_7_8(w_ir_7_8), .w_ir_7_9(w_ir_7_9), .w_ir_7_10(w_ir_7_10), .w_ir_7_11(w_ir_7_11), .w_ir_7_12(w_ir_7_12), .w_ir_7_13(w_ir_7_13), .w_ir_7_14(w_ir_7_14), .w_ir_7_15(w_ir_7_15), .w_ir_7_16(w_ir_7_16), .w_ir_7_17(w_ir_7_17), .w_ir_7_18(w_ir_7_18), .w_ir_7_19(w_ir_7_19), .w_ir_7_20(w_ir_7_20), .w_ir_7_21(w_ir_7_21), .w_ir_7_22(w_ir_7_22), .w_ir_7_23(w_ir_7_23), .w_ir_7_24(w_ir_7_24), .w_ir_7_25(w_ir_7_25), .w_ir_7_26(w_ir_7_26), .w_ir_7_27(w_ir_7_27), .w_ir_7_28(w_ir_7_28), .w_ir_7_29(w_ir_7_29), .w_ir_7_30(w_ir_7_30), .w_ir_7_31(w_ir_7_31), .w_ir_7_32(w_ir_7_32), .w_ir_7_33(w_ir_7_33), .w_ir_7_34(w_ir_7_34), .w_ir_7_35(w_ir_7_35), .w_ir_7_36(w_ir_7_36), .w_ir_7_37(w_ir_7_37), .w_ir_7_38(w_ir_7_38), .w_ir_7_39(w_ir_7_39), .w_ir_7_40(w_ir_7_40), .w_ir_7_41(w_ir_7_41), .w_ir_7_42(w_ir_7_42), .w_ir_7_43(w_ir_7_43), .w_ir_7_44(w_ir_7_44), .w_ir_7_45(w_ir_7_45), .w_ir_7_46(w_ir_7_46), .w_ir_7_47(w_ir_7_47), .w_ir_7_48(w_ir_7_48), .w_ir_7_49(w_ir_7_49), .w_ir_7_50(w_ir_7_50), .w_ir_7_51(w_ir_7_51), .w_ir_7_52(w_ir_7_52), .w_ir_7_53(w_ir_7_53), .w_ir_7_54(w_ir_7_54), .w_ir_7_55(w_ir_7_55), .w_ir_7_56(w_ir_7_56), .w_ir_7_57(w_ir_7_57), .w_ir_7_58(w_ir_7_58), .w_ir_7_59(w_ir_7_59), .w_ir_7_60(w_ir_7_60), .w_ir_7_61(w_ir_7_61), .w_ir_7_62(w_ir_7_62), .w_ir_7_63(w_ir_7_63), .w_ir_7_64(w_ir_7_64), .w_ir_7_65(w_ir_7_65), .w_ir_7_66(w_ir_7_66), .w_ir_7_67(w_ir_7_67), .w_ir_7_68(w_ir_7_68), .w_ir_7_69(w_ir_7_69), .w_ir_7_70(w_ir_7_70), .w_ir_7_71(w_ir_7_71), .w_ir_7_72(w_ir_7_72), .w_ir_7_73(w_ir_7_73), .w_ir_7_74(w_ir_7_74), .w_ir_7_75(w_ir_7_75), .w_ir_7_76(w_ir_7_76), .w_ir_7_77(w_ir_7_77), .w_ir_7_78(w_ir_7_78), .w_ir_7_79(w_ir_7_79), .w_ir_7_80(w_ir_7_80), .w_ir_7_81(w_ir_7_81), .w_ir_7_82(w_ir_7_82), .w_ir_7_83(w_ir_7_83), .w_ir_7_84(w_ir_7_84), .w_ir_7_85(w_ir_7_85), .w_ir_7_86(w_ir_7_86), .w_ir_7_87(w_ir_7_87), .w_ir_7_88(w_ir_7_88), .w_ir_7_89(w_ir_7_89), .w_ir_7_90(w_ir_7_90), .w_ir_7_91(w_ir_7_91), .w_ir_7_92(w_ir_7_92), .w_ir_7_93(w_ir_7_93), .w_ir_7_94(w_ir_7_94), .w_ir_7_95(w_ir_7_95), .w_ir_7_96(w_ir_7_96), .w_ir_7_97(w_ir_7_97), .w_ir_7_98(w_ir_7_98), .w_ir_7_99(w_ir_7_99), .w_ir_7_100(w_ir_7_100), .w_ir_7_101(w_ir_7_101), .w_ir_7_102(w_ir_7_102), .w_ir_7_103(w_ir_7_103), .w_ir_7_104(w_ir_7_104), .w_ir_7_105(w_ir_7_105), .w_ir_7_106(w_ir_7_106), .w_ir_7_107(w_ir_7_107), .w_ir_7_108(w_ir_7_108), .w_ir_7_109(w_ir_7_109), .w_ir_7_110(w_ir_7_110), .w_ir_7_111(w_ir_7_111), .w_ir_7_112(w_ir_7_112), .w_ir_7_113(w_ir_7_113), .w_ir_7_114(w_ir_7_114), .w_ir_7_115(w_ir_7_115), .w_ir_7_116(w_ir_7_116), .w_ir_7_117(w_ir_7_117), .w_ir_7_118(w_ir_7_118), .w_ir_7_119(w_ir_7_119), .w_ir_7_120(w_ir_7_120), .w_ir_7_121(w_ir_7_121), .w_ir_7_122(w_ir_7_122), .w_ir_7_123(w_ir_7_123), .w_ir_7_124(w_ir_7_124), .w_ir_7_125(w_ir_7_125), .w_ir_7_126(w_ir_7_126), .w_ir_7_127(w_ir_7_127), .w_ir_7_128(w_ir_7_128), .w_ir_7_129(w_ir_7_129), .w_ir_7_130(w_ir_7_130), .w_ir_7_131(w_ir_7_131), .w_ir_7_132(w_ir_7_132), .w_ir_7_133(w_ir_7_133), .w_ir_7_134(w_ir_7_134), .w_ir_7_135(w_ir_7_135), .w_ir_7_136(w_ir_7_136), .w_ir_7_137(w_ir_7_137), .w_ir_7_138(w_ir_7_138), .w_ir_7_139(w_ir_7_139), .w_ir_7_140(w_ir_7_140), .w_ir_7_141(w_ir_7_141), .w_ir_7_142(w_ir_7_142), .w_ir_7_143(w_ir_7_143), .w_ir_7_144(w_ir_7_144), .w_ir_7_145(w_ir_7_145), .w_ir_7_146(w_ir_7_146), .w_ir_7_147(w_ir_7_147), .w_ir_7_148(w_ir_7_148), .w_ir_7_149(w_ir_7_149), .w_ir_7_150(w_ir_7_150), .w_ir_7_151(w_ir_7_151), .w_ir_7_152(w_ir_7_152), .w_ir_7_153(w_ir_7_153), .w_ir_7_154(w_ir_7_154), .w_ir_7_155(w_ir_7_155), .w_ir_7_156(w_ir_7_156), .w_ir_7_157(w_ir_7_157), .w_ir_7_158(w_ir_7_158), .w_ir_7_159(w_ir_7_159), .w_ir_7_160(w_ir_7_160), .w_ir_7_161(w_ir_7_161), .w_ir_7_162(w_ir_7_162), .w_ir_7_163(w_ir_7_163), .w_ir_7_164(w_ir_7_164), .w_ir_7_165(w_ir_7_165), .w_ir_7_166(w_ir_7_166), .w_ir_7_167(w_ir_7_167), .w_ir_7_168(w_ir_7_168), .w_ir_7_169(w_ir_7_169), .w_ir_7_170(w_ir_7_170), .w_ir_7_171(w_ir_7_171), .w_ir_7_172(w_ir_7_172), .w_ir_7_173(w_ir_7_173), .w_ir_7_174(w_ir_7_174), .w_ir_7_175(w_ir_7_175), .w_ir_7_176(w_ir_7_176), .w_ir_7_177(w_ir_7_177), .w_ir_7_178(w_ir_7_178), .w_ir_7_179(w_ir_7_179), .w_ir_7_180(w_ir_7_180), .w_ir_7_181(w_ir_7_181), .w_ir_7_182(w_ir_7_182), .w_ir_7_183(w_ir_7_183), .w_ir_7_184(w_ir_7_184), .w_ir_7_185(w_ir_7_185), .w_ir_7_186(w_ir_7_186), .w_ir_7_187(w_ir_7_187), .w_ir_7_188(w_ir_7_188), .w_ir_7_189(w_ir_7_189), .w_ir_7_190(w_ir_7_190), .w_ir_7_191(w_ir_7_191), .w_ir_7_192(w_ir_7_192), .w_ir_7_193(w_ir_7_193), .w_ir_7_194(w_ir_7_194), .w_ir_7_195(w_ir_7_195), .w_ir_7_196(w_ir_7_196), .w_ir_7_197(w_ir_7_197), .w_ir_7_198(w_ir_7_198), .w_ir_7_199(w_ir_7_199), .w_ir_7_200(w_ir_7_200), .w_ir_7_201(w_ir_7_201), .w_ir_7_202(w_ir_7_202), .w_ir_7_203(w_ir_7_203), .w_ir_7_204(w_ir_7_204), .w_ir_7_205(w_ir_7_205), .w_ir_7_206(w_ir_7_206), .w_ir_7_207(w_ir_7_207), .w_ir_7_208(w_ir_7_208), .w_ir_7_209(w_ir_7_209), .w_ir_7_210(w_ir_7_210), .w_ir_7_211(w_ir_7_211), .w_ir_7_212(w_ir_7_212), .w_ir_7_213(w_ir_7_213), .w_ir_7_214(w_ir_7_214), .w_ir_7_215(w_ir_7_215), .w_ir_7_216(w_ir_7_216), .w_ir_7_217(w_ir_7_217), .w_ir_7_218(w_ir_7_218), .w_ir_7_219(w_ir_7_219), .w_ir_7_220(w_ir_7_220), .w_ir_7_221(w_ir_7_221), .w_ir_7_222(w_ir_7_222), .w_ir_7_223(w_ir_7_223), .w_ir_7_224(w_ir_7_224), .w_ir_7_225(w_ir_7_225), .w_ir_7_226(w_ir_7_226), .w_ir_7_227(w_ir_7_227), .w_ir_7_228(w_ir_7_228), .w_ir_7_229(w_ir_7_229), .w_ir_7_230(w_ir_7_230), .w_ir_7_231(w_ir_7_231), .w_ir_7_232(w_ir_7_232), .w_ir_7_233(w_ir_7_233), .w_ir_7_234(w_ir_7_234), .w_ir_7_235(w_ir_7_235), .w_ir_7_236(w_ir_7_236), .w_ir_7_237(w_ir_7_237), .w_ir_7_238(w_ir_7_238), .w_ir_7_239(w_ir_7_239), .w_ir_7_240(w_ir_7_240), .w_ir_7_241(w_ir_7_241), .w_ir_7_242(w_ir_7_242), .w_ir_7_243(w_ir_7_243), .w_ir_7_244(w_ir_7_244), .w_ir_7_245(w_ir_7_245), .w_ir_7_246(w_ir_7_246), .w_ir_7_247(w_ir_7_247), .w_ir_7_248(w_ir_7_248), .w_ir_7_249(w_ir_7_249), .w_ir_7_250(w_ir_7_250), .w_ir_7_251(w_ir_7_251), .w_ir_7_252(w_ir_7_252), .w_ir_7_253(w_ir_7_253), .w_ir_7_254(w_ir_7_254), .w_ir_7_255(w_ir_7_255), 	
.w_iz_0_0(w_iz_0_0), .w_iz_0_1(w_iz_0_1), .w_iz_0_2(w_iz_0_2), .w_iz_0_3(w_iz_0_3), .w_iz_0_4(w_iz_0_4), .w_iz_0_5(w_iz_0_5), .w_iz_0_6(w_iz_0_6), .w_iz_0_7(w_iz_0_7), .w_iz_0_8(w_iz_0_8), .w_iz_0_9(w_iz_0_9), .w_iz_0_10(w_iz_0_10), .w_iz_0_11(w_iz_0_11), .w_iz_0_12(w_iz_0_12), .w_iz_0_13(w_iz_0_13), .w_iz_0_14(w_iz_0_14), .w_iz_0_15(w_iz_0_15), .w_iz_0_16(w_iz_0_16), .w_iz_0_17(w_iz_0_17), .w_iz_0_18(w_iz_0_18), .w_iz_0_19(w_iz_0_19), .w_iz_0_20(w_iz_0_20), .w_iz_0_21(w_iz_0_21), .w_iz_0_22(w_iz_0_22), .w_iz_0_23(w_iz_0_23), .w_iz_0_24(w_iz_0_24), .w_iz_0_25(w_iz_0_25), .w_iz_0_26(w_iz_0_26), .w_iz_0_27(w_iz_0_27), .w_iz_0_28(w_iz_0_28), .w_iz_0_29(w_iz_0_29), .w_iz_0_30(w_iz_0_30), .w_iz_0_31(w_iz_0_31), .w_iz_0_32(w_iz_0_32), .w_iz_0_33(w_iz_0_33), .w_iz_0_34(w_iz_0_34), .w_iz_0_35(w_iz_0_35), .w_iz_0_36(w_iz_0_36), .w_iz_0_37(w_iz_0_37), .w_iz_0_38(w_iz_0_38), .w_iz_0_39(w_iz_0_39), .w_iz_0_40(w_iz_0_40), .w_iz_0_41(w_iz_0_41), .w_iz_0_42(w_iz_0_42), .w_iz_0_43(w_iz_0_43), .w_iz_0_44(w_iz_0_44), .w_iz_0_45(w_iz_0_45), .w_iz_0_46(w_iz_0_46), .w_iz_0_47(w_iz_0_47), .w_iz_0_48(w_iz_0_48), .w_iz_0_49(w_iz_0_49), .w_iz_0_50(w_iz_0_50), .w_iz_0_51(w_iz_0_51), .w_iz_0_52(w_iz_0_52), .w_iz_0_53(w_iz_0_53), .w_iz_0_54(w_iz_0_54), .w_iz_0_55(w_iz_0_55), .w_iz_0_56(w_iz_0_56), .w_iz_0_57(w_iz_0_57), .w_iz_0_58(w_iz_0_58), .w_iz_0_59(w_iz_0_59), .w_iz_0_60(w_iz_0_60), .w_iz_0_61(w_iz_0_61), .w_iz_0_62(w_iz_0_62), .w_iz_0_63(w_iz_0_63), .w_iz_0_64(w_iz_0_64), .w_iz_0_65(w_iz_0_65), .w_iz_0_66(w_iz_0_66), .w_iz_0_67(w_iz_0_67), .w_iz_0_68(w_iz_0_68), .w_iz_0_69(w_iz_0_69), .w_iz_0_70(w_iz_0_70), .w_iz_0_71(w_iz_0_71), .w_iz_0_72(w_iz_0_72), .w_iz_0_73(w_iz_0_73), .w_iz_0_74(w_iz_0_74), .w_iz_0_75(w_iz_0_75), .w_iz_0_76(w_iz_0_76), .w_iz_0_77(w_iz_0_77), .w_iz_0_78(w_iz_0_78), .w_iz_0_79(w_iz_0_79), .w_iz_0_80(w_iz_0_80), .w_iz_0_81(w_iz_0_81), .w_iz_0_82(w_iz_0_82), .w_iz_0_83(w_iz_0_83), .w_iz_0_84(w_iz_0_84), .w_iz_0_85(w_iz_0_85), .w_iz_0_86(w_iz_0_86), .w_iz_0_87(w_iz_0_87), .w_iz_0_88(w_iz_0_88), .w_iz_0_89(w_iz_0_89), .w_iz_0_90(w_iz_0_90), .w_iz_0_91(w_iz_0_91), .w_iz_0_92(w_iz_0_92), .w_iz_0_93(w_iz_0_93), .w_iz_0_94(w_iz_0_94), .w_iz_0_95(w_iz_0_95), .w_iz_0_96(w_iz_0_96), .w_iz_0_97(w_iz_0_97), .w_iz_0_98(w_iz_0_98), .w_iz_0_99(w_iz_0_99), .w_iz_0_100(w_iz_0_100), .w_iz_0_101(w_iz_0_101), .w_iz_0_102(w_iz_0_102), .w_iz_0_103(w_iz_0_103), .w_iz_0_104(w_iz_0_104), .w_iz_0_105(w_iz_0_105), .w_iz_0_106(w_iz_0_106), .w_iz_0_107(w_iz_0_107), .w_iz_0_108(w_iz_0_108), .w_iz_0_109(w_iz_0_109), .w_iz_0_110(w_iz_0_110), .w_iz_0_111(w_iz_0_111), .w_iz_0_112(w_iz_0_112), .w_iz_0_113(w_iz_0_113), .w_iz_0_114(w_iz_0_114), .w_iz_0_115(w_iz_0_115), .w_iz_0_116(w_iz_0_116), .w_iz_0_117(w_iz_0_117), .w_iz_0_118(w_iz_0_118), .w_iz_0_119(w_iz_0_119), .w_iz_0_120(w_iz_0_120), .w_iz_0_121(w_iz_0_121), .w_iz_0_122(w_iz_0_122), .w_iz_0_123(w_iz_0_123), .w_iz_0_124(w_iz_0_124), .w_iz_0_125(w_iz_0_125), .w_iz_0_126(w_iz_0_126), .w_iz_0_127(w_iz_0_127), .w_iz_0_128(w_iz_0_128), .w_iz_0_129(w_iz_0_129), .w_iz_0_130(w_iz_0_130), .w_iz_0_131(w_iz_0_131), .w_iz_0_132(w_iz_0_132), .w_iz_0_133(w_iz_0_133), .w_iz_0_134(w_iz_0_134), .w_iz_0_135(w_iz_0_135), .w_iz_0_136(w_iz_0_136), .w_iz_0_137(w_iz_0_137), .w_iz_0_138(w_iz_0_138), .w_iz_0_139(w_iz_0_139), .w_iz_0_140(w_iz_0_140), .w_iz_0_141(w_iz_0_141), .w_iz_0_142(w_iz_0_142), .w_iz_0_143(w_iz_0_143), .w_iz_0_144(w_iz_0_144), .w_iz_0_145(w_iz_0_145), .w_iz_0_146(w_iz_0_146), .w_iz_0_147(w_iz_0_147), .w_iz_0_148(w_iz_0_148), .w_iz_0_149(w_iz_0_149), .w_iz_0_150(w_iz_0_150), .w_iz_0_151(w_iz_0_151), .w_iz_0_152(w_iz_0_152), .w_iz_0_153(w_iz_0_153), .w_iz_0_154(w_iz_0_154), .w_iz_0_155(w_iz_0_155), .w_iz_0_156(w_iz_0_156), .w_iz_0_157(w_iz_0_157), .w_iz_0_158(w_iz_0_158), .w_iz_0_159(w_iz_0_159), .w_iz_0_160(w_iz_0_160), .w_iz_0_161(w_iz_0_161), .w_iz_0_162(w_iz_0_162), .w_iz_0_163(w_iz_0_163), .w_iz_0_164(w_iz_0_164), .w_iz_0_165(w_iz_0_165), .w_iz_0_166(w_iz_0_166), .w_iz_0_167(w_iz_0_167), .w_iz_0_168(w_iz_0_168), .w_iz_0_169(w_iz_0_169), .w_iz_0_170(w_iz_0_170), .w_iz_0_171(w_iz_0_171), .w_iz_0_172(w_iz_0_172), .w_iz_0_173(w_iz_0_173), .w_iz_0_174(w_iz_0_174), .w_iz_0_175(w_iz_0_175), .w_iz_0_176(w_iz_0_176), .w_iz_0_177(w_iz_0_177), .w_iz_0_178(w_iz_0_178), .w_iz_0_179(w_iz_0_179), .w_iz_0_180(w_iz_0_180), .w_iz_0_181(w_iz_0_181), .w_iz_0_182(w_iz_0_182), .w_iz_0_183(w_iz_0_183), .w_iz_0_184(w_iz_0_184), .w_iz_0_185(w_iz_0_185), .w_iz_0_186(w_iz_0_186), .w_iz_0_187(w_iz_0_187), .w_iz_0_188(w_iz_0_188), .w_iz_0_189(w_iz_0_189), .w_iz_0_190(w_iz_0_190), .w_iz_0_191(w_iz_0_191), .w_iz_0_192(w_iz_0_192), .w_iz_0_193(w_iz_0_193), .w_iz_0_194(w_iz_0_194), .w_iz_0_195(w_iz_0_195), .w_iz_0_196(w_iz_0_196), .w_iz_0_197(w_iz_0_197), .w_iz_0_198(w_iz_0_198), .w_iz_0_199(w_iz_0_199), .w_iz_0_200(w_iz_0_200), .w_iz_0_201(w_iz_0_201), .w_iz_0_202(w_iz_0_202), .w_iz_0_203(w_iz_0_203), .w_iz_0_204(w_iz_0_204), .w_iz_0_205(w_iz_0_205), .w_iz_0_206(w_iz_0_206), .w_iz_0_207(w_iz_0_207), .w_iz_0_208(w_iz_0_208), .w_iz_0_209(w_iz_0_209), .w_iz_0_210(w_iz_0_210), .w_iz_0_211(w_iz_0_211), .w_iz_0_212(w_iz_0_212), .w_iz_0_213(w_iz_0_213), .w_iz_0_214(w_iz_0_214), .w_iz_0_215(w_iz_0_215), .w_iz_0_216(w_iz_0_216), .w_iz_0_217(w_iz_0_217), .w_iz_0_218(w_iz_0_218), .w_iz_0_219(w_iz_0_219), .w_iz_0_220(w_iz_0_220), .w_iz_0_221(w_iz_0_221), .w_iz_0_222(w_iz_0_222), .w_iz_0_223(w_iz_0_223), .w_iz_0_224(w_iz_0_224), .w_iz_0_225(w_iz_0_225), .w_iz_0_226(w_iz_0_226), .w_iz_0_227(w_iz_0_227), .w_iz_0_228(w_iz_0_228), .w_iz_0_229(w_iz_0_229), .w_iz_0_230(w_iz_0_230), .w_iz_0_231(w_iz_0_231), .w_iz_0_232(w_iz_0_232), .w_iz_0_233(w_iz_0_233), .w_iz_0_234(w_iz_0_234), .w_iz_0_235(w_iz_0_235), .w_iz_0_236(w_iz_0_236), .w_iz_0_237(w_iz_0_237), .w_iz_0_238(w_iz_0_238), .w_iz_0_239(w_iz_0_239), .w_iz_0_240(w_iz_0_240), .w_iz_0_241(w_iz_0_241), .w_iz_0_242(w_iz_0_242), .w_iz_0_243(w_iz_0_243), .w_iz_0_244(w_iz_0_244), .w_iz_0_245(w_iz_0_245), .w_iz_0_246(w_iz_0_246), .w_iz_0_247(w_iz_0_247), .w_iz_0_248(w_iz_0_248), .w_iz_0_249(w_iz_0_249), .w_iz_0_250(w_iz_0_250), .w_iz_0_251(w_iz_0_251), .w_iz_0_252(w_iz_0_252), .w_iz_0_253(w_iz_0_253), .w_iz_0_254(w_iz_0_254), .w_iz_0_255(w_iz_0_255), .w_iz_1_0(w_iz_1_0), .w_iz_1_1(w_iz_1_1), .w_iz_1_2(w_iz_1_2), .w_iz_1_3(w_iz_1_3), .w_iz_1_4(w_iz_1_4), .w_iz_1_5(w_iz_1_5), .w_iz_1_6(w_iz_1_6), .w_iz_1_7(w_iz_1_7), .w_iz_1_8(w_iz_1_8), .w_iz_1_9(w_iz_1_9), .w_iz_1_10(w_iz_1_10), .w_iz_1_11(w_iz_1_11), .w_iz_1_12(w_iz_1_12), .w_iz_1_13(w_iz_1_13), .w_iz_1_14(w_iz_1_14), .w_iz_1_15(w_iz_1_15), .w_iz_1_16(w_iz_1_16), .w_iz_1_17(w_iz_1_17), .w_iz_1_18(w_iz_1_18), .w_iz_1_19(w_iz_1_19), .w_iz_1_20(w_iz_1_20), .w_iz_1_21(w_iz_1_21), .w_iz_1_22(w_iz_1_22), .w_iz_1_23(w_iz_1_23), .w_iz_1_24(w_iz_1_24), .w_iz_1_25(w_iz_1_25), .w_iz_1_26(w_iz_1_26), .w_iz_1_27(w_iz_1_27), .w_iz_1_28(w_iz_1_28), .w_iz_1_29(w_iz_1_29), .w_iz_1_30(w_iz_1_30), .w_iz_1_31(w_iz_1_31), .w_iz_1_32(w_iz_1_32), .w_iz_1_33(w_iz_1_33), .w_iz_1_34(w_iz_1_34), .w_iz_1_35(w_iz_1_35), .w_iz_1_36(w_iz_1_36), .w_iz_1_37(w_iz_1_37), .w_iz_1_38(w_iz_1_38), .w_iz_1_39(w_iz_1_39), .w_iz_1_40(w_iz_1_40), .w_iz_1_41(w_iz_1_41), .w_iz_1_42(w_iz_1_42), .w_iz_1_43(w_iz_1_43), .w_iz_1_44(w_iz_1_44), .w_iz_1_45(w_iz_1_45), .w_iz_1_46(w_iz_1_46), .w_iz_1_47(w_iz_1_47), .w_iz_1_48(w_iz_1_48), .w_iz_1_49(w_iz_1_49), .w_iz_1_50(w_iz_1_50), .w_iz_1_51(w_iz_1_51), .w_iz_1_52(w_iz_1_52), .w_iz_1_53(w_iz_1_53), .w_iz_1_54(w_iz_1_54), .w_iz_1_55(w_iz_1_55), .w_iz_1_56(w_iz_1_56), .w_iz_1_57(w_iz_1_57), .w_iz_1_58(w_iz_1_58), .w_iz_1_59(w_iz_1_59), .w_iz_1_60(w_iz_1_60), .w_iz_1_61(w_iz_1_61), .w_iz_1_62(w_iz_1_62), .w_iz_1_63(w_iz_1_63), .w_iz_1_64(w_iz_1_64), .w_iz_1_65(w_iz_1_65), .w_iz_1_66(w_iz_1_66), .w_iz_1_67(w_iz_1_67), .w_iz_1_68(w_iz_1_68), .w_iz_1_69(w_iz_1_69), .w_iz_1_70(w_iz_1_70), .w_iz_1_71(w_iz_1_71), .w_iz_1_72(w_iz_1_72), .w_iz_1_73(w_iz_1_73), .w_iz_1_74(w_iz_1_74), .w_iz_1_75(w_iz_1_75), .w_iz_1_76(w_iz_1_76), .w_iz_1_77(w_iz_1_77), .w_iz_1_78(w_iz_1_78), .w_iz_1_79(w_iz_1_79), .w_iz_1_80(w_iz_1_80), .w_iz_1_81(w_iz_1_81), .w_iz_1_82(w_iz_1_82), .w_iz_1_83(w_iz_1_83), .w_iz_1_84(w_iz_1_84), .w_iz_1_85(w_iz_1_85), .w_iz_1_86(w_iz_1_86), .w_iz_1_87(w_iz_1_87), .w_iz_1_88(w_iz_1_88), .w_iz_1_89(w_iz_1_89), .w_iz_1_90(w_iz_1_90), .w_iz_1_91(w_iz_1_91), .w_iz_1_92(w_iz_1_92), .w_iz_1_93(w_iz_1_93), .w_iz_1_94(w_iz_1_94), .w_iz_1_95(w_iz_1_95), .w_iz_1_96(w_iz_1_96), .w_iz_1_97(w_iz_1_97), .w_iz_1_98(w_iz_1_98), .w_iz_1_99(w_iz_1_99), .w_iz_1_100(w_iz_1_100), .w_iz_1_101(w_iz_1_101), .w_iz_1_102(w_iz_1_102), .w_iz_1_103(w_iz_1_103), .w_iz_1_104(w_iz_1_104), .w_iz_1_105(w_iz_1_105), .w_iz_1_106(w_iz_1_106), .w_iz_1_107(w_iz_1_107), .w_iz_1_108(w_iz_1_108), .w_iz_1_109(w_iz_1_109), .w_iz_1_110(w_iz_1_110), .w_iz_1_111(w_iz_1_111), .w_iz_1_112(w_iz_1_112), .w_iz_1_113(w_iz_1_113), .w_iz_1_114(w_iz_1_114), .w_iz_1_115(w_iz_1_115), .w_iz_1_116(w_iz_1_116), .w_iz_1_117(w_iz_1_117), .w_iz_1_118(w_iz_1_118), .w_iz_1_119(w_iz_1_119), .w_iz_1_120(w_iz_1_120), .w_iz_1_121(w_iz_1_121), .w_iz_1_122(w_iz_1_122), .w_iz_1_123(w_iz_1_123), .w_iz_1_124(w_iz_1_124), .w_iz_1_125(w_iz_1_125), .w_iz_1_126(w_iz_1_126), .w_iz_1_127(w_iz_1_127), .w_iz_1_128(w_iz_1_128), .w_iz_1_129(w_iz_1_129), .w_iz_1_130(w_iz_1_130), .w_iz_1_131(w_iz_1_131), .w_iz_1_132(w_iz_1_132), .w_iz_1_133(w_iz_1_133), .w_iz_1_134(w_iz_1_134), .w_iz_1_135(w_iz_1_135), .w_iz_1_136(w_iz_1_136), .w_iz_1_137(w_iz_1_137), .w_iz_1_138(w_iz_1_138), .w_iz_1_139(w_iz_1_139), .w_iz_1_140(w_iz_1_140), .w_iz_1_141(w_iz_1_141), .w_iz_1_142(w_iz_1_142), .w_iz_1_143(w_iz_1_143), .w_iz_1_144(w_iz_1_144), .w_iz_1_145(w_iz_1_145), .w_iz_1_146(w_iz_1_146), .w_iz_1_147(w_iz_1_147), .w_iz_1_148(w_iz_1_148), .w_iz_1_149(w_iz_1_149), .w_iz_1_150(w_iz_1_150), .w_iz_1_151(w_iz_1_151), .w_iz_1_152(w_iz_1_152), .w_iz_1_153(w_iz_1_153), .w_iz_1_154(w_iz_1_154), .w_iz_1_155(w_iz_1_155), .w_iz_1_156(w_iz_1_156), .w_iz_1_157(w_iz_1_157), .w_iz_1_158(w_iz_1_158), .w_iz_1_159(w_iz_1_159), .w_iz_1_160(w_iz_1_160), .w_iz_1_161(w_iz_1_161), .w_iz_1_162(w_iz_1_162), .w_iz_1_163(w_iz_1_163), .w_iz_1_164(w_iz_1_164), .w_iz_1_165(w_iz_1_165), .w_iz_1_166(w_iz_1_166), .w_iz_1_167(w_iz_1_167), .w_iz_1_168(w_iz_1_168), .w_iz_1_169(w_iz_1_169), .w_iz_1_170(w_iz_1_170), .w_iz_1_171(w_iz_1_171), .w_iz_1_172(w_iz_1_172), .w_iz_1_173(w_iz_1_173), .w_iz_1_174(w_iz_1_174), .w_iz_1_175(w_iz_1_175), .w_iz_1_176(w_iz_1_176), .w_iz_1_177(w_iz_1_177), .w_iz_1_178(w_iz_1_178), .w_iz_1_179(w_iz_1_179), .w_iz_1_180(w_iz_1_180), .w_iz_1_181(w_iz_1_181), .w_iz_1_182(w_iz_1_182), .w_iz_1_183(w_iz_1_183), .w_iz_1_184(w_iz_1_184), .w_iz_1_185(w_iz_1_185), .w_iz_1_186(w_iz_1_186), .w_iz_1_187(w_iz_1_187), .w_iz_1_188(w_iz_1_188), .w_iz_1_189(w_iz_1_189), .w_iz_1_190(w_iz_1_190), .w_iz_1_191(w_iz_1_191), .w_iz_1_192(w_iz_1_192), .w_iz_1_193(w_iz_1_193), .w_iz_1_194(w_iz_1_194), .w_iz_1_195(w_iz_1_195), .w_iz_1_196(w_iz_1_196), .w_iz_1_197(w_iz_1_197), .w_iz_1_198(w_iz_1_198), .w_iz_1_199(w_iz_1_199), .w_iz_1_200(w_iz_1_200), .w_iz_1_201(w_iz_1_201), .w_iz_1_202(w_iz_1_202), .w_iz_1_203(w_iz_1_203), .w_iz_1_204(w_iz_1_204), .w_iz_1_205(w_iz_1_205), .w_iz_1_206(w_iz_1_206), .w_iz_1_207(w_iz_1_207), .w_iz_1_208(w_iz_1_208), .w_iz_1_209(w_iz_1_209), .w_iz_1_210(w_iz_1_210), .w_iz_1_211(w_iz_1_211), .w_iz_1_212(w_iz_1_212), .w_iz_1_213(w_iz_1_213), .w_iz_1_214(w_iz_1_214), .w_iz_1_215(w_iz_1_215), .w_iz_1_216(w_iz_1_216), .w_iz_1_217(w_iz_1_217), .w_iz_1_218(w_iz_1_218), .w_iz_1_219(w_iz_1_219), .w_iz_1_220(w_iz_1_220), .w_iz_1_221(w_iz_1_221), .w_iz_1_222(w_iz_1_222), .w_iz_1_223(w_iz_1_223), .w_iz_1_224(w_iz_1_224), .w_iz_1_225(w_iz_1_225), .w_iz_1_226(w_iz_1_226), .w_iz_1_227(w_iz_1_227), .w_iz_1_228(w_iz_1_228), .w_iz_1_229(w_iz_1_229), .w_iz_1_230(w_iz_1_230), .w_iz_1_231(w_iz_1_231), .w_iz_1_232(w_iz_1_232), .w_iz_1_233(w_iz_1_233), .w_iz_1_234(w_iz_1_234), .w_iz_1_235(w_iz_1_235), .w_iz_1_236(w_iz_1_236), .w_iz_1_237(w_iz_1_237), .w_iz_1_238(w_iz_1_238), .w_iz_1_239(w_iz_1_239), .w_iz_1_240(w_iz_1_240), .w_iz_1_241(w_iz_1_241), .w_iz_1_242(w_iz_1_242), .w_iz_1_243(w_iz_1_243), .w_iz_1_244(w_iz_1_244), .w_iz_1_245(w_iz_1_245), .w_iz_1_246(w_iz_1_246), .w_iz_1_247(w_iz_1_247), .w_iz_1_248(w_iz_1_248), .w_iz_1_249(w_iz_1_249), .w_iz_1_250(w_iz_1_250), .w_iz_1_251(w_iz_1_251), .w_iz_1_252(w_iz_1_252), .w_iz_1_253(w_iz_1_253), .w_iz_1_254(w_iz_1_254), .w_iz_1_255(w_iz_1_255), .w_iz_2_0(w_iz_2_0), .w_iz_2_1(w_iz_2_1), .w_iz_2_2(w_iz_2_2), .w_iz_2_3(w_iz_2_3), .w_iz_2_4(w_iz_2_4), .w_iz_2_5(w_iz_2_5), .w_iz_2_6(w_iz_2_6), .w_iz_2_7(w_iz_2_7), .w_iz_2_8(w_iz_2_8), .w_iz_2_9(w_iz_2_9), .w_iz_2_10(w_iz_2_10), .w_iz_2_11(w_iz_2_11), .w_iz_2_12(w_iz_2_12), .w_iz_2_13(w_iz_2_13), .w_iz_2_14(w_iz_2_14), .w_iz_2_15(w_iz_2_15), .w_iz_2_16(w_iz_2_16), .w_iz_2_17(w_iz_2_17), .w_iz_2_18(w_iz_2_18), .w_iz_2_19(w_iz_2_19), .w_iz_2_20(w_iz_2_20), .w_iz_2_21(w_iz_2_21), .w_iz_2_22(w_iz_2_22), .w_iz_2_23(w_iz_2_23), .w_iz_2_24(w_iz_2_24), .w_iz_2_25(w_iz_2_25), .w_iz_2_26(w_iz_2_26), .w_iz_2_27(w_iz_2_27), .w_iz_2_28(w_iz_2_28), .w_iz_2_29(w_iz_2_29), .w_iz_2_30(w_iz_2_30), .w_iz_2_31(w_iz_2_31), .w_iz_2_32(w_iz_2_32), .w_iz_2_33(w_iz_2_33), .w_iz_2_34(w_iz_2_34), .w_iz_2_35(w_iz_2_35), .w_iz_2_36(w_iz_2_36), .w_iz_2_37(w_iz_2_37), .w_iz_2_38(w_iz_2_38), .w_iz_2_39(w_iz_2_39), .w_iz_2_40(w_iz_2_40), .w_iz_2_41(w_iz_2_41), .w_iz_2_42(w_iz_2_42), .w_iz_2_43(w_iz_2_43), .w_iz_2_44(w_iz_2_44), .w_iz_2_45(w_iz_2_45), .w_iz_2_46(w_iz_2_46), .w_iz_2_47(w_iz_2_47), .w_iz_2_48(w_iz_2_48), .w_iz_2_49(w_iz_2_49), .w_iz_2_50(w_iz_2_50), .w_iz_2_51(w_iz_2_51), .w_iz_2_52(w_iz_2_52), .w_iz_2_53(w_iz_2_53), .w_iz_2_54(w_iz_2_54), .w_iz_2_55(w_iz_2_55), .w_iz_2_56(w_iz_2_56), .w_iz_2_57(w_iz_2_57), .w_iz_2_58(w_iz_2_58), .w_iz_2_59(w_iz_2_59), .w_iz_2_60(w_iz_2_60), .w_iz_2_61(w_iz_2_61), .w_iz_2_62(w_iz_2_62), .w_iz_2_63(w_iz_2_63), .w_iz_2_64(w_iz_2_64), .w_iz_2_65(w_iz_2_65), .w_iz_2_66(w_iz_2_66), .w_iz_2_67(w_iz_2_67), .w_iz_2_68(w_iz_2_68), .w_iz_2_69(w_iz_2_69), .w_iz_2_70(w_iz_2_70), .w_iz_2_71(w_iz_2_71), .w_iz_2_72(w_iz_2_72), .w_iz_2_73(w_iz_2_73), .w_iz_2_74(w_iz_2_74), .w_iz_2_75(w_iz_2_75), .w_iz_2_76(w_iz_2_76), .w_iz_2_77(w_iz_2_77), .w_iz_2_78(w_iz_2_78), .w_iz_2_79(w_iz_2_79), .w_iz_2_80(w_iz_2_80), .w_iz_2_81(w_iz_2_81), .w_iz_2_82(w_iz_2_82), .w_iz_2_83(w_iz_2_83), .w_iz_2_84(w_iz_2_84), .w_iz_2_85(w_iz_2_85), .w_iz_2_86(w_iz_2_86), .w_iz_2_87(w_iz_2_87), .w_iz_2_88(w_iz_2_88), .w_iz_2_89(w_iz_2_89), .w_iz_2_90(w_iz_2_90), .w_iz_2_91(w_iz_2_91), .w_iz_2_92(w_iz_2_92), .w_iz_2_93(w_iz_2_93), .w_iz_2_94(w_iz_2_94), .w_iz_2_95(w_iz_2_95), .w_iz_2_96(w_iz_2_96), .w_iz_2_97(w_iz_2_97), .w_iz_2_98(w_iz_2_98), .w_iz_2_99(w_iz_2_99), .w_iz_2_100(w_iz_2_100), .w_iz_2_101(w_iz_2_101), .w_iz_2_102(w_iz_2_102), .w_iz_2_103(w_iz_2_103), .w_iz_2_104(w_iz_2_104), .w_iz_2_105(w_iz_2_105), .w_iz_2_106(w_iz_2_106), .w_iz_2_107(w_iz_2_107), .w_iz_2_108(w_iz_2_108), .w_iz_2_109(w_iz_2_109), .w_iz_2_110(w_iz_2_110), .w_iz_2_111(w_iz_2_111), .w_iz_2_112(w_iz_2_112), .w_iz_2_113(w_iz_2_113), .w_iz_2_114(w_iz_2_114), .w_iz_2_115(w_iz_2_115), .w_iz_2_116(w_iz_2_116), .w_iz_2_117(w_iz_2_117), .w_iz_2_118(w_iz_2_118), .w_iz_2_119(w_iz_2_119), .w_iz_2_120(w_iz_2_120), .w_iz_2_121(w_iz_2_121), .w_iz_2_122(w_iz_2_122), .w_iz_2_123(w_iz_2_123), .w_iz_2_124(w_iz_2_124), .w_iz_2_125(w_iz_2_125), .w_iz_2_126(w_iz_2_126), .w_iz_2_127(w_iz_2_127), .w_iz_2_128(w_iz_2_128), .w_iz_2_129(w_iz_2_129), .w_iz_2_130(w_iz_2_130), .w_iz_2_131(w_iz_2_131), .w_iz_2_132(w_iz_2_132), .w_iz_2_133(w_iz_2_133), .w_iz_2_134(w_iz_2_134), .w_iz_2_135(w_iz_2_135), .w_iz_2_136(w_iz_2_136), .w_iz_2_137(w_iz_2_137), .w_iz_2_138(w_iz_2_138), .w_iz_2_139(w_iz_2_139), .w_iz_2_140(w_iz_2_140), .w_iz_2_141(w_iz_2_141), .w_iz_2_142(w_iz_2_142), .w_iz_2_143(w_iz_2_143), .w_iz_2_144(w_iz_2_144), .w_iz_2_145(w_iz_2_145), .w_iz_2_146(w_iz_2_146), .w_iz_2_147(w_iz_2_147), .w_iz_2_148(w_iz_2_148), .w_iz_2_149(w_iz_2_149), .w_iz_2_150(w_iz_2_150), .w_iz_2_151(w_iz_2_151), .w_iz_2_152(w_iz_2_152), .w_iz_2_153(w_iz_2_153), .w_iz_2_154(w_iz_2_154), .w_iz_2_155(w_iz_2_155), .w_iz_2_156(w_iz_2_156), .w_iz_2_157(w_iz_2_157), .w_iz_2_158(w_iz_2_158), .w_iz_2_159(w_iz_2_159), .w_iz_2_160(w_iz_2_160), .w_iz_2_161(w_iz_2_161), .w_iz_2_162(w_iz_2_162), .w_iz_2_163(w_iz_2_163), .w_iz_2_164(w_iz_2_164), .w_iz_2_165(w_iz_2_165), .w_iz_2_166(w_iz_2_166), .w_iz_2_167(w_iz_2_167), .w_iz_2_168(w_iz_2_168), .w_iz_2_169(w_iz_2_169), .w_iz_2_170(w_iz_2_170), .w_iz_2_171(w_iz_2_171), .w_iz_2_172(w_iz_2_172), .w_iz_2_173(w_iz_2_173), .w_iz_2_174(w_iz_2_174), .w_iz_2_175(w_iz_2_175), .w_iz_2_176(w_iz_2_176), .w_iz_2_177(w_iz_2_177), .w_iz_2_178(w_iz_2_178), .w_iz_2_179(w_iz_2_179), .w_iz_2_180(w_iz_2_180), .w_iz_2_181(w_iz_2_181), .w_iz_2_182(w_iz_2_182), .w_iz_2_183(w_iz_2_183), .w_iz_2_184(w_iz_2_184), .w_iz_2_185(w_iz_2_185), .w_iz_2_186(w_iz_2_186), .w_iz_2_187(w_iz_2_187), .w_iz_2_188(w_iz_2_188), .w_iz_2_189(w_iz_2_189), .w_iz_2_190(w_iz_2_190), .w_iz_2_191(w_iz_2_191), .w_iz_2_192(w_iz_2_192), .w_iz_2_193(w_iz_2_193), .w_iz_2_194(w_iz_2_194), .w_iz_2_195(w_iz_2_195), .w_iz_2_196(w_iz_2_196), .w_iz_2_197(w_iz_2_197), .w_iz_2_198(w_iz_2_198), .w_iz_2_199(w_iz_2_199), .w_iz_2_200(w_iz_2_200), .w_iz_2_201(w_iz_2_201), .w_iz_2_202(w_iz_2_202), .w_iz_2_203(w_iz_2_203), .w_iz_2_204(w_iz_2_204), .w_iz_2_205(w_iz_2_205), .w_iz_2_206(w_iz_2_206), .w_iz_2_207(w_iz_2_207), .w_iz_2_208(w_iz_2_208), .w_iz_2_209(w_iz_2_209), .w_iz_2_210(w_iz_2_210), .w_iz_2_211(w_iz_2_211), .w_iz_2_212(w_iz_2_212), .w_iz_2_213(w_iz_2_213), .w_iz_2_214(w_iz_2_214), .w_iz_2_215(w_iz_2_215), .w_iz_2_216(w_iz_2_216), .w_iz_2_217(w_iz_2_217), .w_iz_2_218(w_iz_2_218), .w_iz_2_219(w_iz_2_219), .w_iz_2_220(w_iz_2_220), .w_iz_2_221(w_iz_2_221), .w_iz_2_222(w_iz_2_222), .w_iz_2_223(w_iz_2_223), .w_iz_2_224(w_iz_2_224), .w_iz_2_225(w_iz_2_225), .w_iz_2_226(w_iz_2_226), .w_iz_2_227(w_iz_2_227), .w_iz_2_228(w_iz_2_228), .w_iz_2_229(w_iz_2_229), .w_iz_2_230(w_iz_2_230), .w_iz_2_231(w_iz_2_231), .w_iz_2_232(w_iz_2_232), .w_iz_2_233(w_iz_2_233), .w_iz_2_234(w_iz_2_234), .w_iz_2_235(w_iz_2_235), .w_iz_2_236(w_iz_2_236), .w_iz_2_237(w_iz_2_237), .w_iz_2_238(w_iz_2_238), .w_iz_2_239(w_iz_2_239), .w_iz_2_240(w_iz_2_240), .w_iz_2_241(w_iz_2_241), .w_iz_2_242(w_iz_2_242), .w_iz_2_243(w_iz_2_243), .w_iz_2_244(w_iz_2_244), .w_iz_2_245(w_iz_2_245), .w_iz_2_246(w_iz_2_246), .w_iz_2_247(w_iz_2_247), .w_iz_2_248(w_iz_2_248), .w_iz_2_249(w_iz_2_249), .w_iz_2_250(w_iz_2_250), .w_iz_2_251(w_iz_2_251), .w_iz_2_252(w_iz_2_252), .w_iz_2_253(w_iz_2_253), .w_iz_2_254(w_iz_2_254), .w_iz_2_255(w_iz_2_255), .w_iz_3_0(w_iz_3_0), .w_iz_3_1(w_iz_3_1), .w_iz_3_2(w_iz_3_2), .w_iz_3_3(w_iz_3_3), .w_iz_3_4(w_iz_3_4), .w_iz_3_5(w_iz_3_5), .w_iz_3_6(w_iz_3_6), .w_iz_3_7(w_iz_3_7), .w_iz_3_8(w_iz_3_8), .w_iz_3_9(w_iz_3_9), .w_iz_3_10(w_iz_3_10), .w_iz_3_11(w_iz_3_11), .w_iz_3_12(w_iz_3_12), .w_iz_3_13(w_iz_3_13), .w_iz_3_14(w_iz_3_14), .w_iz_3_15(w_iz_3_15), .w_iz_3_16(w_iz_3_16), .w_iz_3_17(w_iz_3_17), .w_iz_3_18(w_iz_3_18), .w_iz_3_19(w_iz_3_19), .w_iz_3_20(w_iz_3_20), .w_iz_3_21(w_iz_3_21), .w_iz_3_22(w_iz_3_22), .w_iz_3_23(w_iz_3_23), .w_iz_3_24(w_iz_3_24), .w_iz_3_25(w_iz_3_25), .w_iz_3_26(w_iz_3_26), .w_iz_3_27(w_iz_3_27), .w_iz_3_28(w_iz_3_28), .w_iz_3_29(w_iz_3_29), .w_iz_3_30(w_iz_3_30), .w_iz_3_31(w_iz_3_31), .w_iz_3_32(w_iz_3_32), .w_iz_3_33(w_iz_3_33), .w_iz_3_34(w_iz_3_34), .w_iz_3_35(w_iz_3_35), .w_iz_3_36(w_iz_3_36), .w_iz_3_37(w_iz_3_37), .w_iz_3_38(w_iz_3_38), .w_iz_3_39(w_iz_3_39), .w_iz_3_40(w_iz_3_40), .w_iz_3_41(w_iz_3_41), .w_iz_3_42(w_iz_3_42), .w_iz_3_43(w_iz_3_43), .w_iz_3_44(w_iz_3_44), .w_iz_3_45(w_iz_3_45), .w_iz_3_46(w_iz_3_46), .w_iz_3_47(w_iz_3_47), .w_iz_3_48(w_iz_3_48), .w_iz_3_49(w_iz_3_49), .w_iz_3_50(w_iz_3_50), .w_iz_3_51(w_iz_3_51), .w_iz_3_52(w_iz_3_52), .w_iz_3_53(w_iz_3_53), .w_iz_3_54(w_iz_3_54), .w_iz_3_55(w_iz_3_55), .w_iz_3_56(w_iz_3_56), .w_iz_3_57(w_iz_3_57), .w_iz_3_58(w_iz_3_58), .w_iz_3_59(w_iz_3_59), .w_iz_3_60(w_iz_3_60), .w_iz_3_61(w_iz_3_61), .w_iz_3_62(w_iz_3_62), .w_iz_3_63(w_iz_3_63), .w_iz_3_64(w_iz_3_64), .w_iz_3_65(w_iz_3_65), .w_iz_3_66(w_iz_3_66), .w_iz_3_67(w_iz_3_67), .w_iz_3_68(w_iz_3_68), .w_iz_3_69(w_iz_3_69), .w_iz_3_70(w_iz_3_70), .w_iz_3_71(w_iz_3_71), .w_iz_3_72(w_iz_3_72), .w_iz_3_73(w_iz_3_73), .w_iz_3_74(w_iz_3_74), .w_iz_3_75(w_iz_3_75), .w_iz_3_76(w_iz_3_76), .w_iz_3_77(w_iz_3_77), .w_iz_3_78(w_iz_3_78), .w_iz_3_79(w_iz_3_79), .w_iz_3_80(w_iz_3_80), .w_iz_3_81(w_iz_3_81), .w_iz_3_82(w_iz_3_82), .w_iz_3_83(w_iz_3_83), .w_iz_3_84(w_iz_3_84), .w_iz_3_85(w_iz_3_85), .w_iz_3_86(w_iz_3_86), .w_iz_3_87(w_iz_3_87), .w_iz_3_88(w_iz_3_88), .w_iz_3_89(w_iz_3_89), .w_iz_3_90(w_iz_3_90), .w_iz_3_91(w_iz_3_91), .w_iz_3_92(w_iz_3_92), .w_iz_3_93(w_iz_3_93), .w_iz_3_94(w_iz_3_94), .w_iz_3_95(w_iz_3_95), .w_iz_3_96(w_iz_3_96), .w_iz_3_97(w_iz_3_97), .w_iz_3_98(w_iz_3_98), .w_iz_3_99(w_iz_3_99), .w_iz_3_100(w_iz_3_100), .w_iz_3_101(w_iz_3_101), .w_iz_3_102(w_iz_3_102), .w_iz_3_103(w_iz_3_103), .w_iz_3_104(w_iz_3_104), .w_iz_3_105(w_iz_3_105), .w_iz_3_106(w_iz_3_106), .w_iz_3_107(w_iz_3_107), .w_iz_3_108(w_iz_3_108), .w_iz_3_109(w_iz_3_109), .w_iz_3_110(w_iz_3_110), .w_iz_3_111(w_iz_3_111), .w_iz_3_112(w_iz_3_112), .w_iz_3_113(w_iz_3_113), .w_iz_3_114(w_iz_3_114), .w_iz_3_115(w_iz_3_115), .w_iz_3_116(w_iz_3_116), .w_iz_3_117(w_iz_3_117), .w_iz_3_118(w_iz_3_118), .w_iz_3_119(w_iz_3_119), .w_iz_3_120(w_iz_3_120), .w_iz_3_121(w_iz_3_121), .w_iz_3_122(w_iz_3_122), .w_iz_3_123(w_iz_3_123), .w_iz_3_124(w_iz_3_124), .w_iz_3_125(w_iz_3_125), .w_iz_3_126(w_iz_3_126), .w_iz_3_127(w_iz_3_127), .w_iz_3_128(w_iz_3_128), .w_iz_3_129(w_iz_3_129), .w_iz_3_130(w_iz_3_130), .w_iz_3_131(w_iz_3_131), .w_iz_3_132(w_iz_3_132), .w_iz_3_133(w_iz_3_133), .w_iz_3_134(w_iz_3_134), .w_iz_3_135(w_iz_3_135), .w_iz_3_136(w_iz_3_136), .w_iz_3_137(w_iz_3_137), .w_iz_3_138(w_iz_3_138), .w_iz_3_139(w_iz_3_139), .w_iz_3_140(w_iz_3_140), .w_iz_3_141(w_iz_3_141), .w_iz_3_142(w_iz_3_142), .w_iz_3_143(w_iz_3_143), .w_iz_3_144(w_iz_3_144), .w_iz_3_145(w_iz_3_145), .w_iz_3_146(w_iz_3_146), .w_iz_3_147(w_iz_3_147), .w_iz_3_148(w_iz_3_148), .w_iz_3_149(w_iz_3_149), .w_iz_3_150(w_iz_3_150), .w_iz_3_151(w_iz_3_151), .w_iz_3_152(w_iz_3_152), .w_iz_3_153(w_iz_3_153), .w_iz_3_154(w_iz_3_154), .w_iz_3_155(w_iz_3_155), .w_iz_3_156(w_iz_3_156), .w_iz_3_157(w_iz_3_157), .w_iz_3_158(w_iz_3_158), .w_iz_3_159(w_iz_3_159), .w_iz_3_160(w_iz_3_160), .w_iz_3_161(w_iz_3_161), .w_iz_3_162(w_iz_3_162), .w_iz_3_163(w_iz_3_163), .w_iz_3_164(w_iz_3_164), .w_iz_3_165(w_iz_3_165), .w_iz_3_166(w_iz_3_166), .w_iz_3_167(w_iz_3_167), .w_iz_3_168(w_iz_3_168), .w_iz_3_169(w_iz_3_169), .w_iz_3_170(w_iz_3_170), .w_iz_3_171(w_iz_3_171), .w_iz_3_172(w_iz_3_172), .w_iz_3_173(w_iz_3_173), .w_iz_3_174(w_iz_3_174), .w_iz_3_175(w_iz_3_175), .w_iz_3_176(w_iz_3_176), .w_iz_3_177(w_iz_3_177), .w_iz_3_178(w_iz_3_178), .w_iz_3_179(w_iz_3_179), .w_iz_3_180(w_iz_3_180), .w_iz_3_181(w_iz_3_181), .w_iz_3_182(w_iz_3_182), .w_iz_3_183(w_iz_3_183), .w_iz_3_184(w_iz_3_184), .w_iz_3_185(w_iz_3_185), .w_iz_3_186(w_iz_3_186), .w_iz_3_187(w_iz_3_187), .w_iz_3_188(w_iz_3_188), .w_iz_3_189(w_iz_3_189), .w_iz_3_190(w_iz_3_190), .w_iz_3_191(w_iz_3_191), .w_iz_3_192(w_iz_3_192), .w_iz_3_193(w_iz_3_193), .w_iz_3_194(w_iz_3_194), .w_iz_3_195(w_iz_3_195), .w_iz_3_196(w_iz_3_196), .w_iz_3_197(w_iz_3_197), .w_iz_3_198(w_iz_3_198), .w_iz_3_199(w_iz_3_199), .w_iz_3_200(w_iz_3_200), .w_iz_3_201(w_iz_3_201), .w_iz_3_202(w_iz_3_202), .w_iz_3_203(w_iz_3_203), .w_iz_3_204(w_iz_3_204), .w_iz_3_205(w_iz_3_205), .w_iz_3_206(w_iz_3_206), .w_iz_3_207(w_iz_3_207), .w_iz_3_208(w_iz_3_208), .w_iz_3_209(w_iz_3_209), .w_iz_3_210(w_iz_3_210), .w_iz_3_211(w_iz_3_211), .w_iz_3_212(w_iz_3_212), .w_iz_3_213(w_iz_3_213), .w_iz_3_214(w_iz_3_214), .w_iz_3_215(w_iz_3_215), .w_iz_3_216(w_iz_3_216), .w_iz_3_217(w_iz_3_217), .w_iz_3_218(w_iz_3_218), .w_iz_3_219(w_iz_3_219), .w_iz_3_220(w_iz_3_220), .w_iz_3_221(w_iz_3_221), .w_iz_3_222(w_iz_3_222), .w_iz_3_223(w_iz_3_223), .w_iz_3_224(w_iz_3_224), .w_iz_3_225(w_iz_3_225), .w_iz_3_226(w_iz_3_226), .w_iz_3_227(w_iz_3_227), .w_iz_3_228(w_iz_3_228), .w_iz_3_229(w_iz_3_229), .w_iz_3_230(w_iz_3_230), .w_iz_3_231(w_iz_3_231), .w_iz_3_232(w_iz_3_232), .w_iz_3_233(w_iz_3_233), .w_iz_3_234(w_iz_3_234), .w_iz_3_235(w_iz_3_235), .w_iz_3_236(w_iz_3_236), .w_iz_3_237(w_iz_3_237), .w_iz_3_238(w_iz_3_238), .w_iz_3_239(w_iz_3_239), .w_iz_3_240(w_iz_3_240), .w_iz_3_241(w_iz_3_241), .w_iz_3_242(w_iz_3_242), .w_iz_3_243(w_iz_3_243), .w_iz_3_244(w_iz_3_244), .w_iz_3_245(w_iz_3_245), .w_iz_3_246(w_iz_3_246), .w_iz_3_247(w_iz_3_247), .w_iz_3_248(w_iz_3_248), .w_iz_3_249(w_iz_3_249), .w_iz_3_250(w_iz_3_250), .w_iz_3_251(w_iz_3_251), .w_iz_3_252(w_iz_3_252), .w_iz_3_253(w_iz_3_253), .w_iz_3_254(w_iz_3_254), .w_iz_3_255(w_iz_3_255), .w_iz_4_0(w_iz_4_0), .w_iz_4_1(w_iz_4_1), .w_iz_4_2(w_iz_4_2), .w_iz_4_3(w_iz_4_3), .w_iz_4_4(w_iz_4_4), .w_iz_4_5(w_iz_4_5), .w_iz_4_6(w_iz_4_6), .w_iz_4_7(w_iz_4_7), .w_iz_4_8(w_iz_4_8), .w_iz_4_9(w_iz_4_9), .w_iz_4_10(w_iz_4_10), .w_iz_4_11(w_iz_4_11), .w_iz_4_12(w_iz_4_12), .w_iz_4_13(w_iz_4_13), .w_iz_4_14(w_iz_4_14), .w_iz_4_15(w_iz_4_15), .w_iz_4_16(w_iz_4_16), .w_iz_4_17(w_iz_4_17), .w_iz_4_18(w_iz_4_18), .w_iz_4_19(w_iz_4_19), .w_iz_4_20(w_iz_4_20), .w_iz_4_21(w_iz_4_21), .w_iz_4_22(w_iz_4_22), .w_iz_4_23(w_iz_4_23), .w_iz_4_24(w_iz_4_24), .w_iz_4_25(w_iz_4_25), .w_iz_4_26(w_iz_4_26), .w_iz_4_27(w_iz_4_27), .w_iz_4_28(w_iz_4_28), .w_iz_4_29(w_iz_4_29), .w_iz_4_30(w_iz_4_30), .w_iz_4_31(w_iz_4_31), .w_iz_4_32(w_iz_4_32), .w_iz_4_33(w_iz_4_33), .w_iz_4_34(w_iz_4_34), .w_iz_4_35(w_iz_4_35), .w_iz_4_36(w_iz_4_36), .w_iz_4_37(w_iz_4_37), .w_iz_4_38(w_iz_4_38), .w_iz_4_39(w_iz_4_39), .w_iz_4_40(w_iz_4_40), .w_iz_4_41(w_iz_4_41), .w_iz_4_42(w_iz_4_42), .w_iz_4_43(w_iz_4_43), .w_iz_4_44(w_iz_4_44), .w_iz_4_45(w_iz_4_45), .w_iz_4_46(w_iz_4_46), .w_iz_4_47(w_iz_4_47), .w_iz_4_48(w_iz_4_48), .w_iz_4_49(w_iz_4_49), .w_iz_4_50(w_iz_4_50), .w_iz_4_51(w_iz_4_51), .w_iz_4_52(w_iz_4_52), .w_iz_4_53(w_iz_4_53), .w_iz_4_54(w_iz_4_54), .w_iz_4_55(w_iz_4_55), .w_iz_4_56(w_iz_4_56), .w_iz_4_57(w_iz_4_57), .w_iz_4_58(w_iz_4_58), .w_iz_4_59(w_iz_4_59), .w_iz_4_60(w_iz_4_60), .w_iz_4_61(w_iz_4_61), .w_iz_4_62(w_iz_4_62), .w_iz_4_63(w_iz_4_63), .w_iz_4_64(w_iz_4_64), .w_iz_4_65(w_iz_4_65), .w_iz_4_66(w_iz_4_66), .w_iz_4_67(w_iz_4_67), .w_iz_4_68(w_iz_4_68), .w_iz_4_69(w_iz_4_69), .w_iz_4_70(w_iz_4_70), .w_iz_4_71(w_iz_4_71), .w_iz_4_72(w_iz_4_72), .w_iz_4_73(w_iz_4_73), .w_iz_4_74(w_iz_4_74), .w_iz_4_75(w_iz_4_75), .w_iz_4_76(w_iz_4_76), .w_iz_4_77(w_iz_4_77), .w_iz_4_78(w_iz_4_78), .w_iz_4_79(w_iz_4_79), .w_iz_4_80(w_iz_4_80), .w_iz_4_81(w_iz_4_81), .w_iz_4_82(w_iz_4_82), .w_iz_4_83(w_iz_4_83), .w_iz_4_84(w_iz_4_84), .w_iz_4_85(w_iz_4_85), .w_iz_4_86(w_iz_4_86), .w_iz_4_87(w_iz_4_87), .w_iz_4_88(w_iz_4_88), .w_iz_4_89(w_iz_4_89), .w_iz_4_90(w_iz_4_90), .w_iz_4_91(w_iz_4_91), .w_iz_4_92(w_iz_4_92), .w_iz_4_93(w_iz_4_93), .w_iz_4_94(w_iz_4_94), .w_iz_4_95(w_iz_4_95), .w_iz_4_96(w_iz_4_96), .w_iz_4_97(w_iz_4_97), .w_iz_4_98(w_iz_4_98), .w_iz_4_99(w_iz_4_99), .w_iz_4_100(w_iz_4_100), .w_iz_4_101(w_iz_4_101), .w_iz_4_102(w_iz_4_102), .w_iz_4_103(w_iz_4_103), .w_iz_4_104(w_iz_4_104), .w_iz_4_105(w_iz_4_105), .w_iz_4_106(w_iz_4_106), .w_iz_4_107(w_iz_4_107), .w_iz_4_108(w_iz_4_108), .w_iz_4_109(w_iz_4_109), .w_iz_4_110(w_iz_4_110), .w_iz_4_111(w_iz_4_111), .w_iz_4_112(w_iz_4_112), .w_iz_4_113(w_iz_4_113), .w_iz_4_114(w_iz_4_114), .w_iz_4_115(w_iz_4_115), .w_iz_4_116(w_iz_4_116), .w_iz_4_117(w_iz_4_117), .w_iz_4_118(w_iz_4_118), .w_iz_4_119(w_iz_4_119), .w_iz_4_120(w_iz_4_120), .w_iz_4_121(w_iz_4_121), .w_iz_4_122(w_iz_4_122), .w_iz_4_123(w_iz_4_123), .w_iz_4_124(w_iz_4_124), .w_iz_4_125(w_iz_4_125), .w_iz_4_126(w_iz_4_126), .w_iz_4_127(w_iz_4_127), .w_iz_4_128(w_iz_4_128), .w_iz_4_129(w_iz_4_129), .w_iz_4_130(w_iz_4_130), .w_iz_4_131(w_iz_4_131), .w_iz_4_132(w_iz_4_132), .w_iz_4_133(w_iz_4_133), .w_iz_4_134(w_iz_4_134), .w_iz_4_135(w_iz_4_135), .w_iz_4_136(w_iz_4_136), .w_iz_4_137(w_iz_4_137), .w_iz_4_138(w_iz_4_138), .w_iz_4_139(w_iz_4_139), .w_iz_4_140(w_iz_4_140), .w_iz_4_141(w_iz_4_141), .w_iz_4_142(w_iz_4_142), .w_iz_4_143(w_iz_4_143), .w_iz_4_144(w_iz_4_144), .w_iz_4_145(w_iz_4_145), .w_iz_4_146(w_iz_4_146), .w_iz_4_147(w_iz_4_147), .w_iz_4_148(w_iz_4_148), .w_iz_4_149(w_iz_4_149), .w_iz_4_150(w_iz_4_150), .w_iz_4_151(w_iz_4_151), .w_iz_4_152(w_iz_4_152), .w_iz_4_153(w_iz_4_153), .w_iz_4_154(w_iz_4_154), .w_iz_4_155(w_iz_4_155), .w_iz_4_156(w_iz_4_156), .w_iz_4_157(w_iz_4_157), .w_iz_4_158(w_iz_4_158), .w_iz_4_159(w_iz_4_159), .w_iz_4_160(w_iz_4_160), .w_iz_4_161(w_iz_4_161), .w_iz_4_162(w_iz_4_162), .w_iz_4_163(w_iz_4_163), .w_iz_4_164(w_iz_4_164), .w_iz_4_165(w_iz_4_165), .w_iz_4_166(w_iz_4_166), .w_iz_4_167(w_iz_4_167), .w_iz_4_168(w_iz_4_168), .w_iz_4_169(w_iz_4_169), .w_iz_4_170(w_iz_4_170), .w_iz_4_171(w_iz_4_171), .w_iz_4_172(w_iz_4_172), .w_iz_4_173(w_iz_4_173), .w_iz_4_174(w_iz_4_174), .w_iz_4_175(w_iz_4_175), .w_iz_4_176(w_iz_4_176), .w_iz_4_177(w_iz_4_177), .w_iz_4_178(w_iz_4_178), .w_iz_4_179(w_iz_4_179), .w_iz_4_180(w_iz_4_180), .w_iz_4_181(w_iz_4_181), .w_iz_4_182(w_iz_4_182), .w_iz_4_183(w_iz_4_183), .w_iz_4_184(w_iz_4_184), .w_iz_4_185(w_iz_4_185), .w_iz_4_186(w_iz_4_186), .w_iz_4_187(w_iz_4_187), .w_iz_4_188(w_iz_4_188), .w_iz_4_189(w_iz_4_189), .w_iz_4_190(w_iz_4_190), .w_iz_4_191(w_iz_4_191), .w_iz_4_192(w_iz_4_192), .w_iz_4_193(w_iz_4_193), .w_iz_4_194(w_iz_4_194), .w_iz_4_195(w_iz_4_195), .w_iz_4_196(w_iz_4_196), .w_iz_4_197(w_iz_4_197), .w_iz_4_198(w_iz_4_198), .w_iz_4_199(w_iz_4_199), .w_iz_4_200(w_iz_4_200), .w_iz_4_201(w_iz_4_201), .w_iz_4_202(w_iz_4_202), .w_iz_4_203(w_iz_4_203), .w_iz_4_204(w_iz_4_204), .w_iz_4_205(w_iz_4_205), .w_iz_4_206(w_iz_4_206), .w_iz_4_207(w_iz_4_207), .w_iz_4_208(w_iz_4_208), .w_iz_4_209(w_iz_4_209), .w_iz_4_210(w_iz_4_210), .w_iz_4_211(w_iz_4_211), .w_iz_4_212(w_iz_4_212), .w_iz_4_213(w_iz_4_213), .w_iz_4_214(w_iz_4_214), .w_iz_4_215(w_iz_4_215), .w_iz_4_216(w_iz_4_216), .w_iz_4_217(w_iz_4_217), .w_iz_4_218(w_iz_4_218), .w_iz_4_219(w_iz_4_219), .w_iz_4_220(w_iz_4_220), .w_iz_4_221(w_iz_4_221), .w_iz_4_222(w_iz_4_222), .w_iz_4_223(w_iz_4_223), .w_iz_4_224(w_iz_4_224), .w_iz_4_225(w_iz_4_225), .w_iz_4_226(w_iz_4_226), .w_iz_4_227(w_iz_4_227), .w_iz_4_228(w_iz_4_228), .w_iz_4_229(w_iz_4_229), .w_iz_4_230(w_iz_4_230), .w_iz_4_231(w_iz_4_231), .w_iz_4_232(w_iz_4_232), .w_iz_4_233(w_iz_4_233), .w_iz_4_234(w_iz_4_234), .w_iz_4_235(w_iz_4_235), .w_iz_4_236(w_iz_4_236), .w_iz_4_237(w_iz_4_237), .w_iz_4_238(w_iz_4_238), .w_iz_4_239(w_iz_4_239), .w_iz_4_240(w_iz_4_240), .w_iz_4_241(w_iz_4_241), .w_iz_4_242(w_iz_4_242), .w_iz_4_243(w_iz_4_243), .w_iz_4_244(w_iz_4_244), .w_iz_4_245(w_iz_4_245), .w_iz_4_246(w_iz_4_246), .w_iz_4_247(w_iz_4_247), .w_iz_4_248(w_iz_4_248), .w_iz_4_249(w_iz_4_249), .w_iz_4_250(w_iz_4_250), .w_iz_4_251(w_iz_4_251), .w_iz_4_252(w_iz_4_252), .w_iz_4_253(w_iz_4_253), .w_iz_4_254(w_iz_4_254), .w_iz_4_255(w_iz_4_255), .w_iz_5_0(w_iz_5_0), .w_iz_5_1(w_iz_5_1), .w_iz_5_2(w_iz_5_2), .w_iz_5_3(w_iz_5_3), .w_iz_5_4(w_iz_5_4), .w_iz_5_5(w_iz_5_5), .w_iz_5_6(w_iz_5_6), .w_iz_5_7(w_iz_5_7), .w_iz_5_8(w_iz_5_8), .w_iz_5_9(w_iz_5_9), .w_iz_5_10(w_iz_5_10), .w_iz_5_11(w_iz_5_11), .w_iz_5_12(w_iz_5_12), .w_iz_5_13(w_iz_5_13), .w_iz_5_14(w_iz_5_14), .w_iz_5_15(w_iz_5_15), .w_iz_5_16(w_iz_5_16), .w_iz_5_17(w_iz_5_17), .w_iz_5_18(w_iz_5_18), .w_iz_5_19(w_iz_5_19), .w_iz_5_20(w_iz_5_20), .w_iz_5_21(w_iz_5_21), .w_iz_5_22(w_iz_5_22), .w_iz_5_23(w_iz_5_23), .w_iz_5_24(w_iz_5_24), .w_iz_5_25(w_iz_5_25), .w_iz_5_26(w_iz_5_26), .w_iz_5_27(w_iz_5_27), .w_iz_5_28(w_iz_5_28), .w_iz_5_29(w_iz_5_29), .w_iz_5_30(w_iz_5_30), .w_iz_5_31(w_iz_5_31), .w_iz_5_32(w_iz_5_32), .w_iz_5_33(w_iz_5_33), .w_iz_5_34(w_iz_5_34), .w_iz_5_35(w_iz_5_35), .w_iz_5_36(w_iz_5_36), .w_iz_5_37(w_iz_5_37), .w_iz_5_38(w_iz_5_38), .w_iz_5_39(w_iz_5_39), .w_iz_5_40(w_iz_5_40), .w_iz_5_41(w_iz_5_41), .w_iz_5_42(w_iz_5_42), .w_iz_5_43(w_iz_5_43), .w_iz_5_44(w_iz_5_44), .w_iz_5_45(w_iz_5_45), .w_iz_5_46(w_iz_5_46), .w_iz_5_47(w_iz_5_47), .w_iz_5_48(w_iz_5_48), .w_iz_5_49(w_iz_5_49), .w_iz_5_50(w_iz_5_50), .w_iz_5_51(w_iz_5_51), .w_iz_5_52(w_iz_5_52), .w_iz_5_53(w_iz_5_53), .w_iz_5_54(w_iz_5_54), .w_iz_5_55(w_iz_5_55), .w_iz_5_56(w_iz_5_56), .w_iz_5_57(w_iz_5_57), .w_iz_5_58(w_iz_5_58), .w_iz_5_59(w_iz_5_59), .w_iz_5_60(w_iz_5_60), .w_iz_5_61(w_iz_5_61), .w_iz_5_62(w_iz_5_62), .w_iz_5_63(w_iz_5_63), .w_iz_5_64(w_iz_5_64), .w_iz_5_65(w_iz_5_65), .w_iz_5_66(w_iz_5_66), .w_iz_5_67(w_iz_5_67), .w_iz_5_68(w_iz_5_68), .w_iz_5_69(w_iz_5_69), .w_iz_5_70(w_iz_5_70), .w_iz_5_71(w_iz_5_71), .w_iz_5_72(w_iz_5_72), .w_iz_5_73(w_iz_5_73), .w_iz_5_74(w_iz_5_74), .w_iz_5_75(w_iz_5_75), .w_iz_5_76(w_iz_5_76), .w_iz_5_77(w_iz_5_77), .w_iz_5_78(w_iz_5_78), .w_iz_5_79(w_iz_5_79), .w_iz_5_80(w_iz_5_80), .w_iz_5_81(w_iz_5_81), .w_iz_5_82(w_iz_5_82), .w_iz_5_83(w_iz_5_83), .w_iz_5_84(w_iz_5_84), .w_iz_5_85(w_iz_5_85), .w_iz_5_86(w_iz_5_86), .w_iz_5_87(w_iz_5_87), .w_iz_5_88(w_iz_5_88), .w_iz_5_89(w_iz_5_89), .w_iz_5_90(w_iz_5_90), .w_iz_5_91(w_iz_5_91), .w_iz_5_92(w_iz_5_92), .w_iz_5_93(w_iz_5_93), .w_iz_5_94(w_iz_5_94), .w_iz_5_95(w_iz_5_95), .w_iz_5_96(w_iz_5_96), .w_iz_5_97(w_iz_5_97), .w_iz_5_98(w_iz_5_98), .w_iz_5_99(w_iz_5_99), .w_iz_5_100(w_iz_5_100), .w_iz_5_101(w_iz_5_101), .w_iz_5_102(w_iz_5_102), .w_iz_5_103(w_iz_5_103), .w_iz_5_104(w_iz_5_104), .w_iz_5_105(w_iz_5_105), .w_iz_5_106(w_iz_5_106), .w_iz_5_107(w_iz_5_107), .w_iz_5_108(w_iz_5_108), .w_iz_5_109(w_iz_5_109), .w_iz_5_110(w_iz_5_110), .w_iz_5_111(w_iz_5_111), .w_iz_5_112(w_iz_5_112), .w_iz_5_113(w_iz_5_113), .w_iz_5_114(w_iz_5_114), .w_iz_5_115(w_iz_5_115), .w_iz_5_116(w_iz_5_116), .w_iz_5_117(w_iz_5_117), .w_iz_5_118(w_iz_5_118), .w_iz_5_119(w_iz_5_119), .w_iz_5_120(w_iz_5_120), .w_iz_5_121(w_iz_5_121), .w_iz_5_122(w_iz_5_122), .w_iz_5_123(w_iz_5_123), .w_iz_5_124(w_iz_5_124), .w_iz_5_125(w_iz_5_125), .w_iz_5_126(w_iz_5_126), .w_iz_5_127(w_iz_5_127), .w_iz_5_128(w_iz_5_128), .w_iz_5_129(w_iz_5_129), .w_iz_5_130(w_iz_5_130), .w_iz_5_131(w_iz_5_131), .w_iz_5_132(w_iz_5_132), .w_iz_5_133(w_iz_5_133), .w_iz_5_134(w_iz_5_134), .w_iz_5_135(w_iz_5_135), .w_iz_5_136(w_iz_5_136), .w_iz_5_137(w_iz_5_137), .w_iz_5_138(w_iz_5_138), .w_iz_5_139(w_iz_5_139), .w_iz_5_140(w_iz_5_140), .w_iz_5_141(w_iz_5_141), .w_iz_5_142(w_iz_5_142), .w_iz_5_143(w_iz_5_143), .w_iz_5_144(w_iz_5_144), .w_iz_5_145(w_iz_5_145), .w_iz_5_146(w_iz_5_146), .w_iz_5_147(w_iz_5_147), .w_iz_5_148(w_iz_5_148), .w_iz_5_149(w_iz_5_149), .w_iz_5_150(w_iz_5_150), .w_iz_5_151(w_iz_5_151), .w_iz_5_152(w_iz_5_152), .w_iz_5_153(w_iz_5_153), .w_iz_5_154(w_iz_5_154), .w_iz_5_155(w_iz_5_155), .w_iz_5_156(w_iz_5_156), .w_iz_5_157(w_iz_5_157), .w_iz_5_158(w_iz_5_158), .w_iz_5_159(w_iz_5_159), .w_iz_5_160(w_iz_5_160), .w_iz_5_161(w_iz_5_161), .w_iz_5_162(w_iz_5_162), .w_iz_5_163(w_iz_5_163), .w_iz_5_164(w_iz_5_164), .w_iz_5_165(w_iz_5_165), .w_iz_5_166(w_iz_5_166), .w_iz_5_167(w_iz_5_167), .w_iz_5_168(w_iz_5_168), .w_iz_5_169(w_iz_5_169), .w_iz_5_170(w_iz_5_170), .w_iz_5_171(w_iz_5_171), .w_iz_5_172(w_iz_5_172), .w_iz_5_173(w_iz_5_173), .w_iz_5_174(w_iz_5_174), .w_iz_5_175(w_iz_5_175), .w_iz_5_176(w_iz_5_176), .w_iz_5_177(w_iz_5_177), .w_iz_5_178(w_iz_5_178), .w_iz_5_179(w_iz_5_179), .w_iz_5_180(w_iz_5_180), .w_iz_5_181(w_iz_5_181), .w_iz_5_182(w_iz_5_182), .w_iz_5_183(w_iz_5_183), .w_iz_5_184(w_iz_5_184), .w_iz_5_185(w_iz_5_185), .w_iz_5_186(w_iz_5_186), .w_iz_5_187(w_iz_5_187), .w_iz_5_188(w_iz_5_188), .w_iz_5_189(w_iz_5_189), .w_iz_5_190(w_iz_5_190), .w_iz_5_191(w_iz_5_191), .w_iz_5_192(w_iz_5_192), .w_iz_5_193(w_iz_5_193), .w_iz_5_194(w_iz_5_194), .w_iz_5_195(w_iz_5_195), .w_iz_5_196(w_iz_5_196), .w_iz_5_197(w_iz_5_197), .w_iz_5_198(w_iz_5_198), .w_iz_5_199(w_iz_5_199), .w_iz_5_200(w_iz_5_200), .w_iz_5_201(w_iz_5_201), .w_iz_5_202(w_iz_5_202), .w_iz_5_203(w_iz_5_203), .w_iz_5_204(w_iz_5_204), .w_iz_5_205(w_iz_5_205), .w_iz_5_206(w_iz_5_206), .w_iz_5_207(w_iz_5_207), .w_iz_5_208(w_iz_5_208), .w_iz_5_209(w_iz_5_209), .w_iz_5_210(w_iz_5_210), .w_iz_5_211(w_iz_5_211), .w_iz_5_212(w_iz_5_212), .w_iz_5_213(w_iz_5_213), .w_iz_5_214(w_iz_5_214), .w_iz_5_215(w_iz_5_215), .w_iz_5_216(w_iz_5_216), .w_iz_5_217(w_iz_5_217), .w_iz_5_218(w_iz_5_218), .w_iz_5_219(w_iz_5_219), .w_iz_5_220(w_iz_5_220), .w_iz_5_221(w_iz_5_221), .w_iz_5_222(w_iz_5_222), .w_iz_5_223(w_iz_5_223), .w_iz_5_224(w_iz_5_224), .w_iz_5_225(w_iz_5_225), .w_iz_5_226(w_iz_5_226), .w_iz_5_227(w_iz_5_227), .w_iz_5_228(w_iz_5_228), .w_iz_5_229(w_iz_5_229), .w_iz_5_230(w_iz_5_230), .w_iz_5_231(w_iz_5_231), .w_iz_5_232(w_iz_5_232), .w_iz_5_233(w_iz_5_233), .w_iz_5_234(w_iz_5_234), .w_iz_5_235(w_iz_5_235), .w_iz_5_236(w_iz_5_236), .w_iz_5_237(w_iz_5_237), .w_iz_5_238(w_iz_5_238), .w_iz_5_239(w_iz_5_239), .w_iz_5_240(w_iz_5_240), .w_iz_5_241(w_iz_5_241), .w_iz_5_242(w_iz_5_242), .w_iz_5_243(w_iz_5_243), .w_iz_5_244(w_iz_5_244), .w_iz_5_245(w_iz_5_245), .w_iz_5_246(w_iz_5_246), .w_iz_5_247(w_iz_5_247), .w_iz_5_248(w_iz_5_248), .w_iz_5_249(w_iz_5_249), .w_iz_5_250(w_iz_5_250), .w_iz_5_251(w_iz_5_251), .w_iz_5_252(w_iz_5_252), .w_iz_5_253(w_iz_5_253), .w_iz_5_254(w_iz_5_254), .w_iz_5_255(w_iz_5_255), .w_iz_6_0(w_iz_6_0), .w_iz_6_1(w_iz_6_1), .w_iz_6_2(w_iz_6_2), .w_iz_6_3(w_iz_6_3), .w_iz_6_4(w_iz_6_4), .w_iz_6_5(w_iz_6_5), .w_iz_6_6(w_iz_6_6), .w_iz_6_7(w_iz_6_7), .w_iz_6_8(w_iz_6_8), .w_iz_6_9(w_iz_6_9), .w_iz_6_10(w_iz_6_10), .w_iz_6_11(w_iz_6_11), .w_iz_6_12(w_iz_6_12), .w_iz_6_13(w_iz_6_13), .w_iz_6_14(w_iz_6_14), .w_iz_6_15(w_iz_6_15), .w_iz_6_16(w_iz_6_16), .w_iz_6_17(w_iz_6_17), .w_iz_6_18(w_iz_6_18), .w_iz_6_19(w_iz_6_19), .w_iz_6_20(w_iz_6_20), .w_iz_6_21(w_iz_6_21), .w_iz_6_22(w_iz_6_22), .w_iz_6_23(w_iz_6_23), .w_iz_6_24(w_iz_6_24), .w_iz_6_25(w_iz_6_25), .w_iz_6_26(w_iz_6_26), .w_iz_6_27(w_iz_6_27), .w_iz_6_28(w_iz_6_28), .w_iz_6_29(w_iz_6_29), .w_iz_6_30(w_iz_6_30), .w_iz_6_31(w_iz_6_31), .w_iz_6_32(w_iz_6_32), .w_iz_6_33(w_iz_6_33), .w_iz_6_34(w_iz_6_34), .w_iz_6_35(w_iz_6_35), .w_iz_6_36(w_iz_6_36), .w_iz_6_37(w_iz_6_37), .w_iz_6_38(w_iz_6_38), .w_iz_6_39(w_iz_6_39), .w_iz_6_40(w_iz_6_40), .w_iz_6_41(w_iz_6_41), .w_iz_6_42(w_iz_6_42), .w_iz_6_43(w_iz_6_43), .w_iz_6_44(w_iz_6_44), .w_iz_6_45(w_iz_6_45), .w_iz_6_46(w_iz_6_46), .w_iz_6_47(w_iz_6_47), .w_iz_6_48(w_iz_6_48), .w_iz_6_49(w_iz_6_49), .w_iz_6_50(w_iz_6_50), .w_iz_6_51(w_iz_6_51), .w_iz_6_52(w_iz_6_52), .w_iz_6_53(w_iz_6_53), .w_iz_6_54(w_iz_6_54), .w_iz_6_55(w_iz_6_55), .w_iz_6_56(w_iz_6_56), .w_iz_6_57(w_iz_6_57), .w_iz_6_58(w_iz_6_58), .w_iz_6_59(w_iz_6_59), .w_iz_6_60(w_iz_6_60), .w_iz_6_61(w_iz_6_61), .w_iz_6_62(w_iz_6_62), .w_iz_6_63(w_iz_6_63), .w_iz_6_64(w_iz_6_64), .w_iz_6_65(w_iz_6_65), .w_iz_6_66(w_iz_6_66), .w_iz_6_67(w_iz_6_67), .w_iz_6_68(w_iz_6_68), .w_iz_6_69(w_iz_6_69), .w_iz_6_70(w_iz_6_70), .w_iz_6_71(w_iz_6_71), .w_iz_6_72(w_iz_6_72), .w_iz_6_73(w_iz_6_73), .w_iz_6_74(w_iz_6_74), .w_iz_6_75(w_iz_6_75), .w_iz_6_76(w_iz_6_76), .w_iz_6_77(w_iz_6_77), .w_iz_6_78(w_iz_6_78), .w_iz_6_79(w_iz_6_79), .w_iz_6_80(w_iz_6_80), .w_iz_6_81(w_iz_6_81), .w_iz_6_82(w_iz_6_82), .w_iz_6_83(w_iz_6_83), .w_iz_6_84(w_iz_6_84), .w_iz_6_85(w_iz_6_85), .w_iz_6_86(w_iz_6_86), .w_iz_6_87(w_iz_6_87), .w_iz_6_88(w_iz_6_88), .w_iz_6_89(w_iz_6_89), .w_iz_6_90(w_iz_6_90), .w_iz_6_91(w_iz_6_91), .w_iz_6_92(w_iz_6_92), .w_iz_6_93(w_iz_6_93), .w_iz_6_94(w_iz_6_94), .w_iz_6_95(w_iz_6_95), .w_iz_6_96(w_iz_6_96), .w_iz_6_97(w_iz_6_97), .w_iz_6_98(w_iz_6_98), .w_iz_6_99(w_iz_6_99), .w_iz_6_100(w_iz_6_100), .w_iz_6_101(w_iz_6_101), .w_iz_6_102(w_iz_6_102), .w_iz_6_103(w_iz_6_103), .w_iz_6_104(w_iz_6_104), .w_iz_6_105(w_iz_6_105), .w_iz_6_106(w_iz_6_106), .w_iz_6_107(w_iz_6_107), .w_iz_6_108(w_iz_6_108), .w_iz_6_109(w_iz_6_109), .w_iz_6_110(w_iz_6_110), .w_iz_6_111(w_iz_6_111), .w_iz_6_112(w_iz_6_112), .w_iz_6_113(w_iz_6_113), .w_iz_6_114(w_iz_6_114), .w_iz_6_115(w_iz_6_115), .w_iz_6_116(w_iz_6_116), .w_iz_6_117(w_iz_6_117), .w_iz_6_118(w_iz_6_118), .w_iz_6_119(w_iz_6_119), .w_iz_6_120(w_iz_6_120), .w_iz_6_121(w_iz_6_121), .w_iz_6_122(w_iz_6_122), .w_iz_6_123(w_iz_6_123), .w_iz_6_124(w_iz_6_124), .w_iz_6_125(w_iz_6_125), .w_iz_6_126(w_iz_6_126), .w_iz_6_127(w_iz_6_127), .w_iz_6_128(w_iz_6_128), .w_iz_6_129(w_iz_6_129), .w_iz_6_130(w_iz_6_130), .w_iz_6_131(w_iz_6_131), .w_iz_6_132(w_iz_6_132), .w_iz_6_133(w_iz_6_133), .w_iz_6_134(w_iz_6_134), .w_iz_6_135(w_iz_6_135), .w_iz_6_136(w_iz_6_136), .w_iz_6_137(w_iz_6_137), .w_iz_6_138(w_iz_6_138), .w_iz_6_139(w_iz_6_139), .w_iz_6_140(w_iz_6_140), .w_iz_6_141(w_iz_6_141), .w_iz_6_142(w_iz_6_142), .w_iz_6_143(w_iz_6_143), .w_iz_6_144(w_iz_6_144), .w_iz_6_145(w_iz_6_145), .w_iz_6_146(w_iz_6_146), .w_iz_6_147(w_iz_6_147), .w_iz_6_148(w_iz_6_148), .w_iz_6_149(w_iz_6_149), .w_iz_6_150(w_iz_6_150), .w_iz_6_151(w_iz_6_151), .w_iz_6_152(w_iz_6_152), .w_iz_6_153(w_iz_6_153), .w_iz_6_154(w_iz_6_154), .w_iz_6_155(w_iz_6_155), .w_iz_6_156(w_iz_6_156), .w_iz_6_157(w_iz_6_157), .w_iz_6_158(w_iz_6_158), .w_iz_6_159(w_iz_6_159), .w_iz_6_160(w_iz_6_160), .w_iz_6_161(w_iz_6_161), .w_iz_6_162(w_iz_6_162), .w_iz_6_163(w_iz_6_163), .w_iz_6_164(w_iz_6_164), .w_iz_6_165(w_iz_6_165), .w_iz_6_166(w_iz_6_166), .w_iz_6_167(w_iz_6_167), .w_iz_6_168(w_iz_6_168), .w_iz_6_169(w_iz_6_169), .w_iz_6_170(w_iz_6_170), .w_iz_6_171(w_iz_6_171), .w_iz_6_172(w_iz_6_172), .w_iz_6_173(w_iz_6_173), .w_iz_6_174(w_iz_6_174), .w_iz_6_175(w_iz_6_175), .w_iz_6_176(w_iz_6_176), .w_iz_6_177(w_iz_6_177), .w_iz_6_178(w_iz_6_178), .w_iz_6_179(w_iz_6_179), .w_iz_6_180(w_iz_6_180), .w_iz_6_181(w_iz_6_181), .w_iz_6_182(w_iz_6_182), .w_iz_6_183(w_iz_6_183), .w_iz_6_184(w_iz_6_184), .w_iz_6_185(w_iz_6_185), .w_iz_6_186(w_iz_6_186), .w_iz_6_187(w_iz_6_187), .w_iz_6_188(w_iz_6_188), .w_iz_6_189(w_iz_6_189), .w_iz_6_190(w_iz_6_190), .w_iz_6_191(w_iz_6_191), .w_iz_6_192(w_iz_6_192), .w_iz_6_193(w_iz_6_193), .w_iz_6_194(w_iz_6_194), .w_iz_6_195(w_iz_6_195), .w_iz_6_196(w_iz_6_196), .w_iz_6_197(w_iz_6_197), .w_iz_6_198(w_iz_6_198), .w_iz_6_199(w_iz_6_199), .w_iz_6_200(w_iz_6_200), .w_iz_6_201(w_iz_6_201), .w_iz_6_202(w_iz_6_202), .w_iz_6_203(w_iz_6_203), .w_iz_6_204(w_iz_6_204), .w_iz_6_205(w_iz_6_205), .w_iz_6_206(w_iz_6_206), .w_iz_6_207(w_iz_6_207), .w_iz_6_208(w_iz_6_208), .w_iz_6_209(w_iz_6_209), .w_iz_6_210(w_iz_6_210), .w_iz_6_211(w_iz_6_211), .w_iz_6_212(w_iz_6_212), .w_iz_6_213(w_iz_6_213), .w_iz_6_214(w_iz_6_214), .w_iz_6_215(w_iz_6_215), .w_iz_6_216(w_iz_6_216), .w_iz_6_217(w_iz_6_217), .w_iz_6_218(w_iz_6_218), .w_iz_6_219(w_iz_6_219), .w_iz_6_220(w_iz_6_220), .w_iz_6_221(w_iz_6_221), .w_iz_6_222(w_iz_6_222), .w_iz_6_223(w_iz_6_223), .w_iz_6_224(w_iz_6_224), .w_iz_6_225(w_iz_6_225), .w_iz_6_226(w_iz_6_226), .w_iz_6_227(w_iz_6_227), .w_iz_6_228(w_iz_6_228), .w_iz_6_229(w_iz_6_229), .w_iz_6_230(w_iz_6_230), .w_iz_6_231(w_iz_6_231), .w_iz_6_232(w_iz_6_232), .w_iz_6_233(w_iz_6_233), .w_iz_6_234(w_iz_6_234), .w_iz_6_235(w_iz_6_235), .w_iz_6_236(w_iz_6_236), .w_iz_6_237(w_iz_6_237), .w_iz_6_238(w_iz_6_238), .w_iz_6_239(w_iz_6_239), .w_iz_6_240(w_iz_6_240), .w_iz_6_241(w_iz_6_241), .w_iz_6_242(w_iz_6_242), .w_iz_6_243(w_iz_6_243), .w_iz_6_244(w_iz_6_244), .w_iz_6_245(w_iz_6_245), .w_iz_6_246(w_iz_6_246), .w_iz_6_247(w_iz_6_247), .w_iz_6_248(w_iz_6_248), .w_iz_6_249(w_iz_6_249), .w_iz_6_250(w_iz_6_250), .w_iz_6_251(w_iz_6_251), .w_iz_6_252(w_iz_6_252), .w_iz_6_253(w_iz_6_253), .w_iz_6_254(w_iz_6_254), .w_iz_6_255(w_iz_6_255), .w_iz_7_0(w_iz_7_0), .w_iz_7_1(w_iz_7_1), .w_iz_7_2(w_iz_7_2), .w_iz_7_3(w_iz_7_3), .w_iz_7_4(w_iz_7_4), .w_iz_7_5(w_iz_7_5), .w_iz_7_6(w_iz_7_6), .w_iz_7_7(w_iz_7_7), .w_iz_7_8(w_iz_7_8), .w_iz_7_9(w_iz_7_9), .w_iz_7_10(w_iz_7_10), .w_iz_7_11(w_iz_7_11), .w_iz_7_12(w_iz_7_12), .w_iz_7_13(w_iz_7_13), .w_iz_7_14(w_iz_7_14), .w_iz_7_15(w_iz_7_15), .w_iz_7_16(w_iz_7_16), .w_iz_7_17(w_iz_7_17), .w_iz_7_18(w_iz_7_18), .w_iz_7_19(w_iz_7_19), .w_iz_7_20(w_iz_7_20), .w_iz_7_21(w_iz_7_21), .w_iz_7_22(w_iz_7_22), .w_iz_7_23(w_iz_7_23), .w_iz_7_24(w_iz_7_24), .w_iz_7_25(w_iz_7_25), .w_iz_7_26(w_iz_7_26), .w_iz_7_27(w_iz_7_27), .w_iz_7_28(w_iz_7_28), .w_iz_7_29(w_iz_7_29), .w_iz_7_30(w_iz_7_30), .w_iz_7_31(w_iz_7_31), .w_iz_7_32(w_iz_7_32), .w_iz_7_33(w_iz_7_33), .w_iz_7_34(w_iz_7_34), .w_iz_7_35(w_iz_7_35), .w_iz_7_36(w_iz_7_36), .w_iz_7_37(w_iz_7_37), .w_iz_7_38(w_iz_7_38), .w_iz_7_39(w_iz_7_39), .w_iz_7_40(w_iz_7_40), .w_iz_7_41(w_iz_7_41), .w_iz_7_42(w_iz_7_42), .w_iz_7_43(w_iz_7_43), .w_iz_7_44(w_iz_7_44), .w_iz_7_45(w_iz_7_45), .w_iz_7_46(w_iz_7_46), .w_iz_7_47(w_iz_7_47), .w_iz_7_48(w_iz_7_48), .w_iz_7_49(w_iz_7_49), .w_iz_7_50(w_iz_7_50), .w_iz_7_51(w_iz_7_51), .w_iz_7_52(w_iz_7_52), .w_iz_7_53(w_iz_7_53), .w_iz_7_54(w_iz_7_54), .w_iz_7_55(w_iz_7_55), .w_iz_7_56(w_iz_7_56), .w_iz_7_57(w_iz_7_57), .w_iz_7_58(w_iz_7_58), .w_iz_7_59(w_iz_7_59), .w_iz_7_60(w_iz_7_60), .w_iz_7_61(w_iz_7_61), .w_iz_7_62(w_iz_7_62), .w_iz_7_63(w_iz_7_63), .w_iz_7_64(w_iz_7_64), .w_iz_7_65(w_iz_7_65), .w_iz_7_66(w_iz_7_66), .w_iz_7_67(w_iz_7_67), .w_iz_7_68(w_iz_7_68), .w_iz_7_69(w_iz_7_69), .w_iz_7_70(w_iz_7_70), .w_iz_7_71(w_iz_7_71), .w_iz_7_72(w_iz_7_72), .w_iz_7_73(w_iz_7_73), .w_iz_7_74(w_iz_7_74), .w_iz_7_75(w_iz_7_75), .w_iz_7_76(w_iz_7_76), .w_iz_7_77(w_iz_7_77), .w_iz_7_78(w_iz_7_78), .w_iz_7_79(w_iz_7_79), .w_iz_7_80(w_iz_7_80), .w_iz_7_81(w_iz_7_81), .w_iz_7_82(w_iz_7_82), .w_iz_7_83(w_iz_7_83), .w_iz_7_84(w_iz_7_84), .w_iz_7_85(w_iz_7_85), .w_iz_7_86(w_iz_7_86), .w_iz_7_87(w_iz_7_87), .w_iz_7_88(w_iz_7_88), .w_iz_7_89(w_iz_7_89), .w_iz_7_90(w_iz_7_90), .w_iz_7_91(w_iz_7_91), .w_iz_7_92(w_iz_7_92), .w_iz_7_93(w_iz_7_93), .w_iz_7_94(w_iz_7_94), .w_iz_7_95(w_iz_7_95), .w_iz_7_96(w_iz_7_96), .w_iz_7_97(w_iz_7_97), .w_iz_7_98(w_iz_7_98), .w_iz_7_99(w_iz_7_99), .w_iz_7_100(w_iz_7_100), .w_iz_7_101(w_iz_7_101), .w_iz_7_102(w_iz_7_102), .w_iz_7_103(w_iz_7_103), .w_iz_7_104(w_iz_7_104), .w_iz_7_105(w_iz_7_105), .w_iz_7_106(w_iz_7_106), .w_iz_7_107(w_iz_7_107), .w_iz_7_108(w_iz_7_108), .w_iz_7_109(w_iz_7_109), .w_iz_7_110(w_iz_7_110), .w_iz_7_111(w_iz_7_111), .w_iz_7_112(w_iz_7_112), .w_iz_7_113(w_iz_7_113), .w_iz_7_114(w_iz_7_114), .w_iz_7_115(w_iz_7_115), .w_iz_7_116(w_iz_7_116), .w_iz_7_117(w_iz_7_117), .w_iz_7_118(w_iz_7_118), .w_iz_7_119(w_iz_7_119), .w_iz_7_120(w_iz_7_120), .w_iz_7_121(w_iz_7_121), .w_iz_7_122(w_iz_7_122), .w_iz_7_123(w_iz_7_123), .w_iz_7_124(w_iz_7_124), .w_iz_7_125(w_iz_7_125), .w_iz_7_126(w_iz_7_126), .w_iz_7_127(w_iz_7_127), .w_iz_7_128(w_iz_7_128), .w_iz_7_129(w_iz_7_129), .w_iz_7_130(w_iz_7_130), .w_iz_7_131(w_iz_7_131), .w_iz_7_132(w_iz_7_132), .w_iz_7_133(w_iz_7_133), .w_iz_7_134(w_iz_7_134), .w_iz_7_135(w_iz_7_135), .w_iz_7_136(w_iz_7_136), .w_iz_7_137(w_iz_7_137), .w_iz_7_138(w_iz_7_138), .w_iz_7_139(w_iz_7_139), .w_iz_7_140(w_iz_7_140), .w_iz_7_141(w_iz_7_141), .w_iz_7_142(w_iz_7_142), .w_iz_7_143(w_iz_7_143), .w_iz_7_144(w_iz_7_144), .w_iz_7_145(w_iz_7_145), .w_iz_7_146(w_iz_7_146), .w_iz_7_147(w_iz_7_147), .w_iz_7_148(w_iz_7_148), .w_iz_7_149(w_iz_7_149), .w_iz_7_150(w_iz_7_150), .w_iz_7_151(w_iz_7_151), .w_iz_7_152(w_iz_7_152), .w_iz_7_153(w_iz_7_153), .w_iz_7_154(w_iz_7_154), .w_iz_7_155(w_iz_7_155), .w_iz_7_156(w_iz_7_156), .w_iz_7_157(w_iz_7_157), .w_iz_7_158(w_iz_7_158), .w_iz_7_159(w_iz_7_159), .w_iz_7_160(w_iz_7_160), .w_iz_7_161(w_iz_7_161), .w_iz_7_162(w_iz_7_162), .w_iz_7_163(w_iz_7_163), .w_iz_7_164(w_iz_7_164), .w_iz_7_165(w_iz_7_165), .w_iz_7_166(w_iz_7_166), .w_iz_7_167(w_iz_7_167), .w_iz_7_168(w_iz_7_168), .w_iz_7_169(w_iz_7_169), .w_iz_7_170(w_iz_7_170), .w_iz_7_171(w_iz_7_171), .w_iz_7_172(w_iz_7_172), .w_iz_7_173(w_iz_7_173), .w_iz_7_174(w_iz_7_174), .w_iz_7_175(w_iz_7_175), .w_iz_7_176(w_iz_7_176), .w_iz_7_177(w_iz_7_177), .w_iz_7_178(w_iz_7_178), .w_iz_7_179(w_iz_7_179), .w_iz_7_180(w_iz_7_180), .w_iz_7_181(w_iz_7_181), .w_iz_7_182(w_iz_7_182), .w_iz_7_183(w_iz_7_183), .w_iz_7_184(w_iz_7_184), .w_iz_7_185(w_iz_7_185), .w_iz_7_186(w_iz_7_186), .w_iz_7_187(w_iz_7_187), .w_iz_7_188(w_iz_7_188), .w_iz_7_189(w_iz_7_189), .w_iz_7_190(w_iz_7_190), .w_iz_7_191(w_iz_7_191), .w_iz_7_192(w_iz_7_192), .w_iz_7_193(w_iz_7_193), .w_iz_7_194(w_iz_7_194), .w_iz_7_195(w_iz_7_195), .w_iz_7_196(w_iz_7_196), .w_iz_7_197(w_iz_7_197), .w_iz_7_198(w_iz_7_198), .w_iz_7_199(w_iz_7_199), .w_iz_7_200(w_iz_7_200), .w_iz_7_201(w_iz_7_201), .w_iz_7_202(w_iz_7_202), .w_iz_7_203(w_iz_7_203), .w_iz_7_204(w_iz_7_204), .w_iz_7_205(w_iz_7_205), .w_iz_7_206(w_iz_7_206), .w_iz_7_207(w_iz_7_207), .w_iz_7_208(w_iz_7_208), .w_iz_7_209(w_iz_7_209), .w_iz_7_210(w_iz_7_210), .w_iz_7_211(w_iz_7_211), .w_iz_7_212(w_iz_7_212), .w_iz_7_213(w_iz_7_213), .w_iz_7_214(w_iz_7_214), .w_iz_7_215(w_iz_7_215), .w_iz_7_216(w_iz_7_216), .w_iz_7_217(w_iz_7_217), .w_iz_7_218(w_iz_7_218), .w_iz_7_219(w_iz_7_219), .w_iz_7_220(w_iz_7_220), .w_iz_7_221(w_iz_7_221), .w_iz_7_222(w_iz_7_222), .w_iz_7_223(w_iz_7_223), .w_iz_7_224(w_iz_7_224), .w_iz_7_225(w_iz_7_225), .w_iz_7_226(w_iz_7_226), .w_iz_7_227(w_iz_7_227), .w_iz_7_228(w_iz_7_228), .w_iz_7_229(w_iz_7_229), .w_iz_7_230(w_iz_7_230), .w_iz_7_231(w_iz_7_231), .w_iz_7_232(w_iz_7_232), .w_iz_7_233(w_iz_7_233), .w_iz_7_234(w_iz_7_234), .w_iz_7_235(w_iz_7_235), .w_iz_7_236(w_iz_7_236), .w_iz_7_237(w_iz_7_237), .w_iz_7_238(w_iz_7_238), .w_iz_7_239(w_iz_7_239), .w_iz_7_240(w_iz_7_240), .w_iz_7_241(w_iz_7_241), .w_iz_7_242(w_iz_7_242), .w_iz_7_243(w_iz_7_243), .w_iz_7_244(w_iz_7_244), .w_iz_7_245(w_iz_7_245), .w_iz_7_246(w_iz_7_246), .w_iz_7_247(w_iz_7_247), .w_iz_7_248(w_iz_7_248), .w_iz_7_249(w_iz_7_249), .w_iz_7_250(w_iz_7_250), .w_iz_7_251(w_iz_7_251), .w_iz_7_252(w_iz_7_252), .w_iz_7_253(w_iz_7_253), .w_iz_7_254(w_iz_7_254), .w_iz_7_255(w_iz_7_255), 
.w_in_0_0(w_in_0_0), .w_in_0_1(w_in_0_1), .w_in_0_2(w_in_0_2), .w_in_0_3(w_in_0_3), .w_in_0_4(w_in_0_4), .w_in_0_5(w_in_0_5), .w_in_0_6(w_in_0_6), .w_in_0_7(w_in_0_7), .w_in_0_8(w_in_0_8), .w_in_0_9(w_in_0_9), .w_in_0_10(w_in_0_10), .w_in_0_11(w_in_0_11), .w_in_0_12(w_in_0_12), .w_in_0_13(w_in_0_13), .w_in_0_14(w_in_0_14), .w_in_0_15(w_in_0_15), .w_in_0_16(w_in_0_16), .w_in_0_17(w_in_0_17), .w_in_0_18(w_in_0_18), .w_in_0_19(w_in_0_19), .w_in_0_20(w_in_0_20), .w_in_0_21(w_in_0_21), .w_in_0_22(w_in_0_22), .w_in_0_23(w_in_0_23), .w_in_0_24(w_in_0_24), .w_in_0_25(w_in_0_25), .w_in_0_26(w_in_0_26), .w_in_0_27(w_in_0_27), .w_in_0_28(w_in_0_28), .w_in_0_29(w_in_0_29), .w_in_0_30(w_in_0_30), .w_in_0_31(w_in_0_31), .w_in_0_32(w_in_0_32), .w_in_0_33(w_in_0_33), .w_in_0_34(w_in_0_34), .w_in_0_35(w_in_0_35), .w_in_0_36(w_in_0_36), .w_in_0_37(w_in_0_37), .w_in_0_38(w_in_0_38), .w_in_0_39(w_in_0_39), .w_in_0_40(w_in_0_40), .w_in_0_41(w_in_0_41), .w_in_0_42(w_in_0_42), .w_in_0_43(w_in_0_43), .w_in_0_44(w_in_0_44), .w_in_0_45(w_in_0_45), .w_in_0_46(w_in_0_46), .w_in_0_47(w_in_0_47), .w_in_0_48(w_in_0_48), .w_in_0_49(w_in_0_49), .w_in_0_50(w_in_0_50), .w_in_0_51(w_in_0_51), .w_in_0_52(w_in_0_52), .w_in_0_53(w_in_0_53), .w_in_0_54(w_in_0_54), .w_in_0_55(w_in_0_55), .w_in_0_56(w_in_0_56), .w_in_0_57(w_in_0_57), .w_in_0_58(w_in_0_58), .w_in_0_59(w_in_0_59), .w_in_0_60(w_in_0_60), .w_in_0_61(w_in_0_61), .w_in_0_62(w_in_0_62), .w_in_0_63(w_in_0_63), .w_in_0_64(w_in_0_64), .w_in_0_65(w_in_0_65), .w_in_0_66(w_in_0_66), .w_in_0_67(w_in_0_67), .w_in_0_68(w_in_0_68), .w_in_0_69(w_in_0_69), .w_in_0_70(w_in_0_70), .w_in_0_71(w_in_0_71), .w_in_0_72(w_in_0_72), .w_in_0_73(w_in_0_73), .w_in_0_74(w_in_0_74), .w_in_0_75(w_in_0_75), .w_in_0_76(w_in_0_76), .w_in_0_77(w_in_0_77), .w_in_0_78(w_in_0_78), .w_in_0_79(w_in_0_79), .w_in_0_80(w_in_0_80), .w_in_0_81(w_in_0_81), .w_in_0_82(w_in_0_82), .w_in_0_83(w_in_0_83), .w_in_0_84(w_in_0_84), .w_in_0_85(w_in_0_85), .w_in_0_86(w_in_0_86), .w_in_0_87(w_in_0_87), .w_in_0_88(w_in_0_88), .w_in_0_89(w_in_0_89), .w_in_0_90(w_in_0_90), .w_in_0_91(w_in_0_91), .w_in_0_92(w_in_0_92), .w_in_0_93(w_in_0_93), .w_in_0_94(w_in_0_94), .w_in_0_95(w_in_0_95), .w_in_0_96(w_in_0_96), .w_in_0_97(w_in_0_97), .w_in_0_98(w_in_0_98), .w_in_0_99(w_in_0_99), .w_in_0_100(w_in_0_100), .w_in_0_101(w_in_0_101), .w_in_0_102(w_in_0_102), .w_in_0_103(w_in_0_103), .w_in_0_104(w_in_0_104), .w_in_0_105(w_in_0_105), .w_in_0_106(w_in_0_106), .w_in_0_107(w_in_0_107), .w_in_0_108(w_in_0_108), .w_in_0_109(w_in_0_109), .w_in_0_110(w_in_0_110), .w_in_0_111(w_in_0_111), .w_in_0_112(w_in_0_112), .w_in_0_113(w_in_0_113), .w_in_0_114(w_in_0_114), .w_in_0_115(w_in_0_115), .w_in_0_116(w_in_0_116), .w_in_0_117(w_in_0_117), .w_in_0_118(w_in_0_118), .w_in_0_119(w_in_0_119), .w_in_0_120(w_in_0_120), .w_in_0_121(w_in_0_121), .w_in_0_122(w_in_0_122), .w_in_0_123(w_in_0_123), .w_in_0_124(w_in_0_124), .w_in_0_125(w_in_0_125), .w_in_0_126(w_in_0_126), .w_in_0_127(w_in_0_127), .w_in_0_128(w_in_0_128), .w_in_0_129(w_in_0_129), .w_in_0_130(w_in_0_130), .w_in_0_131(w_in_0_131), .w_in_0_132(w_in_0_132), .w_in_0_133(w_in_0_133), .w_in_0_134(w_in_0_134), .w_in_0_135(w_in_0_135), .w_in_0_136(w_in_0_136), .w_in_0_137(w_in_0_137), .w_in_0_138(w_in_0_138), .w_in_0_139(w_in_0_139), .w_in_0_140(w_in_0_140), .w_in_0_141(w_in_0_141), .w_in_0_142(w_in_0_142), .w_in_0_143(w_in_0_143), .w_in_0_144(w_in_0_144), .w_in_0_145(w_in_0_145), .w_in_0_146(w_in_0_146), .w_in_0_147(w_in_0_147), .w_in_0_148(w_in_0_148), .w_in_0_149(w_in_0_149), .w_in_0_150(w_in_0_150), .w_in_0_151(w_in_0_151), .w_in_0_152(w_in_0_152), .w_in_0_153(w_in_0_153), .w_in_0_154(w_in_0_154), .w_in_0_155(w_in_0_155), .w_in_0_156(w_in_0_156), .w_in_0_157(w_in_0_157), .w_in_0_158(w_in_0_158), .w_in_0_159(w_in_0_159), .w_in_0_160(w_in_0_160), .w_in_0_161(w_in_0_161), .w_in_0_162(w_in_0_162), .w_in_0_163(w_in_0_163), .w_in_0_164(w_in_0_164), .w_in_0_165(w_in_0_165), .w_in_0_166(w_in_0_166), .w_in_0_167(w_in_0_167), .w_in_0_168(w_in_0_168), .w_in_0_169(w_in_0_169), .w_in_0_170(w_in_0_170), .w_in_0_171(w_in_0_171), .w_in_0_172(w_in_0_172), .w_in_0_173(w_in_0_173), .w_in_0_174(w_in_0_174), .w_in_0_175(w_in_0_175), .w_in_0_176(w_in_0_176), .w_in_0_177(w_in_0_177), .w_in_0_178(w_in_0_178), .w_in_0_179(w_in_0_179), .w_in_0_180(w_in_0_180), .w_in_0_181(w_in_0_181), .w_in_0_182(w_in_0_182), .w_in_0_183(w_in_0_183), .w_in_0_184(w_in_0_184), .w_in_0_185(w_in_0_185), .w_in_0_186(w_in_0_186), .w_in_0_187(w_in_0_187), .w_in_0_188(w_in_0_188), .w_in_0_189(w_in_0_189), .w_in_0_190(w_in_0_190), .w_in_0_191(w_in_0_191), .w_in_0_192(w_in_0_192), .w_in_0_193(w_in_0_193), .w_in_0_194(w_in_0_194), .w_in_0_195(w_in_0_195), .w_in_0_196(w_in_0_196), .w_in_0_197(w_in_0_197), .w_in_0_198(w_in_0_198), .w_in_0_199(w_in_0_199), .w_in_0_200(w_in_0_200), .w_in_0_201(w_in_0_201), .w_in_0_202(w_in_0_202), .w_in_0_203(w_in_0_203), .w_in_0_204(w_in_0_204), .w_in_0_205(w_in_0_205), .w_in_0_206(w_in_0_206), .w_in_0_207(w_in_0_207), .w_in_0_208(w_in_0_208), .w_in_0_209(w_in_0_209), .w_in_0_210(w_in_0_210), .w_in_0_211(w_in_0_211), .w_in_0_212(w_in_0_212), .w_in_0_213(w_in_0_213), .w_in_0_214(w_in_0_214), .w_in_0_215(w_in_0_215), .w_in_0_216(w_in_0_216), .w_in_0_217(w_in_0_217), .w_in_0_218(w_in_0_218), .w_in_0_219(w_in_0_219), .w_in_0_220(w_in_0_220), .w_in_0_221(w_in_0_221), .w_in_0_222(w_in_0_222), .w_in_0_223(w_in_0_223), .w_in_0_224(w_in_0_224), .w_in_0_225(w_in_0_225), .w_in_0_226(w_in_0_226), .w_in_0_227(w_in_0_227), .w_in_0_228(w_in_0_228), .w_in_0_229(w_in_0_229), .w_in_0_230(w_in_0_230), .w_in_0_231(w_in_0_231), .w_in_0_232(w_in_0_232), .w_in_0_233(w_in_0_233), .w_in_0_234(w_in_0_234), .w_in_0_235(w_in_0_235), .w_in_0_236(w_in_0_236), .w_in_0_237(w_in_0_237), .w_in_0_238(w_in_0_238), .w_in_0_239(w_in_0_239), .w_in_0_240(w_in_0_240), .w_in_0_241(w_in_0_241), .w_in_0_242(w_in_0_242), .w_in_0_243(w_in_0_243), .w_in_0_244(w_in_0_244), .w_in_0_245(w_in_0_245), .w_in_0_246(w_in_0_246), .w_in_0_247(w_in_0_247), .w_in_0_248(w_in_0_248), .w_in_0_249(w_in_0_249), .w_in_0_250(w_in_0_250), .w_in_0_251(w_in_0_251), .w_in_0_252(w_in_0_252), .w_in_0_253(w_in_0_253), .w_in_0_254(w_in_0_254), .w_in_0_255(w_in_0_255), .w_in_1_0(w_in_1_0), .w_in_1_1(w_in_1_1), .w_in_1_2(w_in_1_2), .w_in_1_3(w_in_1_3), .w_in_1_4(w_in_1_4), .w_in_1_5(w_in_1_5), .w_in_1_6(w_in_1_6), .w_in_1_7(w_in_1_7), .w_in_1_8(w_in_1_8), .w_in_1_9(w_in_1_9), .w_in_1_10(w_in_1_10), .w_in_1_11(w_in_1_11), .w_in_1_12(w_in_1_12), .w_in_1_13(w_in_1_13), .w_in_1_14(w_in_1_14), .w_in_1_15(w_in_1_15), .w_in_1_16(w_in_1_16), .w_in_1_17(w_in_1_17), .w_in_1_18(w_in_1_18), .w_in_1_19(w_in_1_19), .w_in_1_20(w_in_1_20), .w_in_1_21(w_in_1_21), .w_in_1_22(w_in_1_22), .w_in_1_23(w_in_1_23), .w_in_1_24(w_in_1_24), .w_in_1_25(w_in_1_25), .w_in_1_26(w_in_1_26), .w_in_1_27(w_in_1_27), .w_in_1_28(w_in_1_28), .w_in_1_29(w_in_1_29), .w_in_1_30(w_in_1_30), .w_in_1_31(w_in_1_31), .w_in_1_32(w_in_1_32), .w_in_1_33(w_in_1_33), .w_in_1_34(w_in_1_34), .w_in_1_35(w_in_1_35), .w_in_1_36(w_in_1_36), .w_in_1_37(w_in_1_37), .w_in_1_38(w_in_1_38), .w_in_1_39(w_in_1_39), .w_in_1_40(w_in_1_40), .w_in_1_41(w_in_1_41), .w_in_1_42(w_in_1_42), .w_in_1_43(w_in_1_43), .w_in_1_44(w_in_1_44), .w_in_1_45(w_in_1_45), .w_in_1_46(w_in_1_46), .w_in_1_47(w_in_1_47), .w_in_1_48(w_in_1_48), .w_in_1_49(w_in_1_49), .w_in_1_50(w_in_1_50), .w_in_1_51(w_in_1_51), .w_in_1_52(w_in_1_52), .w_in_1_53(w_in_1_53), .w_in_1_54(w_in_1_54), .w_in_1_55(w_in_1_55), .w_in_1_56(w_in_1_56), .w_in_1_57(w_in_1_57), .w_in_1_58(w_in_1_58), .w_in_1_59(w_in_1_59), .w_in_1_60(w_in_1_60), .w_in_1_61(w_in_1_61), .w_in_1_62(w_in_1_62), .w_in_1_63(w_in_1_63), .w_in_1_64(w_in_1_64), .w_in_1_65(w_in_1_65), .w_in_1_66(w_in_1_66), .w_in_1_67(w_in_1_67), .w_in_1_68(w_in_1_68), .w_in_1_69(w_in_1_69), .w_in_1_70(w_in_1_70), .w_in_1_71(w_in_1_71), .w_in_1_72(w_in_1_72), .w_in_1_73(w_in_1_73), .w_in_1_74(w_in_1_74), .w_in_1_75(w_in_1_75), .w_in_1_76(w_in_1_76), .w_in_1_77(w_in_1_77), .w_in_1_78(w_in_1_78), .w_in_1_79(w_in_1_79), .w_in_1_80(w_in_1_80), .w_in_1_81(w_in_1_81), .w_in_1_82(w_in_1_82), .w_in_1_83(w_in_1_83), .w_in_1_84(w_in_1_84), .w_in_1_85(w_in_1_85), .w_in_1_86(w_in_1_86), .w_in_1_87(w_in_1_87), .w_in_1_88(w_in_1_88), .w_in_1_89(w_in_1_89), .w_in_1_90(w_in_1_90), .w_in_1_91(w_in_1_91), .w_in_1_92(w_in_1_92), .w_in_1_93(w_in_1_93), .w_in_1_94(w_in_1_94), .w_in_1_95(w_in_1_95), .w_in_1_96(w_in_1_96), .w_in_1_97(w_in_1_97), .w_in_1_98(w_in_1_98), .w_in_1_99(w_in_1_99), .w_in_1_100(w_in_1_100), .w_in_1_101(w_in_1_101), .w_in_1_102(w_in_1_102), .w_in_1_103(w_in_1_103), .w_in_1_104(w_in_1_104), .w_in_1_105(w_in_1_105), .w_in_1_106(w_in_1_106), .w_in_1_107(w_in_1_107), .w_in_1_108(w_in_1_108), .w_in_1_109(w_in_1_109), .w_in_1_110(w_in_1_110), .w_in_1_111(w_in_1_111), .w_in_1_112(w_in_1_112), .w_in_1_113(w_in_1_113), .w_in_1_114(w_in_1_114), .w_in_1_115(w_in_1_115), .w_in_1_116(w_in_1_116), .w_in_1_117(w_in_1_117), .w_in_1_118(w_in_1_118), .w_in_1_119(w_in_1_119), .w_in_1_120(w_in_1_120), .w_in_1_121(w_in_1_121), .w_in_1_122(w_in_1_122), .w_in_1_123(w_in_1_123), .w_in_1_124(w_in_1_124), .w_in_1_125(w_in_1_125), .w_in_1_126(w_in_1_126), .w_in_1_127(w_in_1_127), .w_in_1_128(w_in_1_128), .w_in_1_129(w_in_1_129), .w_in_1_130(w_in_1_130), .w_in_1_131(w_in_1_131), .w_in_1_132(w_in_1_132), .w_in_1_133(w_in_1_133), .w_in_1_134(w_in_1_134), .w_in_1_135(w_in_1_135), .w_in_1_136(w_in_1_136), .w_in_1_137(w_in_1_137), .w_in_1_138(w_in_1_138), .w_in_1_139(w_in_1_139), .w_in_1_140(w_in_1_140), .w_in_1_141(w_in_1_141), .w_in_1_142(w_in_1_142), .w_in_1_143(w_in_1_143), .w_in_1_144(w_in_1_144), .w_in_1_145(w_in_1_145), .w_in_1_146(w_in_1_146), .w_in_1_147(w_in_1_147), .w_in_1_148(w_in_1_148), .w_in_1_149(w_in_1_149), .w_in_1_150(w_in_1_150), .w_in_1_151(w_in_1_151), .w_in_1_152(w_in_1_152), .w_in_1_153(w_in_1_153), .w_in_1_154(w_in_1_154), .w_in_1_155(w_in_1_155), .w_in_1_156(w_in_1_156), .w_in_1_157(w_in_1_157), .w_in_1_158(w_in_1_158), .w_in_1_159(w_in_1_159), .w_in_1_160(w_in_1_160), .w_in_1_161(w_in_1_161), .w_in_1_162(w_in_1_162), .w_in_1_163(w_in_1_163), .w_in_1_164(w_in_1_164), .w_in_1_165(w_in_1_165), .w_in_1_166(w_in_1_166), .w_in_1_167(w_in_1_167), .w_in_1_168(w_in_1_168), .w_in_1_169(w_in_1_169), .w_in_1_170(w_in_1_170), .w_in_1_171(w_in_1_171), .w_in_1_172(w_in_1_172), .w_in_1_173(w_in_1_173), .w_in_1_174(w_in_1_174), .w_in_1_175(w_in_1_175), .w_in_1_176(w_in_1_176), .w_in_1_177(w_in_1_177), .w_in_1_178(w_in_1_178), .w_in_1_179(w_in_1_179), .w_in_1_180(w_in_1_180), .w_in_1_181(w_in_1_181), .w_in_1_182(w_in_1_182), .w_in_1_183(w_in_1_183), .w_in_1_184(w_in_1_184), .w_in_1_185(w_in_1_185), .w_in_1_186(w_in_1_186), .w_in_1_187(w_in_1_187), .w_in_1_188(w_in_1_188), .w_in_1_189(w_in_1_189), .w_in_1_190(w_in_1_190), .w_in_1_191(w_in_1_191), .w_in_1_192(w_in_1_192), .w_in_1_193(w_in_1_193), .w_in_1_194(w_in_1_194), .w_in_1_195(w_in_1_195), .w_in_1_196(w_in_1_196), .w_in_1_197(w_in_1_197), .w_in_1_198(w_in_1_198), .w_in_1_199(w_in_1_199), .w_in_1_200(w_in_1_200), .w_in_1_201(w_in_1_201), .w_in_1_202(w_in_1_202), .w_in_1_203(w_in_1_203), .w_in_1_204(w_in_1_204), .w_in_1_205(w_in_1_205), .w_in_1_206(w_in_1_206), .w_in_1_207(w_in_1_207), .w_in_1_208(w_in_1_208), .w_in_1_209(w_in_1_209), .w_in_1_210(w_in_1_210), .w_in_1_211(w_in_1_211), .w_in_1_212(w_in_1_212), .w_in_1_213(w_in_1_213), .w_in_1_214(w_in_1_214), .w_in_1_215(w_in_1_215), .w_in_1_216(w_in_1_216), .w_in_1_217(w_in_1_217), .w_in_1_218(w_in_1_218), .w_in_1_219(w_in_1_219), .w_in_1_220(w_in_1_220), .w_in_1_221(w_in_1_221), .w_in_1_222(w_in_1_222), .w_in_1_223(w_in_1_223), .w_in_1_224(w_in_1_224), .w_in_1_225(w_in_1_225), .w_in_1_226(w_in_1_226), .w_in_1_227(w_in_1_227), .w_in_1_228(w_in_1_228), .w_in_1_229(w_in_1_229), .w_in_1_230(w_in_1_230), .w_in_1_231(w_in_1_231), .w_in_1_232(w_in_1_232), .w_in_1_233(w_in_1_233), .w_in_1_234(w_in_1_234), .w_in_1_235(w_in_1_235), .w_in_1_236(w_in_1_236), .w_in_1_237(w_in_1_237), .w_in_1_238(w_in_1_238), .w_in_1_239(w_in_1_239), .w_in_1_240(w_in_1_240), .w_in_1_241(w_in_1_241), .w_in_1_242(w_in_1_242), .w_in_1_243(w_in_1_243), .w_in_1_244(w_in_1_244), .w_in_1_245(w_in_1_245), .w_in_1_246(w_in_1_246), .w_in_1_247(w_in_1_247), .w_in_1_248(w_in_1_248), .w_in_1_249(w_in_1_249), .w_in_1_250(w_in_1_250), .w_in_1_251(w_in_1_251), .w_in_1_252(w_in_1_252), .w_in_1_253(w_in_1_253), .w_in_1_254(w_in_1_254), .w_in_1_255(w_in_1_255), .w_in_2_0(w_in_2_0), .w_in_2_1(w_in_2_1), .w_in_2_2(w_in_2_2), .w_in_2_3(w_in_2_3), .w_in_2_4(w_in_2_4), .w_in_2_5(w_in_2_5), .w_in_2_6(w_in_2_6), .w_in_2_7(w_in_2_7), .w_in_2_8(w_in_2_8), .w_in_2_9(w_in_2_9), .w_in_2_10(w_in_2_10), .w_in_2_11(w_in_2_11), .w_in_2_12(w_in_2_12), .w_in_2_13(w_in_2_13), .w_in_2_14(w_in_2_14), .w_in_2_15(w_in_2_15), .w_in_2_16(w_in_2_16), .w_in_2_17(w_in_2_17), .w_in_2_18(w_in_2_18), .w_in_2_19(w_in_2_19), .w_in_2_20(w_in_2_20), .w_in_2_21(w_in_2_21), .w_in_2_22(w_in_2_22), .w_in_2_23(w_in_2_23), .w_in_2_24(w_in_2_24), .w_in_2_25(w_in_2_25), .w_in_2_26(w_in_2_26), .w_in_2_27(w_in_2_27), .w_in_2_28(w_in_2_28), .w_in_2_29(w_in_2_29), .w_in_2_30(w_in_2_30), .w_in_2_31(w_in_2_31), .w_in_2_32(w_in_2_32), .w_in_2_33(w_in_2_33), .w_in_2_34(w_in_2_34), .w_in_2_35(w_in_2_35), .w_in_2_36(w_in_2_36), .w_in_2_37(w_in_2_37), .w_in_2_38(w_in_2_38), .w_in_2_39(w_in_2_39), .w_in_2_40(w_in_2_40), .w_in_2_41(w_in_2_41), .w_in_2_42(w_in_2_42), .w_in_2_43(w_in_2_43), .w_in_2_44(w_in_2_44), .w_in_2_45(w_in_2_45), .w_in_2_46(w_in_2_46), .w_in_2_47(w_in_2_47), .w_in_2_48(w_in_2_48), .w_in_2_49(w_in_2_49), .w_in_2_50(w_in_2_50), .w_in_2_51(w_in_2_51), .w_in_2_52(w_in_2_52), .w_in_2_53(w_in_2_53), .w_in_2_54(w_in_2_54), .w_in_2_55(w_in_2_55), .w_in_2_56(w_in_2_56), .w_in_2_57(w_in_2_57), .w_in_2_58(w_in_2_58), .w_in_2_59(w_in_2_59), .w_in_2_60(w_in_2_60), .w_in_2_61(w_in_2_61), .w_in_2_62(w_in_2_62), .w_in_2_63(w_in_2_63), .w_in_2_64(w_in_2_64), .w_in_2_65(w_in_2_65), .w_in_2_66(w_in_2_66), .w_in_2_67(w_in_2_67), .w_in_2_68(w_in_2_68), .w_in_2_69(w_in_2_69), .w_in_2_70(w_in_2_70), .w_in_2_71(w_in_2_71), .w_in_2_72(w_in_2_72), .w_in_2_73(w_in_2_73), .w_in_2_74(w_in_2_74), .w_in_2_75(w_in_2_75), .w_in_2_76(w_in_2_76), .w_in_2_77(w_in_2_77), .w_in_2_78(w_in_2_78), .w_in_2_79(w_in_2_79), .w_in_2_80(w_in_2_80), .w_in_2_81(w_in_2_81), .w_in_2_82(w_in_2_82), .w_in_2_83(w_in_2_83), .w_in_2_84(w_in_2_84), .w_in_2_85(w_in_2_85), .w_in_2_86(w_in_2_86), .w_in_2_87(w_in_2_87), .w_in_2_88(w_in_2_88), .w_in_2_89(w_in_2_89), .w_in_2_90(w_in_2_90), .w_in_2_91(w_in_2_91), .w_in_2_92(w_in_2_92), .w_in_2_93(w_in_2_93), .w_in_2_94(w_in_2_94), .w_in_2_95(w_in_2_95), .w_in_2_96(w_in_2_96), .w_in_2_97(w_in_2_97), .w_in_2_98(w_in_2_98), .w_in_2_99(w_in_2_99), .w_in_2_100(w_in_2_100), .w_in_2_101(w_in_2_101), .w_in_2_102(w_in_2_102), .w_in_2_103(w_in_2_103), .w_in_2_104(w_in_2_104), .w_in_2_105(w_in_2_105), .w_in_2_106(w_in_2_106), .w_in_2_107(w_in_2_107), .w_in_2_108(w_in_2_108), .w_in_2_109(w_in_2_109), .w_in_2_110(w_in_2_110), .w_in_2_111(w_in_2_111), .w_in_2_112(w_in_2_112), .w_in_2_113(w_in_2_113), .w_in_2_114(w_in_2_114), .w_in_2_115(w_in_2_115), .w_in_2_116(w_in_2_116), .w_in_2_117(w_in_2_117), .w_in_2_118(w_in_2_118), .w_in_2_119(w_in_2_119), .w_in_2_120(w_in_2_120), .w_in_2_121(w_in_2_121), .w_in_2_122(w_in_2_122), .w_in_2_123(w_in_2_123), .w_in_2_124(w_in_2_124), .w_in_2_125(w_in_2_125), .w_in_2_126(w_in_2_126), .w_in_2_127(w_in_2_127), .w_in_2_128(w_in_2_128), .w_in_2_129(w_in_2_129), .w_in_2_130(w_in_2_130), .w_in_2_131(w_in_2_131), .w_in_2_132(w_in_2_132), .w_in_2_133(w_in_2_133), .w_in_2_134(w_in_2_134), .w_in_2_135(w_in_2_135), .w_in_2_136(w_in_2_136), .w_in_2_137(w_in_2_137), .w_in_2_138(w_in_2_138), .w_in_2_139(w_in_2_139), .w_in_2_140(w_in_2_140), .w_in_2_141(w_in_2_141), .w_in_2_142(w_in_2_142), .w_in_2_143(w_in_2_143), .w_in_2_144(w_in_2_144), .w_in_2_145(w_in_2_145), .w_in_2_146(w_in_2_146), .w_in_2_147(w_in_2_147), .w_in_2_148(w_in_2_148), .w_in_2_149(w_in_2_149), .w_in_2_150(w_in_2_150), .w_in_2_151(w_in_2_151), .w_in_2_152(w_in_2_152), .w_in_2_153(w_in_2_153), .w_in_2_154(w_in_2_154), .w_in_2_155(w_in_2_155), .w_in_2_156(w_in_2_156), .w_in_2_157(w_in_2_157), .w_in_2_158(w_in_2_158), .w_in_2_159(w_in_2_159), .w_in_2_160(w_in_2_160), .w_in_2_161(w_in_2_161), .w_in_2_162(w_in_2_162), .w_in_2_163(w_in_2_163), .w_in_2_164(w_in_2_164), .w_in_2_165(w_in_2_165), .w_in_2_166(w_in_2_166), .w_in_2_167(w_in_2_167), .w_in_2_168(w_in_2_168), .w_in_2_169(w_in_2_169), .w_in_2_170(w_in_2_170), .w_in_2_171(w_in_2_171), .w_in_2_172(w_in_2_172), .w_in_2_173(w_in_2_173), .w_in_2_174(w_in_2_174), .w_in_2_175(w_in_2_175), .w_in_2_176(w_in_2_176), .w_in_2_177(w_in_2_177), .w_in_2_178(w_in_2_178), .w_in_2_179(w_in_2_179), .w_in_2_180(w_in_2_180), .w_in_2_181(w_in_2_181), .w_in_2_182(w_in_2_182), .w_in_2_183(w_in_2_183), .w_in_2_184(w_in_2_184), .w_in_2_185(w_in_2_185), .w_in_2_186(w_in_2_186), .w_in_2_187(w_in_2_187), .w_in_2_188(w_in_2_188), .w_in_2_189(w_in_2_189), .w_in_2_190(w_in_2_190), .w_in_2_191(w_in_2_191), .w_in_2_192(w_in_2_192), .w_in_2_193(w_in_2_193), .w_in_2_194(w_in_2_194), .w_in_2_195(w_in_2_195), .w_in_2_196(w_in_2_196), .w_in_2_197(w_in_2_197), .w_in_2_198(w_in_2_198), .w_in_2_199(w_in_2_199), .w_in_2_200(w_in_2_200), .w_in_2_201(w_in_2_201), .w_in_2_202(w_in_2_202), .w_in_2_203(w_in_2_203), .w_in_2_204(w_in_2_204), .w_in_2_205(w_in_2_205), .w_in_2_206(w_in_2_206), .w_in_2_207(w_in_2_207), .w_in_2_208(w_in_2_208), .w_in_2_209(w_in_2_209), .w_in_2_210(w_in_2_210), .w_in_2_211(w_in_2_211), .w_in_2_212(w_in_2_212), .w_in_2_213(w_in_2_213), .w_in_2_214(w_in_2_214), .w_in_2_215(w_in_2_215), .w_in_2_216(w_in_2_216), .w_in_2_217(w_in_2_217), .w_in_2_218(w_in_2_218), .w_in_2_219(w_in_2_219), .w_in_2_220(w_in_2_220), .w_in_2_221(w_in_2_221), .w_in_2_222(w_in_2_222), .w_in_2_223(w_in_2_223), .w_in_2_224(w_in_2_224), .w_in_2_225(w_in_2_225), .w_in_2_226(w_in_2_226), .w_in_2_227(w_in_2_227), .w_in_2_228(w_in_2_228), .w_in_2_229(w_in_2_229), .w_in_2_230(w_in_2_230), .w_in_2_231(w_in_2_231), .w_in_2_232(w_in_2_232), .w_in_2_233(w_in_2_233), .w_in_2_234(w_in_2_234), .w_in_2_235(w_in_2_235), .w_in_2_236(w_in_2_236), .w_in_2_237(w_in_2_237), .w_in_2_238(w_in_2_238), .w_in_2_239(w_in_2_239), .w_in_2_240(w_in_2_240), .w_in_2_241(w_in_2_241), .w_in_2_242(w_in_2_242), .w_in_2_243(w_in_2_243), .w_in_2_244(w_in_2_244), .w_in_2_245(w_in_2_245), .w_in_2_246(w_in_2_246), .w_in_2_247(w_in_2_247), .w_in_2_248(w_in_2_248), .w_in_2_249(w_in_2_249), .w_in_2_250(w_in_2_250), .w_in_2_251(w_in_2_251), .w_in_2_252(w_in_2_252), .w_in_2_253(w_in_2_253), .w_in_2_254(w_in_2_254), .w_in_2_255(w_in_2_255), .w_in_3_0(w_in_3_0), .w_in_3_1(w_in_3_1), .w_in_3_2(w_in_3_2), .w_in_3_3(w_in_3_3), .w_in_3_4(w_in_3_4), .w_in_3_5(w_in_3_5), .w_in_3_6(w_in_3_6), .w_in_3_7(w_in_3_7), .w_in_3_8(w_in_3_8), .w_in_3_9(w_in_3_9), .w_in_3_10(w_in_3_10), .w_in_3_11(w_in_3_11), .w_in_3_12(w_in_3_12), .w_in_3_13(w_in_3_13), .w_in_3_14(w_in_3_14), .w_in_3_15(w_in_3_15), .w_in_3_16(w_in_3_16), .w_in_3_17(w_in_3_17), .w_in_3_18(w_in_3_18), .w_in_3_19(w_in_3_19), .w_in_3_20(w_in_3_20), .w_in_3_21(w_in_3_21), .w_in_3_22(w_in_3_22), .w_in_3_23(w_in_3_23), .w_in_3_24(w_in_3_24), .w_in_3_25(w_in_3_25), .w_in_3_26(w_in_3_26), .w_in_3_27(w_in_3_27), .w_in_3_28(w_in_3_28), .w_in_3_29(w_in_3_29), .w_in_3_30(w_in_3_30), .w_in_3_31(w_in_3_31), .w_in_3_32(w_in_3_32), .w_in_3_33(w_in_3_33), .w_in_3_34(w_in_3_34), .w_in_3_35(w_in_3_35), .w_in_3_36(w_in_3_36), .w_in_3_37(w_in_3_37), .w_in_3_38(w_in_3_38), .w_in_3_39(w_in_3_39), .w_in_3_40(w_in_3_40), .w_in_3_41(w_in_3_41), .w_in_3_42(w_in_3_42), .w_in_3_43(w_in_3_43), .w_in_3_44(w_in_3_44), .w_in_3_45(w_in_3_45), .w_in_3_46(w_in_3_46), .w_in_3_47(w_in_3_47), .w_in_3_48(w_in_3_48), .w_in_3_49(w_in_3_49), .w_in_3_50(w_in_3_50), .w_in_3_51(w_in_3_51), .w_in_3_52(w_in_3_52), .w_in_3_53(w_in_3_53), .w_in_3_54(w_in_3_54), .w_in_3_55(w_in_3_55), .w_in_3_56(w_in_3_56), .w_in_3_57(w_in_3_57), .w_in_3_58(w_in_3_58), .w_in_3_59(w_in_3_59), .w_in_3_60(w_in_3_60), .w_in_3_61(w_in_3_61), .w_in_3_62(w_in_3_62), .w_in_3_63(w_in_3_63), .w_in_3_64(w_in_3_64), .w_in_3_65(w_in_3_65), .w_in_3_66(w_in_3_66), .w_in_3_67(w_in_3_67), .w_in_3_68(w_in_3_68), .w_in_3_69(w_in_3_69), .w_in_3_70(w_in_3_70), .w_in_3_71(w_in_3_71), .w_in_3_72(w_in_3_72), .w_in_3_73(w_in_3_73), .w_in_3_74(w_in_3_74), .w_in_3_75(w_in_3_75), .w_in_3_76(w_in_3_76), .w_in_3_77(w_in_3_77), .w_in_3_78(w_in_3_78), .w_in_3_79(w_in_3_79), .w_in_3_80(w_in_3_80), .w_in_3_81(w_in_3_81), .w_in_3_82(w_in_3_82), .w_in_3_83(w_in_3_83), .w_in_3_84(w_in_3_84), .w_in_3_85(w_in_3_85), .w_in_3_86(w_in_3_86), .w_in_3_87(w_in_3_87), .w_in_3_88(w_in_3_88), .w_in_3_89(w_in_3_89), .w_in_3_90(w_in_3_90), .w_in_3_91(w_in_3_91), .w_in_3_92(w_in_3_92), .w_in_3_93(w_in_3_93), .w_in_3_94(w_in_3_94), .w_in_3_95(w_in_3_95), .w_in_3_96(w_in_3_96), .w_in_3_97(w_in_3_97), .w_in_3_98(w_in_3_98), .w_in_3_99(w_in_3_99), .w_in_3_100(w_in_3_100), .w_in_3_101(w_in_3_101), .w_in_3_102(w_in_3_102), .w_in_3_103(w_in_3_103), .w_in_3_104(w_in_3_104), .w_in_3_105(w_in_3_105), .w_in_3_106(w_in_3_106), .w_in_3_107(w_in_3_107), .w_in_3_108(w_in_3_108), .w_in_3_109(w_in_3_109), .w_in_3_110(w_in_3_110), .w_in_3_111(w_in_3_111), .w_in_3_112(w_in_3_112), .w_in_3_113(w_in_3_113), .w_in_3_114(w_in_3_114), .w_in_3_115(w_in_3_115), .w_in_3_116(w_in_3_116), .w_in_3_117(w_in_3_117), .w_in_3_118(w_in_3_118), .w_in_3_119(w_in_3_119), .w_in_3_120(w_in_3_120), .w_in_3_121(w_in_3_121), .w_in_3_122(w_in_3_122), .w_in_3_123(w_in_3_123), .w_in_3_124(w_in_3_124), .w_in_3_125(w_in_3_125), .w_in_3_126(w_in_3_126), .w_in_3_127(w_in_3_127), .w_in_3_128(w_in_3_128), .w_in_3_129(w_in_3_129), .w_in_3_130(w_in_3_130), .w_in_3_131(w_in_3_131), .w_in_3_132(w_in_3_132), .w_in_3_133(w_in_3_133), .w_in_3_134(w_in_3_134), .w_in_3_135(w_in_3_135), .w_in_3_136(w_in_3_136), .w_in_3_137(w_in_3_137), .w_in_3_138(w_in_3_138), .w_in_3_139(w_in_3_139), .w_in_3_140(w_in_3_140), .w_in_3_141(w_in_3_141), .w_in_3_142(w_in_3_142), .w_in_3_143(w_in_3_143), .w_in_3_144(w_in_3_144), .w_in_3_145(w_in_3_145), .w_in_3_146(w_in_3_146), .w_in_3_147(w_in_3_147), .w_in_3_148(w_in_3_148), .w_in_3_149(w_in_3_149), .w_in_3_150(w_in_3_150), .w_in_3_151(w_in_3_151), .w_in_3_152(w_in_3_152), .w_in_3_153(w_in_3_153), .w_in_3_154(w_in_3_154), .w_in_3_155(w_in_3_155), .w_in_3_156(w_in_3_156), .w_in_3_157(w_in_3_157), .w_in_3_158(w_in_3_158), .w_in_3_159(w_in_3_159), .w_in_3_160(w_in_3_160), .w_in_3_161(w_in_3_161), .w_in_3_162(w_in_3_162), .w_in_3_163(w_in_3_163), .w_in_3_164(w_in_3_164), .w_in_3_165(w_in_3_165), .w_in_3_166(w_in_3_166), .w_in_3_167(w_in_3_167), .w_in_3_168(w_in_3_168), .w_in_3_169(w_in_3_169), .w_in_3_170(w_in_3_170), .w_in_3_171(w_in_3_171), .w_in_3_172(w_in_3_172), .w_in_3_173(w_in_3_173), .w_in_3_174(w_in_3_174), .w_in_3_175(w_in_3_175), .w_in_3_176(w_in_3_176), .w_in_3_177(w_in_3_177), .w_in_3_178(w_in_3_178), .w_in_3_179(w_in_3_179), .w_in_3_180(w_in_3_180), .w_in_3_181(w_in_3_181), .w_in_3_182(w_in_3_182), .w_in_3_183(w_in_3_183), .w_in_3_184(w_in_3_184), .w_in_3_185(w_in_3_185), .w_in_3_186(w_in_3_186), .w_in_3_187(w_in_3_187), .w_in_3_188(w_in_3_188), .w_in_3_189(w_in_3_189), .w_in_3_190(w_in_3_190), .w_in_3_191(w_in_3_191), .w_in_3_192(w_in_3_192), .w_in_3_193(w_in_3_193), .w_in_3_194(w_in_3_194), .w_in_3_195(w_in_3_195), .w_in_3_196(w_in_3_196), .w_in_3_197(w_in_3_197), .w_in_3_198(w_in_3_198), .w_in_3_199(w_in_3_199), .w_in_3_200(w_in_3_200), .w_in_3_201(w_in_3_201), .w_in_3_202(w_in_3_202), .w_in_3_203(w_in_3_203), .w_in_3_204(w_in_3_204), .w_in_3_205(w_in_3_205), .w_in_3_206(w_in_3_206), .w_in_3_207(w_in_3_207), .w_in_3_208(w_in_3_208), .w_in_3_209(w_in_3_209), .w_in_3_210(w_in_3_210), .w_in_3_211(w_in_3_211), .w_in_3_212(w_in_3_212), .w_in_3_213(w_in_3_213), .w_in_3_214(w_in_3_214), .w_in_3_215(w_in_3_215), .w_in_3_216(w_in_3_216), .w_in_3_217(w_in_3_217), .w_in_3_218(w_in_3_218), .w_in_3_219(w_in_3_219), .w_in_3_220(w_in_3_220), .w_in_3_221(w_in_3_221), .w_in_3_222(w_in_3_222), .w_in_3_223(w_in_3_223), .w_in_3_224(w_in_3_224), .w_in_3_225(w_in_3_225), .w_in_3_226(w_in_3_226), .w_in_3_227(w_in_3_227), .w_in_3_228(w_in_3_228), .w_in_3_229(w_in_3_229), .w_in_3_230(w_in_3_230), .w_in_3_231(w_in_3_231), .w_in_3_232(w_in_3_232), .w_in_3_233(w_in_3_233), .w_in_3_234(w_in_3_234), .w_in_3_235(w_in_3_235), .w_in_3_236(w_in_3_236), .w_in_3_237(w_in_3_237), .w_in_3_238(w_in_3_238), .w_in_3_239(w_in_3_239), .w_in_3_240(w_in_3_240), .w_in_3_241(w_in_3_241), .w_in_3_242(w_in_3_242), .w_in_3_243(w_in_3_243), .w_in_3_244(w_in_3_244), .w_in_3_245(w_in_3_245), .w_in_3_246(w_in_3_246), .w_in_3_247(w_in_3_247), .w_in_3_248(w_in_3_248), .w_in_3_249(w_in_3_249), .w_in_3_250(w_in_3_250), .w_in_3_251(w_in_3_251), .w_in_3_252(w_in_3_252), .w_in_3_253(w_in_3_253), .w_in_3_254(w_in_3_254), .w_in_3_255(w_in_3_255), .w_in_4_0(w_in_4_0), .w_in_4_1(w_in_4_1), .w_in_4_2(w_in_4_2), .w_in_4_3(w_in_4_3), .w_in_4_4(w_in_4_4), .w_in_4_5(w_in_4_5), .w_in_4_6(w_in_4_6), .w_in_4_7(w_in_4_7), .w_in_4_8(w_in_4_8), .w_in_4_9(w_in_4_9), .w_in_4_10(w_in_4_10), .w_in_4_11(w_in_4_11), .w_in_4_12(w_in_4_12), .w_in_4_13(w_in_4_13), .w_in_4_14(w_in_4_14), .w_in_4_15(w_in_4_15), .w_in_4_16(w_in_4_16), .w_in_4_17(w_in_4_17), .w_in_4_18(w_in_4_18), .w_in_4_19(w_in_4_19), .w_in_4_20(w_in_4_20), .w_in_4_21(w_in_4_21), .w_in_4_22(w_in_4_22), .w_in_4_23(w_in_4_23), .w_in_4_24(w_in_4_24), .w_in_4_25(w_in_4_25), .w_in_4_26(w_in_4_26), .w_in_4_27(w_in_4_27), .w_in_4_28(w_in_4_28), .w_in_4_29(w_in_4_29), .w_in_4_30(w_in_4_30), .w_in_4_31(w_in_4_31), .w_in_4_32(w_in_4_32), .w_in_4_33(w_in_4_33), .w_in_4_34(w_in_4_34), .w_in_4_35(w_in_4_35), .w_in_4_36(w_in_4_36), .w_in_4_37(w_in_4_37), .w_in_4_38(w_in_4_38), .w_in_4_39(w_in_4_39), .w_in_4_40(w_in_4_40), .w_in_4_41(w_in_4_41), .w_in_4_42(w_in_4_42), .w_in_4_43(w_in_4_43), .w_in_4_44(w_in_4_44), .w_in_4_45(w_in_4_45), .w_in_4_46(w_in_4_46), .w_in_4_47(w_in_4_47), .w_in_4_48(w_in_4_48), .w_in_4_49(w_in_4_49), .w_in_4_50(w_in_4_50), .w_in_4_51(w_in_4_51), .w_in_4_52(w_in_4_52), .w_in_4_53(w_in_4_53), .w_in_4_54(w_in_4_54), .w_in_4_55(w_in_4_55), .w_in_4_56(w_in_4_56), .w_in_4_57(w_in_4_57), .w_in_4_58(w_in_4_58), .w_in_4_59(w_in_4_59), .w_in_4_60(w_in_4_60), .w_in_4_61(w_in_4_61), .w_in_4_62(w_in_4_62), .w_in_4_63(w_in_4_63), .w_in_4_64(w_in_4_64), .w_in_4_65(w_in_4_65), .w_in_4_66(w_in_4_66), .w_in_4_67(w_in_4_67), .w_in_4_68(w_in_4_68), .w_in_4_69(w_in_4_69), .w_in_4_70(w_in_4_70), .w_in_4_71(w_in_4_71), .w_in_4_72(w_in_4_72), .w_in_4_73(w_in_4_73), .w_in_4_74(w_in_4_74), .w_in_4_75(w_in_4_75), .w_in_4_76(w_in_4_76), .w_in_4_77(w_in_4_77), .w_in_4_78(w_in_4_78), .w_in_4_79(w_in_4_79), .w_in_4_80(w_in_4_80), .w_in_4_81(w_in_4_81), .w_in_4_82(w_in_4_82), .w_in_4_83(w_in_4_83), .w_in_4_84(w_in_4_84), .w_in_4_85(w_in_4_85), .w_in_4_86(w_in_4_86), .w_in_4_87(w_in_4_87), .w_in_4_88(w_in_4_88), .w_in_4_89(w_in_4_89), .w_in_4_90(w_in_4_90), .w_in_4_91(w_in_4_91), .w_in_4_92(w_in_4_92), .w_in_4_93(w_in_4_93), .w_in_4_94(w_in_4_94), .w_in_4_95(w_in_4_95), .w_in_4_96(w_in_4_96), .w_in_4_97(w_in_4_97), .w_in_4_98(w_in_4_98), .w_in_4_99(w_in_4_99), .w_in_4_100(w_in_4_100), .w_in_4_101(w_in_4_101), .w_in_4_102(w_in_4_102), .w_in_4_103(w_in_4_103), .w_in_4_104(w_in_4_104), .w_in_4_105(w_in_4_105), .w_in_4_106(w_in_4_106), .w_in_4_107(w_in_4_107), .w_in_4_108(w_in_4_108), .w_in_4_109(w_in_4_109), .w_in_4_110(w_in_4_110), .w_in_4_111(w_in_4_111), .w_in_4_112(w_in_4_112), .w_in_4_113(w_in_4_113), .w_in_4_114(w_in_4_114), .w_in_4_115(w_in_4_115), .w_in_4_116(w_in_4_116), .w_in_4_117(w_in_4_117), .w_in_4_118(w_in_4_118), .w_in_4_119(w_in_4_119), .w_in_4_120(w_in_4_120), .w_in_4_121(w_in_4_121), .w_in_4_122(w_in_4_122), .w_in_4_123(w_in_4_123), .w_in_4_124(w_in_4_124), .w_in_4_125(w_in_4_125), .w_in_4_126(w_in_4_126), .w_in_4_127(w_in_4_127), .w_in_4_128(w_in_4_128), .w_in_4_129(w_in_4_129), .w_in_4_130(w_in_4_130), .w_in_4_131(w_in_4_131), .w_in_4_132(w_in_4_132), .w_in_4_133(w_in_4_133), .w_in_4_134(w_in_4_134), .w_in_4_135(w_in_4_135), .w_in_4_136(w_in_4_136), .w_in_4_137(w_in_4_137), .w_in_4_138(w_in_4_138), .w_in_4_139(w_in_4_139), .w_in_4_140(w_in_4_140), .w_in_4_141(w_in_4_141), .w_in_4_142(w_in_4_142), .w_in_4_143(w_in_4_143), .w_in_4_144(w_in_4_144), .w_in_4_145(w_in_4_145), .w_in_4_146(w_in_4_146), .w_in_4_147(w_in_4_147), .w_in_4_148(w_in_4_148), .w_in_4_149(w_in_4_149), .w_in_4_150(w_in_4_150), .w_in_4_151(w_in_4_151), .w_in_4_152(w_in_4_152), .w_in_4_153(w_in_4_153), .w_in_4_154(w_in_4_154), .w_in_4_155(w_in_4_155), .w_in_4_156(w_in_4_156), .w_in_4_157(w_in_4_157), .w_in_4_158(w_in_4_158), .w_in_4_159(w_in_4_159), .w_in_4_160(w_in_4_160), .w_in_4_161(w_in_4_161), .w_in_4_162(w_in_4_162), .w_in_4_163(w_in_4_163), .w_in_4_164(w_in_4_164), .w_in_4_165(w_in_4_165), .w_in_4_166(w_in_4_166), .w_in_4_167(w_in_4_167), .w_in_4_168(w_in_4_168), .w_in_4_169(w_in_4_169), .w_in_4_170(w_in_4_170), .w_in_4_171(w_in_4_171), .w_in_4_172(w_in_4_172), .w_in_4_173(w_in_4_173), .w_in_4_174(w_in_4_174), .w_in_4_175(w_in_4_175), .w_in_4_176(w_in_4_176), .w_in_4_177(w_in_4_177), .w_in_4_178(w_in_4_178), .w_in_4_179(w_in_4_179), .w_in_4_180(w_in_4_180), .w_in_4_181(w_in_4_181), .w_in_4_182(w_in_4_182), .w_in_4_183(w_in_4_183), .w_in_4_184(w_in_4_184), .w_in_4_185(w_in_4_185), .w_in_4_186(w_in_4_186), .w_in_4_187(w_in_4_187), .w_in_4_188(w_in_4_188), .w_in_4_189(w_in_4_189), .w_in_4_190(w_in_4_190), .w_in_4_191(w_in_4_191), .w_in_4_192(w_in_4_192), .w_in_4_193(w_in_4_193), .w_in_4_194(w_in_4_194), .w_in_4_195(w_in_4_195), .w_in_4_196(w_in_4_196), .w_in_4_197(w_in_4_197), .w_in_4_198(w_in_4_198), .w_in_4_199(w_in_4_199), .w_in_4_200(w_in_4_200), .w_in_4_201(w_in_4_201), .w_in_4_202(w_in_4_202), .w_in_4_203(w_in_4_203), .w_in_4_204(w_in_4_204), .w_in_4_205(w_in_4_205), .w_in_4_206(w_in_4_206), .w_in_4_207(w_in_4_207), .w_in_4_208(w_in_4_208), .w_in_4_209(w_in_4_209), .w_in_4_210(w_in_4_210), .w_in_4_211(w_in_4_211), .w_in_4_212(w_in_4_212), .w_in_4_213(w_in_4_213), .w_in_4_214(w_in_4_214), .w_in_4_215(w_in_4_215), .w_in_4_216(w_in_4_216), .w_in_4_217(w_in_4_217), .w_in_4_218(w_in_4_218), .w_in_4_219(w_in_4_219), .w_in_4_220(w_in_4_220), .w_in_4_221(w_in_4_221), .w_in_4_222(w_in_4_222), .w_in_4_223(w_in_4_223), .w_in_4_224(w_in_4_224), .w_in_4_225(w_in_4_225), .w_in_4_226(w_in_4_226), .w_in_4_227(w_in_4_227), .w_in_4_228(w_in_4_228), .w_in_4_229(w_in_4_229), .w_in_4_230(w_in_4_230), .w_in_4_231(w_in_4_231), .w_in_4_232(w_in_4_232), .w_in_4_233(w_in_4_233), .w_in_4_234(w_in_4_234), .w_in_4_235(w_in_4_235), .w_in_4_236(w_in_4_236), .w_in_4_237(w_in_4_237), .w_in_4_238(w_in_4_238), .w_in_4_239(w_in_4_239), .w_in_4_240(w_in_4_240), .w_in_4_241(w_in_4_241), .w_in_4_242(w_in_4_242), .w_in_4_243(w_in_4_243), .w_in_4_244(w_in_4_244), .w_in_4_245(w_in_4_245), .w_in_4_246(w_in_4_246), .w_in_4_247(w_in_4_247), .w_in_4_248(w_in_4_248), .w_in_4_249(w_in_4_249), .w_in_4_250(w_in_4_250), .w_in_4_251(w_in_4_251), .w_in_4_252(w_in_4_252), .w_in_4_253(w_in_4_253), .w_in_4_254(w_in_4_254), .w_in_4_255(w_in_4_255), .w_in_5_0(w_in_5_0), .w_in_5_1(w_in_5_1), .w_in_5_2(w_in_5_2), .w_in_5_3(w_in_5_3), .w_in_5_4(w_in_5_4), .w_in_5_5(w_in_5_5), .w_in_5_6(w_in_5_6), .w_in_5_7(w_in_5_7), .w_in_5_8(w_in_5_8), .w_in_5_9(w_in_5_9), .w_in_5_10(w_in_5_10), .w_in_5_11(w_in_5_11), .w_in_5_12(w_in_5_12), .w_in_5_13(w_in_5_13), .w_in_5_14(w_in_5_14), .w_in_5_15(w_in_5_15), .w_in_5_16(w_in_5_16), .w_in_5_17(w_in_5_17), .w_in_5_18(w_in_5_18), .w_in_5_19(w_in_5_19), .w_in_5_20(w_in_5_20), .w_in_5_21(w_in_5_21), .w_in_5_22(w_in_5_22), .w_in_5_23(w_in_5_23), .w_in_5_24(w_in_5_24), .w_in_5_25(w_in_5_25), .w_in_5_26(w_in_5_26), .w_in_5_27(w_in_5_27), .w_in_5_28(w_in_5_28), .w_in_5_29(w_in_5_29), .w_in_5_30(w_in_5_30), .w_in_5_31(w_in_5_31), .w_in_5_32(w_in_5_32), .w_in_5_33(w_in_5_33), .w_in_5_34(w_in_5_34), .w_in_5_35(w_in_5_35), .w_in_5_36(w_in_5_36), .w_in_5_37(w_in_5_37), .w_in_5_38(w_in_5_38), .w_in_5_39(w_in_5_39), .w_in_5_40(w_in_5_40), .w_in_5_41(w_in_5_41), .w_in_5_42(w_in_5_42), .w_in_5_43(w_in_5_43), .w_in_5_44(w_in_5_44), .w_in_5_45(w_in_5_45), .w_in_5_46(w_in_5_46), .w_in_5_47(w_in_5_47), .w_in_5_48(w_in_5_48), .w_in_5_49(w_in_5_49), .w_in_5_50(w_in_5_50), .w_in_5_51(w_in_5_51), .w_in_5_52(w_in_5_52), .w_in_5_53(w_in_5_53), .w_in_5_54(w_in_5_54), .w_in_5_55(w_in_5_55), .w_in_5_56(w_in_5_56), .w_in_5_57(w_in_5_57), .w_in_5_58(w_in_5_58), .w_in_5_59(w_in_5_59), .w_in_5_60(w_in_5_60), .w_in_5_61(w_in_5_61), .w_in_5_62(w_in_5_62), .w_in_5_63(w_in_5_63), .w_in_5_64(w_in_5_64), .w_in_5_65(w_in_5_65), .w_in_5_66(w_in_5_66), .w_in_5_67(w_in_5_67), .w_in_5_68(w_in_5_68), .w_in_5_69(w_in_5_69), .w_in_5_70(w_in_5_70), .w_in_5_71(w_in_5_71), .w_in_5_72(w_in_5_72), .w_in_5_73(w_in_5_73), .w_in_5_74(w_in_5_74), .w_in_5_75(w_in_5_75), .w_in_5_76(w_in_5_76), .w_in_5_77(w_in_5_77), .w_in_5_78(w_in_5_78), .w_in_5_79(w_in_5_79), .w_in_5_80(w_in_5_80), .w_in_5_81(w_in_5_81), .w_in_5_82(w_in_5_82), .w_in_5_83(w_in_5_83), .w_in_5_84(w_in_5_84), .w_in_5_85(w_in_5_85), .w_in_5_86(w_in_5_86), .w_in_5_87(w_in_5_87), .w_in_5_88(w_in_5_88), .w_in_5_89(w_in_5_89), .w_in_5_90(w_in_5_90), .w_in_5_91(w_in_5_91), .w_in_5_92(w_in_5_92), .w_in_5_93(w_in_5_93), .w_in_5_94(w_in_5_94), .w_in_5_95(w_in_5_95), .w_in_5_96(w_in_5_96), .w_in_5_97(w_in_5_97), .w_in_5_98(w_in_5_98), .w_in_5_99(w_in_5_99), .w_in_5_100(w_in_5_100), .w_in_5_101(w_in_5_101), .w_in_5_102(w_in_5_102), .w_in_5_103(w_in_5_103), .w_in_5_104(w_in_5_104), .w_in_5_105(w_in_5_105), .w_in_5_106(w_in_5_106), .w_in_5_107(w_in_5_107), .w_in_5_108(w_in_5_108), .w_in_5_109(w_in_5_109), .w_in_5_110(w_in_5_110), .w_in_5_111(w_in_5_111), .w_in_5_112(w_in_5_112), .w_in_5_113(w_in_5_113), .w_in_5_114(w_in_5_114), .w_in_5_115(w_in_5_115), .w_in_5_116(w_in_5_116), .w_in_5_117(w_in_5_117), .w_in_5_118(w_in_5_118), .w_in_5_119(w_in_5_119), .w_in_5_120(w_in_5_120), .w_in_5_121(w_in_5_121), .w_in_5_122(w_in_5_122), .w_in_5_123(w_in_5_123), .w_in_5_124(w_in_5_124), .w_in_5_125(w_in_5_125), .w_in_5_126(w_in_5_126), .w_in_5_127(w_in_5_127), .w_in_5_128(w_in_5_128), .w_in_5_129(w_in_5_129), .w_in_5_130(w_in_5_130), .w_in_5_131(w_in_5_131), .w_in_5_132(w_in_5_132), .w_in_5_133(w_in_5_133), .w_in_5_134(w_in_5_134), .w_in_5_135(w_in_5_135), .w_in_5_136(w_in_5_136), .w_in_5_137(w_in_5_137), .w_in_5_138(w_in_5_138), .w_in_5_139(w_in_5_139), .w_in_5_140(w_in_5_140), .w_in_5_141(w_in_5_141), .w_in_5_142(w_in_5_142), .w_in_5_143(w_in_5_143), .w_in_5_144(w_in_5_144), .w_in_5_145(w_in_5_145), .w_in_5_146(w_in_5_146), .w_in_5_147(w_in_5_147), .w_in_5_148(w_in_5_148), .w_in_5_149(w_in_5_149), .w_in_5_150(w_in_5_150), .w_in_5_151(w_in_5_151), .w_in_5_152(w_in_5_152), .w_in_5_153(w_in_5_153), .w_in_5_154(w_in_5_154), .w_in_5_155(w_in_5_155), .w_in_5_156(w_in_5_156), .w_in_5_157(w_in_5_157), .w_in_5_158(w_in_5_158), .w_in_5_159(w_in_5_159), .w_in_5_160(w_in_5_160), .w_in_5_161(w_in_5_161), .w_in_5_162(w_in_5_162), .w_in_5_163(w_in_5_163), .w_in_5_164(w_in_5_164), .w_in_5_165(w_in_5_165), .w_in_5_166(w_in_5_166), .w_in_5_167(w_in_5_167), .w_in_5_168(w_in_5_168), .w_in_5_169(w_in_5_169), .w_in_5_170(w_in_5_170), .w_in_5_171(w_in_5_171), .w_in_5_172(w_in_5_172), .w_in_5_173(w_in_5_173), .w_in_5_174(w_in_5_174), .w_in_5_175(w_in_5_175), .w_in_5_176(w_in_5_176), .w_in_5_177(w_in_5_177), .w_in_5_178(w_in_5_178), .w_in_5_179(w_in_5_179), .w_in_5_180(w_in_5_180), .w_in_5_181(w_in_5_181), .w_in_5_182(w_in_5_182), .w_in_5_183(w_in_5_183), .w_in_5_184(w_in_5_184), .w_in_5_185(w_in_5_185), .w_in_5_186(w_in_5_186), .w_in_5_187(w_in_5_187), .w_in_5_188(w_in_5_188), .w_in_5_189(w_in_5_189), .w_in_5_190(w_in_5_190), .w_in_5_191(w_in_5_191), .w_in_5_192(w_in_5_192), .w_in_5_193(w_in_5_193), .w_in_5_194(w_in_5_194), .w_in_5_195(w_in_5_195), .w_in_5_196(w_in_5_196), .w_in_5_197(w_in_5_197), .w_in_5_198(w_in_5_198), .w_in_5_199(w_in_5_199), .w_in_5_200(w_in_5_200), .w_in_5_201(w_in_5_201), .w_in_5_202(w_in_5_202), .w_in_5_203(w_in_5_203), .w_in_5_204(w_in_5_204), .w_in_5_205(w_in_5_205), .w_in_5_206(w_in_5_206), .w_in_5_207(w_in_5_207), .w_in_5_208(w_in_5_208), .w_in_5_209(w_in_5_209), .w_in_5_210(w_in_5_210), .w_in_5_211(w_in_5_211), .w_in_5_212(w_in_5_212), .w_in_5_213(w_in_5_213), .w_in_5_214(w_in_5_214), .w_in_5_215(w_in_5_215), .w_in_5_216(w_in_5_216), .w_in_5_217(w_in_5_217), .w_in_5_218(w_in_5_218), .w_in_5_219(w_in_5_219), .w_in_5_220(w_in_5_220), .w_in_5_221(w_in_5_221), .w_in_5_222(w_in_5_222), .w_in_5_223(w_in_5_223), .w_in_5_224(w_in_5_224), .w_in_5_225(w_in_5_225), .w_in_5_226(w_in_5_226), .w_in_5_227(w_in_5_227), .w_in_5_228(w_in_5_228), .w_in_5_229(w_in_5_229), .w_in_5_230(w_in_5_230), .w_in_5_231(w_in_5_231), .w_in_5_232(w_in_5_232), .w_in_5_233(w_in_5_233), .w_in_5_234(w_in_5_234), .w_in_5_235(w_in_5_235), .w_in_5_236(w_in_5_236), .w_in_5_237(w_in_5_237), .w_in_5_238(w_in_5_238), .w_in_5_239(w_in_5_239), .w_in_5_240(w_in_5_240), .w_in_5_241(w_in_5_241), .w_in_5_242(w_in_5_242), .w_in_5_243(w_in_5_243), .w_in_5_244(w_in_5_244), .w_in_5_245(w_in_5_245), .w_in_5_246(w_in_5_246), .w_in_5_247(w_in_5_247), .w_in_5_248(w_in_5_248), .w_in_5_249(w_in_5_249), .w_in_5_250(w_in_5_250), .w_in_5_251(w_in_5_251), .w_in_5_252(w_in_5_252), .w_in_5_253(w_in_5_253), .w_in_5_254(w_in_5_254), .w_in_5_255(w_in_5_255), .w_in_6_0(w_in_6_0), .w_in_6_1(w_in_6_1), .w_in_6_2(w_in_6_2), .w_in_6_3(w_in_6_3), .w_in_6_4(w_in_6_4), .w_in_6_5(w_in_6_5), .w_in_6_6(w_in_6_6), .w_in_6_7(w_in_6_7), .w_in_6_8(w_in_6_8), .w_in_6_9(w_in_6_9), .w_in_6_10(w_in_6_10), .w_in_6_11(w_in_6_11), .w_in_6_12(w_in_6_12), .w_in_6_13(w_in_6_13), .w_in_6_14(w_in_6_14), .w_in_6_15(w_in_6_15), .w_in_6_16(w_in_6_16), .w_in_6_17(w_in_6_17), .w_in_6_18(w_in_6_18), .w_in_6_19(w_in_6_19), .w_in_6_20(w_in_6_20), .w_in_6_21(w_in_6_21), .w_in_6_22(w_in_6_22), .w_in_6_23(w_in_6_23), .w_in_6_24(w_in_6_24), .w_in_6_25(w_in_6_25), .w_in_6_26(w_in_6_26), .w_in_6_27(w_in_6_27), .w_in_6_28(w_in_6_28), .w_in_6_29(w_in_6_29), .w_in_6_30(w_in_6_30), .w_in_6_31(w_in_6_31), .w_in_6_32(w_in_6_32), .w_in_6_33(w_in_6_33), .w_in_6_34(w_in_6_34), .w_in_6_35(w_in_6_35), .w_in_6_36(w_in_6_36), .w_in_6_37(w_in_6_37), .w_in_6_38(w_in_6_38), .w_in_6_39(w_in_6_39), .w_in_6_40(w_in_6_40), .w_in_6_41(w_in_6_41), .w_in_6_42(w_in_6_42), .w_in_6_43(w_in_6_43), .w_in_6_44(w_in_6_44), .w_in_6_45(w_in_6_45), .w_in_6_46(w_in_6_46), .w_in_6_47(w_in_6_47), .w_in_6_48(w_in_6_48), .w_in_6_49(w_in_6_49), .w_in_6_50(w_in_6_50), .w_in_6_51(w_in_6_51), .w_in_6_52(w_in_6_52), .w_in_6_53(w_in_6_53), .w_in_6_54(w_in_6_54), .w_in_6_55(w_in_6_55), .w_in_6_56(w_in_6_56), .w_in_6_57(w_in_6_57), .w_in_6_58(w_in_6_58), .w_in_6_59(w_in_6_59), .w_in_6_60(w_in_6_60), .w_in_6_61(w_in_6_61), .w_in_6_62(w_in_6_62), .w_in_6_63(w_in_6_63), .w_in_6_64(w_in_6_64), .w_in_6_65(w_in_6_65), .w_in_6_66(w_in_6_66), .w_in_6_67(w_in_6_67), .w_in_6_68(w_in_6_68), .w_in_6_69(w_in_6_69), .w_in_6_70(w_in_6_70), .w_in_6_71(w_in_6_71), .w_in_6_72(w_in_6_72), .w_in_6_73(w_in_6_73), .w_in_6_74(w_in_6_74), .w_in_6_75(w_in_6_75), .w_in_6_76(w_in_6_76), .w_in_6_77(w_in_6_77), .w_in_6_78(w_in_6_78), .w_in_6_79(w_in_6_79), .w_in_6_80(w_in_6_80), .w_in_6_81(w_in_6_81), .w_in_6_82(w_in_6_82), .w_in_6_83(w_in_6_83), .w_in_6_84(w_in_6_84), .w_in_6_85(w_in_6_85), .w_in_6_86(w_in_6_86), .w_in_6_87(w_in_6_87), .w_in_6_88(w_in_6_88), .w_in_6_89(w_in_6_89), .w_in_6_90(w_in_6_90), .w_in_6_91(w_in_6_91), .w_in_6_92(w_in_6_92), .w_in_6_93(w_in_6_93), .w_in_6_94(w_in_6_94), .w_in_6_95(w_in_6_95), .w_in_6_96(w_in_6_96), .w_in_6_97(w_in_6_97), .w_in_6_98(w_in_6_98), .w_in_6_99(w_in_6_99), .w_in_6_100(w_in_6_100), .w_in_6_101(w_in_6_101), .w_in_6_102(w_in_6_102), .w_in_6_103(w_in_6_103), .w_in_6_104(w_in_6_104), .w_in_6_105(w_in_6_105), .w_in_6_106(w_in_6_106), .w_in_6_107(w_in_6_107), .w_in_6_108(w_in_6_108), .w_in_6_109(w_in_6_109), .w_in_6_110(w_in_6_110), .w_in_6_111(w_in_6_111), .w_in_6_112(w_in_6_112), .w_in_6_113(w_in_6_113), .w_in_6_114(w_in_6_114), .w_in_6_115(w_in_6_115), .w_in_6_116(w_in_6_116), .w_in_6_117(w_in_6_117), .w_in_6_118(w_in_6_118), .w_in_6_119(w_in_6_119), .w_in_6_120(w_in_6_120), .w_in_6_121(w_in_6_121), .w_in_6_122(w_in_6_122), .w_in_6_123(w_in_6_123), .w_in_6_124(w_in_6_124), .w_in_6_125(w_in_6_125), .w_in_6_126(w_in_6_126), .w_in_6_127(w_in_6_127), .w_in_6_128(w_in_6_128), .w_in_6_129(w_in_6_129), .w_in_6_130(w_in_6_130), .w_in_6_131(w_in_6_131), .w_in_6_132(w_in_6_132), .w_in_6_133(w_in_6_133), .w_in_6_134(w_in_6_134), .w_in_6_135(w_in_6_135), .w_in_6_136(w_in_6_136), .w_in_6_137(w_in_6_137), .w_in_6_138(w_in_6_138), .w_in_6_139(w_in_6_139), .w_in_6_140(w_in_6_140), .w_in_6_141(w_in_6_141), .w_in_6_142(w_in_6_142), .w_in_6_143(w_in_6_143), .w_in_6_144(w_in_6_144), .w_in_6_145(w_in_6_145), .w_in_6_146(w_in_6_146), .w_in_6_147(w_in_6_147), .w_in_6_148(w_in_6_148), .w_in_6_149(w_in_6_149), .w_in_6_150(w_in_6_150), .w_in_6_151(w_in_6_151), .w_in_6_152(w_in_6_152), .w_in_6_153(w_in_6_153), .w_in_6_154(w_in_6_154), .w_in_6_155(w_in_6_155), .w_in_6_156(w_in_6_156), .w_in_6_157(w_in_6_157), .w_in_6_158(w_in_6_158), .w_in_6_159(w_in_6_159), .w_in_6_160(w_in_6_160), .w_in_6_161(w_in_6_161), .w_in_6_162(w_in_6_162), .w_in_6_163(w_in_6_163), .w_in_6_164(w_in_6_164), .w_in_6_165(w_in_6_165), .w_in_6_166(w_in_6_166), .w_in_6_167(w_in_6_167), .w_in_6_168(w_in_6_168), .w_in_6_169(w_in_6_169), .w_in_6_170(w_in_6_170), .w_in_6_171(w_in_6_171), .w_in_6_172(w_in_6_172), .w_in_6_173(w_in_6_173), .w_in_6_174(w_in_6_174), .w_in_6_175(w_in_6_175), .w_in_6_176(w_in_6_176), .w_in_6_177(w_in_6_177), .w_in_6_178(w_in_6_178), .w_in_6_179(w_in_6_179), .w_in_6_180(w_in_6_180), .w_in_6_181(w_in_6_181), .w_in_6_182(w_in_6_182), .w_in_6_183(w_in_6_183), .w_in_6_184(w_in_6_184), .w_in_6_185(w_in_6_185), .w_in_6_186(w_in_6_186), .w_in_6_187(w_in_6_187), .w_in_6_188(w_in_6_188), .w_in_6_189(w_in_6_189), .w_in_6_190(w_in_6_190), .w_in_6_191(w_in_6_191), .w_in_6_192(w_in_6_192), .w_in_6_193(w_in_6_193), .w_in_6_194(w_in_6_194), .w_in_6_195(w_in_6_195), .w_in_6_196(w_in_6_196), .w_in_6_197(w_in_6_197), .w_in_6_198(w_in_6_198), .w_in_6_199(w_in_6_199), .w_in_6_200(w_in_6_200), .w_in_6_201(w_in_6_201), .w_in_6_202(w_in_6_202), .w_in_6_203(w_in_6_203), .w_in_6_204(w_in_6_204), .w_in_6_205(w_in_6_205), .w_in_6_206(w_in_6_206), .w_in_6_207(w_in_6_207), .w_in_6_208(w_in_6_208), .w_in_6_209(w_in_6_209), .w_in_6_210(w_in_6_210), .w_in_6_211(w_in_6_211), .w_in_6_212(w_in_6_212), .w_in_6_213(w_in_6_213), .w_in_6_214(w_in_6_214), .w_in_6_215(w_in_6_215), .w_in_6_216(w_in_6_216), .w_in_6_217(w_in_6_217), .w_in_6_218(w_in_6_218), .w_in_6_219(w_in_6_219), .w_in_6_220(w_in_6_220), .w_in_6_221(w_in_6_221), .w_in_6_222(w_in_6_222), .w_in_6_223(w_in_6_223), .w_in_6_224(w_in_6_224), .w_in_6_225(w_in_6_225), .w_in_6_226(w_in_6_226), .w_in_6_227(w_in_6_227), .w_in_6_228(w_in_6_228), .w_in_6_229(w_in_6_229), .w_in_6_230(w_in_6_230), .w_in_6_231(w_in_6_231), .w_in_6_232(w_in_6_232), .w_in_6_233(w_in_6_233), .w_in_6_234(w_in_6_234), .w_in_6_235(w_in_6_235), .w_in_6_236(w_in_6_236), .w_in_6_237(w_in_6_237), .w_in_6_238(w_in_6_238), .w_in_6_239(w_in_6_239), .w_in_6_240(w_in_6_240), .w_in_6_241(w_in_6_241), .w_in_6_242(w_in_6_242), .w_in_6_243(w_in_6_243), .w_in_6_244(w_in_6_244), .w_in_6_245(w_in_6_245), .w_in_6_246(w_in_6_246), .w_in_6_247(w_in_6_247), .w_in_6_248(w_in_6_248), .w_in_6_249(w_in_6_249), .w_in_6_250(w_in_6_250), .w_in_6_251(w_in_6_251), .w_in_6_252(w_in_6_252), .w_in_6_253(w_in_6_253), .w_in_6_254(w_in_6_254), .w_in_6_255(w_in_6_255), .w_in_7_0(w_in_7_0), .w_in_7_1(w_in_7_1), .w_in_7_2(w_in_7_2), .w_in_7_3(w_in_7_3), .w_in_7_4(w_in_7_4), .w_in_7_5(w_in_7_5), .w_in_7_6(w_in_7_6), .w_in_7_7(w_in_7_7), .w_in_7_8(w_in_7_8), .w_in_7_9(w_in_7_9), .w_in_7_10(w_in_7_10), .w_in_7_11(w_in_7_11), .w_in_7_12(w_in_7_12), .w_in_7_13(w_in_7_13), .w_in_7_14(w_in_7_14), .w_in_7_15(w_in_7_15), .w_in_7_16(w_in_7_16), .w_in_7_17(w_in_7_17), .w_in_7_18(w_in_7_18), .w_in_7_19(w_in_7_19), .w_in_7_20(w_in_7_20), .w_in_7_21(w_in_7_21), .w_in_7_22(w_in_7_22), .w_in_7_23(w_in_7_23), .w_in_7_24(w_in_7_24), .w_in_7_25(w_in_7_25), .w_in_7_26(w_in_7_26), .w_in_7_27(w_in_7_27), .w_in_7_28(w_in_7_28), .w_in_7_29(w_in_7_29), .w_in_7_30(w_in_7_30), .w_in_7_31(w_in_7_31), .w_in_7_32(w_in_7_32), .w_in_7_33(w_in_7_33), .w_in_7_34(w_in_7_34), .w_in_7_35(w_in_7_35), .w_in_7_36(w_in_7_36), .w_in_7_37(w_in_7_37), .w_in_7_38(w_in_7_38), .w_in_7_39(w_in_7_39), .w_in_7_40(w_in_7_40), .w_in_7_41(w_in_7_41), .w_in_7_42(w_in_7_42), .w_in_7_43(w_in_7_43), .w_in_7_44(w_in_7_44), .w_in_7_45(w_in_7_45), .w_in_7_46(w_in_7_46), .w_in_7_47(w_in_7_47), .w_in_7_48(w_in_7_48), .w_in_7_49(w_in_7_49), .w_in_7_50(w_in_7_50), .w_in_7_51(w_in_7_51), .w_in_7_52(w_in_7_52), .w_in_7_53(w_in_7_53), .w_in_7_54(w_in_7_54), .w_in_7_55(w_in_7_55), .w_in_7_56(w_in_7_56), .w_in_7_57(w_in_7_57), .w_in_7_58(w_in_7_58), .w_in_7_59(w_in_7_59), .w_in_7_60(w_in_7_60), .w_in_7_61(w_in_7_61), .w_in_7_62(w_in_7_62), .w_in_7_63(w_in_7_63), .w_in_7_64(w_in_7_64), .w_in_7_65(w_in_7_65), .w_in_7_66(w_in_7_66), .w_in_7_67(w_in_7_67), .w_in_7_68(w_in_7_68), .w_in_7_69(w_in_7_69), .w_in_7_70(w_in_7_70), .w_in_7_71(w_in_7_71), .w_in_7_72(w_in_7_72), .w_in_7_73(w_in_7_73), .w_in_7_74(w_in_7_74), .w_in_7_75(w_in_7_75), .w_in_7_76(w_in_7_76), .w_in_7_77(w_in_7_77), .w_in_7_78(w_in_7_78), .w_in_7_79(w_in_7_79), .w_in_7_80(w_in_7_80), .w_in_7_81(w_in_7_81), .w_in_7_82(w_in_7_82), .w_in_7_83(w_in_7_83), .w_in_7_84(w_in_7_84), .w_in_7_85(w_in_7_85), .w_in_7_86(w_in_7_86), .w_in_7_87(w_in_7_87), .w_in_7_88(w_in_7_88), .w_in_7_89(w_in_7_89), .w_in_7_90(w_in_7_90), .w_in_7_91(w_in_7_91), .w_in_7_92(w_in_7_92), .w_in_7_93(w_in_7_93), .w_in_7_94(w_in_7_94), .w_in_7_95(w_in_7_95), .w_in_7_96(w_in_7_96), .w_in_7_97(w_in_7_97), .w_in_7_98(w_in_7_98), .w_in_7_99(w_in_7_99), .w_in_7_100(w_in_7_100), .w_in_7_101(w_in_7_101), .w_in_7_102(w_in_7_102), .w_in_7_103(w_in_7_103), .w_in_7_104(w_in_7_104), .w_in_7_105(w_in_7_105), .w_in_7_106(w_in_7_106), .w_in_7_107(w_in_7_107), .w_in_7_108(w_in_7_108), .w_in_7_109(w_in_7_109), .w_in_7_110(w_in_7_110), .w_in_7_111(w_in_7_111), .w_in_7_112(w_in_7_112), .w_in_7_113(w_in_7_113), .w_in_7_114(w_in_7_114), .w_in_7_115(w_in_7_115), .w_in_7_116(w_in_7_116), .w_in_7_117(w_in_7_117), .w_in_7_118(w_in_7_118), .w_in_7_119(w_in_7_119), .w_in_7_120(w_in_7_120), .w_in_7_121(w_in_7_121), .w_in_7_122(w_in_7_122), .w_in_7_123(w_in_7_123), .w_in_7_124(w_in_7_124), .w_in_7_125(w_in_7_125), .w_in_7_126(w_in_7_126), .w_in_7_127(w_in_7_127), .w_in_7_128(w_in_7_128), .w_in_7_129(w_in_7_129), .w_in_7_130(w_in_7_130), .w_in_7_131(w_in_7_131), .w_in_7_132(w_in_7_132), .w_in_7_133(w_in_7_133), .w_in_7_134(w_in_7_134), .w_in_7_135(w_in_7_135), .w_in_7_136(w_in_7_136), .w_in_7_137(w_in_7_137), .w_in_7_138(w_in_7_138), .w_in_7_139(w_in_7_139), .w_in_7_140(w_in_7_140), .w_in_7_141(w_in_7_141), .w_in_7_142(w_in_7_142), .w_in_7_143(w_in_7_143), .w_in_7_144(w_in_7_144), .w_in_7_145(w_in_7_145), .w_in_7_146(w_in_7_146), .w_in_7_147(w_in_7_147), .w_in_7_148(w_in_7_148), .w_in_7_149(w_in_7_149), .w_in_7_150(w_in_7_150), .w_in_7_151(w_in_7_151), .w_in_7_152(w_in_7_152), .w_in_7_153(w_in_7_153), .w_in_7_154(w_in_7_154), .w_in_7_155(w_in_7_155), .w_in_7_156(w_in_7_156), .w_in_7_157(w_in_7_157), .w_in_7_158(w_in_7_158), .w_in_7_159(w_in_7_159), .w_in_7_160(w_in_7_160), .w_in_7_161(w_in_7_161), .w_in_7_162(w_in_7_162), .w_in_7_163(w_in_7_163), .w_in_7_164(w_in_7_164), .w_in_7_165(w_in_7_165), .w_in_7_166(w_in_7_166), .w_in_7_167(w_in_7_167), .w_in_7_168(w_in_7_168), .w_in_7_169(w_in_7_169), .w_in_7_170(w_in_7_170), .w_in_7_171(w_in_7_171), .w_in_7_172(w_in_7_172), .w_in_7_173(w_in_7_173), .w_in_7_174(w_in_7_174), .w_in_7_175(w_in_7_175), .w_in_7_176(w_in_7_176), .w_in_7_177(w_in_7_177), .w_in_7_178(w_in_7_178), .w_in_7_179(w_in_7_179), .w_in_7_180(w_in_7_180), .w_in_7_181(w_in_7_181), .w_in_7_182(w_in_7_182), .w_in_7_183(w_in_7_183), .w_in_7_184(w_in_7_184), .w_in_7_185(w_in_7_185), .w_in_7_186(w_in_7_186), .w_in_7_187(w_in_7_187), .w_in_7_188(w_in_7_188), .w_in_7_189(w_in_7_189), .w_in_7_190(w_in_7_190), .w_in_7_191(w_in_7_191), .w_in_7_192(w_in_7_192), .w_in_7_193(w_in_7_193), .w_in_7_194(w_in_7_194), .w_in_7_195(w_in_7_195), .w_in_7_196(w_in_7_196), .w_in_7_197(w_in_7_197), .w_in_7_198(w_in_7_198), .w_in_7_199(w_in_7_199), .w_in_7_200(w_in_7_200), .w_in_7_201(w_in_7_201), .w_in_7_202(w_in_7_202), .w_in_7_203(w_in_7_203), .w_in_7_204(w_in_7_204), .w_in_7_205(w_in_7_205), .w_in_7_206(w_in_7_206), .w_in_7_207(w_in_7_207), .w_in_7_208(w_in_7_208), .w_in_7_209(w_in_7_209), .w_in_7_210(w_in_7_210), .w_in_7_211(w_in_7_211), .w_in_7_212(w_in_7_212), .w_in_7_213(w_in_7_213), .w_in_7_214(w_in_7_214), .w_in_7_215(w_in_7_215), .w_in_7_216(w_in_7_216), .w_in_7_217(w_in_7_217), .w_in_7_218(w_in_7_218), .w_in_7_219(w_in_7_219), .w_in_7_220(w_in_7_220), .w_in_7_221(w_in_7_221), .w_in_7_222(w_in_7_222), .w_in_7_223(w_in_7_223), .w_in_7_224(w_in_7_224), .w_in_7_225(w_in_7_225), .w_in_7_226(w_in_7_226), .w_in_7_227(w_in_7_227), .w_in_7_228(w_in_7_228), .w_in_7_229(w_in_7_229), .w_in_7_230(w_in_7_230), .w_in_7_231(w_in_7_231), .w_in_7_232(w_in_7_232), .w_in_7_233(w_in_7_233), .w_in_7_234(w_in_7_234), .w_in_7_235(w_in_7_235), .w_in_7_236(w_in_7_236), .w_in_7_237(w_in_7_237), .w_in_7_238(w_in_7_238), .w_in_7_239(w_in_7_239), .w_in_7_240(w_in_7_240), .w_in_7_241(w_in_7_241), .w_in_7_242(w_in_7_242), .w_in_7_243(w_in_7_243), .w_in_7_244(w_in_7_244), .w_in_7_245(w_in_7_245), .w_in_7_246(w_in_7_246), .w_in_7_247(w_in_7_247), .w_in_7_248(w_in_7_248), .w_in_7_249(w_in_7_249), .w_in_7_250(w_in_7_250), .w_in_7_251(w_in_7_251), .w_in_7_252(w_in_7_252), .w_in_7_253(w_in_7_253), .w_in_7_254(w_in_7_254), .w_in_7_255(w_in_7_255), 
.w_hr_0_0(w_hr_0_0), .w_hr_0_1(w_hr_0_1), .w_hr_0_2(w_hr_0_2), .w_hr_0_3(w_hr_0_3), .w_hr_0_4(w_hr_0_4), .w_hr_0_5(w_hr_0_5), .w_hr_0_6(w_hr_0_6), .w_hr_0_7(w_hr_0_7), .w_hr_1_0(w_hr_1_0), .w_hr_1_1(w_hr_1_1), .w_hr_1_2(w_hr_1_2), .w_hr_1_3(w_hr_1_3), .w_hr_1_4(w_hr_1_4), .w_hr_1_5(w_hr_1_5), .w_hr_1_6(w_hr_1_6), .w_hr_1_7(w_hr_1_7), .w_hr_2_0(w_hr_2_0), .w_hr_2_1(w_hr_2_1), .w_hr_2_2(w_hr_2_2), .w_hr_2_3(w_hr_2_3), .w_hr_2_4(w_hr_2_4), .w_hr_2_5(w_hr_2_5), .w_hr_2_6(w_hr_2_6), .w_hr_2_7(w_hr_2_7), .w_hr_3_0(w_hr_3_0), .w_hr_3_1(w_hr_3_1), .w_hr_3_2(w_hr_3_2), .w_hr_3_3(w_hr_3_3), .w_hr_3_4(w_hr_3_4), .w_hr_3_5(w_hr_3_5), .w_hr_3_6(w_hr_3_6), .w_hr_3_7(w_hr_3_7), .w_hr_4_0(w_hr_4_0), .w_hr_4_1(w_hr_4_1), .w_hr_4_2(w_hr_4_2), .w_hr_4_3(w_hr_4_3), .w_hr_4_4(w_hr_4_4), .w_hr_4_5(w_hr_4_5), .w_hr_4_6(w_hr_4_6), .w_hr_4_7(w_hr_4_7), .w_hr_5_0(w_hr_5_0), .w_hr_5_1(w_hr_5_1), .w_hr_5_2(w_hr_5_2), .w_hr_5_3(w_hr_5_3), .w_hr_5_4(w_hr_5_4), .w_hr_5_5(w_hr_5_5), .w_hr_5_6(w_hr_5_6), .w_hr_5_7(w_hr_5_7), .w_hr_6_0(w_hr_6_0), .w_hr_6_1(w_hr_6_1), .w_hr_6_2(w_hr_6_2), .w_hr_6_3(w_hr_6_3), .w_hr_6_4(w_hr_6_4), .w_hr_6_5(w_hr_6_5), .w_hr_6_6(w_hr_6_6), .w_hr_6_7(w_hr_6_7), .w_hr_7_0(w_hr_7_0), .w_hr_7_1(w_hr_7_1), .w_hr_7_2(w_hr_7_2), .w_hr_7_3(w_hr_7_3), .w_hr_7_4(w_hr_7_4), .w_hr_7_5(w_hr_7_5), .w_hr_7_6(w_hr_7_6), .w_hr_7_7(w_hr_7_7), 
.w_hz_0_0(w_hz_0_0), .w_hz_0_1(w_hz_0_1), .w_hz_0_2(w_hz_0_2), .w_hz_0_3(w_hz_0_3), .w_hz_0_4(w_hz_0_4), .w_hz_0_5(w_hz_0_5), .w_hz_0_6(w_hz_0_6), .w_hz_0_7(w_hz_0_7), .w_hz_1_0(w_hz_1_0), .w_hz_1_1(w_hz_1_1), .w_hz_1_2(w_hz_1_2), .w_hz_1_3(w_hz_1_3), .w_hz_1_4(w_hz_1_4), .w_hz_1_5(w_hz_1_5), .w_hz_1_6(w_hz_1_6), .w_hz_1_7(w_hz_1_7), .w_hz_2_0(w_hz_2_0), .w_hz_2_1(w_hz_2_1), .w_hz_2_2(w_hz_2_2), .w_hz_2_3(w_hz_2_3), .w_hz_2_4(w_hz_2_4), .w_hz_2_5(w_hz_2_5), .w_hz_2_6(w_hz_2_6), .w_hz_2_7(w_hz_2_7), .w_hz_3_0(w_hz_3_0), .w_hz_3_1(w_hz_3_1), .w_hz_3_2(w_hz_3_2), .w_hz_3_3(w_hz_3_3), .w_hz_3_4(w_hz_3_4), .w_hz_3_5(w_hz_3_5), .w_hz_3_6(w_hz_3_6), .w_hz_3_7(w_hz_3_7), .w_hz_4_0(w_hz_4_0), .w_hz_4_1(w_hz_4_1), .w_hz_4_2(w_hz_4_2), .w_hz_4_3(w_hz_4_3), .w_hz_4_4(w_hz_4_4), .w_hz_4_5(w_hz_4_5), .w_hz_4_6(w_hz_4_6), .w_hz_4_7(w_hz_4_7), .w_hz_5_0(w_hz_5_0), .w_hz_5_1(w_hz_5_1), .w_hz_5_2(w_hz_5_2), .w_hz_5_3(w_hz_5_3), .w_hz_5_4(w_hz_5_4), .w_hz_5_5(w_hz_5_5), .w_hz_5_6(w_hz_5_6), .w_hz_5_7(w_hz_5_7), .w_hz_6_0(w_hz_6_0), .w_hz_6_1(w_hz_6_1), .w_hz_6_2(w_hz_6_2), .w_hz_6_3(w_hz_6_3), .w_hz_6_4(w_hz_6_4), .w_hz_6_5(w_hz_6_5), .w_hz_6_6(w_hz_6_6), .w_hz_6_7(w_hz_6_7), .w_hz_7_0(w_hz_7_0), .w_hz_7_1(w_hz_7_1), .w_hz_7_2(w_hz_7_2), .w_hz_7_3(w_hz_7_3), .w_hz_7_4(w_hz_7_4), .w_hz_7_5(w_hz_7_5), .w_hz_7_6(w_hz_7_6), .w_hz_7_7(w_hz_7_7), 
.w_hn_0_0(w_hn_0_0), .w_hn_0_1(w_hn_0_1), .w_hn_0_2(w_hn_0_2), .w_hn_0_3(w_hn_0_3), .w_hn_0_4(w_hn_0_4), .w_hn_0_5(w_hn_0_5), .w_hn_0_6(w_hn_0_6), .w_hn_0_7(w_hn_0_7), .w_hn_1_0(w_hn_1_0), .w_hn_1_1(w_hn_1_1), .w_hn_1_2(w_hn_1_2), .w_hn_1_3(w_hn_1_3), .w_hn_1_4(w_hn_1_4), .w_hn_1_5(w_hn_1_5), .w_hn_1_6(w_hn_1_6), .w_hn_1_7(w_hn_1_7), .w_hn_2_0(w_hn_2_0), .w_hn_2_1(w_hn_2_1), .w_hn_2_2(w_hn_2_2), .w_hn_2_3(w_hn_2_3), .w_hn_2_4(w_hn_2_4), .w_hn_2_5(w_hn_2_5), .w_hn_2_6(w_hn_2_6), .w_hn_2_7(w_hn_2_7), .w_hn_3_0(w_hn_3_0), .w_hn_3_1(w_hn_3_1), .w_hn_3_2(w_hn_3_2), .w_hn_3_3(w_hn_3_3), .w_hn_3_4(w_hn_3_4), .w_hn_3_5(w_hn_3_5), .w_hn_3_6(w_hn_3_6), .w_hn_3_7(w_hn_3_7), .w_hn_4_0(w_hn_4_0), .w_hn_4_1(w_hn_4_1), .w_hn_4_2(w_hn_4_2), .w_hn_4_3(w_hn_4_3), .w_hn_4_4(w_hn_4_4), .w_hn_4_5(w_hn_4_5), .w_hn_4_6(w_hn_4_6), .w_hn_4_7(w_hn_4_7), .w_hn_5_0(w_hn_5_0), .w_hn_5_1(w_hn_5_1), .w_hn_5_2(w_hn_5_2), .w_hn_5_3(w_hn_5_3), .w_hn_5_4(w_hn_5_4), .w_hn_5_5(w_hn_5_5), .w_hn_5_6(w_hn_5_6), .w_hn_5_7(w_hn_5_7), .w_hn_6_0(w_hn_6_0), .w_hn_6_1(w_hn_6_1), .w_hn_6_2(w_hn_6_2), .w_hn_6_3(w_hn_6_3), .w_hn_6_4(w_hn_6_4), .w_hn_6_5(w_hn_6_5), .w_hn_6_6(w_hn_6_6), .w_hn_6_7(w_hn_6_7), .w_hn_7_0(w_hn_7_0), .w_hn_7_1(w_hn_7_1), .w_hn_7_2(w_hn_7_2), .w_hn_7_3(w_hn_7_3), .w_hn_7_4(w_hn_7_4), .w_hn_7_5(w_hn_7_5), .w_hn_7_6(w_hn_7_6), .w_hn_7_7(w_hn_7_7), 
.b_ir_0(b_ir_0), .b_ir_1(b_ir_1), .b_ir_2(b_ir_2), .b_ir_3(b_ir_3), .b_ir_4(b_ir_4), .b_ir_5(b_ir_5), .b_ir_6(b_ir_6), .b_ir_7(b_ir_7), 
.b_iz_0(b_iz_0), .b_iz_1(b_iz_1), .b_iz_2(b_iz_2), .b_iz_3(b_iz_3), .b_iz_4(b_iz_4), .b_iz_5(b_iz_5), .b_iz_6(b_iz_6), .b_iz_7(b_iz_7), 
.b_in_0(b_in_0), .b_in_1(b_in_1), .b_in_2(b_in_2), .b_in_3(b_in_3), .b_in_4(b_in_4), .b_in_5(b_in_5), .b_in_6(b_in_6), .b_in_7(b_in_7), 
.b_hr_0(b_hr_0), .b_hr_1(b_hr_1), .b_hr_2(b_hr_2), .b_hr_3(b_hr_3), .b_hr_4(b_hr_4), .b_hr_5(b_hr_5), .b_hr_6(b_hr_6), .b_hr_7(b_hr_7), 
.b_hz_0(b_hz_0), .b_hz_1(b_hz_1), .b_hz_2(b_hz_2), .b_hz_3(b_hz_3), .b_hz_4(b_hz_4), .b_hz_5(b_hz_5), .b_hz_6(b_hz_6), .b_hz_7(b_hz_7), 
.b_hn_0(b_hn_0), .b_hn_1(b_hn_1), .b_hn_2(b_hn_2), .b_hn_3(b_hn_3), .b_hn_4(b_hn_4), .b_hn_5(b_hn_5), .b_hn_6(b_hn_6), .b_hn_7(b_hn_7), 
.y_0(y_0), .y_1(y_1), .y_2(y_2), .y_3(y_3), .y_4(y_4), .y_5(y_5), .y_6(y_6), .y_7(y_7)
);

    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end
    
    initial begin
        // Open file for writing (overwrite existing)
        integer fd;
        fd = $fopen("../../../../../output_d256_h8_int4_frac5.txt", "w+");
        if (fd == 0) begin
            $display("ERROR: Failed to open file!");
            $finish;
        end
        x_0 = 'b000100100;
    x_1 = 'b000110111;
    x_2 = 'b001000001;
    x_3 = 'b001001001;
    x_4 = 'b000111011;
    x_5 = 'b000110110;
    x_6 = 'b000100111;
    x_7 = 'b000100101;
    x_8 = 'b000111100;
    x_9 = 'b001001000;
    x_10 = 'b001001011;
    x_11 = 'b001001001;
    x_12 = 'b001000111;
    x_13 = 'b000101101;
    x_14 = 'b000111011;
    x_15 = 'b001000110;
    x_16 = 'b001001010;
    x_17 = 'b001001101;
    x_18 = 'b001001111;
    x_19 = 'b001001110;
    x_20 = 'b000110111;
    x_21 = 'b000010001;
    x_22 = 'b000010100;
    x_23 = 'b000010111;
    x_24 = 'b000001100;
    x_25 = 'b000001110;
    x_26 = 'b000101001;
    x_27 = 'b000011100;
    x_28 = 'b000011110;
    x_29 = 'b000001100;
    x_30 = 'b000011000;
    x_31 = 'b000110010;
    x_32 = 'b000111110;
    x_33 = 'b000111110;
    x_34 = 'b000111000;
    x_35 = 'b000101111;
    x_36 = 'b000101000;
    x_37 = 'b000010100;
    x_38 = 'b000010111;
    x_39 = 'b000100100;
    x_40 = 'b000101010;
    x_41 = 'b000110100;
    x_42 = 'b000100000;
    x_43 = 'b000011011;
    x_44 = 'b000110001;
    x_45 = 'b000010111;
    x_46 = 'b000111011;
    x_47 = 'b001000011;
    x_48 = 'b000111111;
    x_49 = 'b001000110;
    x_50 = 'b001010001;
    x_51 = 'b001010101;
    x_52 = 'b001010001;
    x_53 = 'b001000110;
    x_54 = 'b000110111;
    x_55 = 'b000110111;
    x_56 = 'b001000011;
    x_57 = 'b001000110;
    x_58 = 'b001001001;
    x_59 = 'b000101111;
    x_60 = 'b000110000;
    x_61 = 'b000110011;
    x_62 = 'b000100101;
    x_63 = 'b000110000;
    x_64 = 'b000100100;
    x_65 = 'b000110111;
    x_66 = 'b001000001;
    x_67 = 'b001001001;
    x_68 = 'b000111011;
    x_69 = 'b000110110;
    x_70 = 'b000100111;
    x_71 = 'b000100101;
    x_72 = 'b000111100;
    x_73 = 'b001001000;
    x_74 = 'b001001011;
    x_75 = 'b001001001;
    x_76 = 'b001000111;
    x_77 = 'b000101101;
    x_78 = 'b000111011;
    x_79 = 'b001000110;
    x_80 = 'b001001010;
    x_81 = 'b001001101;
    x_82 = 'b001001111;
    x_83 = 'b001001110;
    x_84 = 'b000110111;
    x_85 = 'b000010001;
    x_86 = 'b000010100;
    x_87 = 'b000010111;
    x_88 = 'b000001100;
    x_89 = 'b000001110;
    x_90 = 'b000101001;
    x_91 = 'b000011100;
    x_92 = 'b000011110;
    x_93 = 'b000001100;
    x_94 = 'b000011000;
    x_95 = 'b000110010;
    x_96 = 'b000111110;
    x_97 = 'b000111110;
    x_98 = 'b000111000;
    x_99 = 'b000101111;
    x_100 = 'b000101000;
    x_101 = 'b000010100;
    x_102 = 'b000010111;
    x_103 = 'b000100100;
    x_104 = 'b000101010;
    x_105 = 'b000110100;
    x_106 = 'b000100000;
    x_107 = 'b000011011;
    x_108 = 'b000110001;
    x_109 = 'b000010111;
    x_110 = 'b000111011;
    x_111 = 'b001000011;
    x_112 = 'b000111111;
    x_113 = 'b001000110;
    x_114 = 'b001010001;
    x_115 = 'b001010101;
    x_116 = 'b001010001;
    x_117 = 'b001000110;
    x_118 = 'b000110111;
    x_119 = 'b000110111;
    x_120 = 'b001000011;
    x_121 = 'b001000110;
    x_122 = 'b001001001;
    x_123 = 'b000101111;
    x_124 = 'b000110000;
    x_125 = 'b000110011;
    x_126 = 'b000100101;
    x_127 = 'b000110000;
    x_128 = 'b000100100;
    x_129 = 'b000110111;
    x_130 = 'b001000001;
    x_131 = 'b001001001;
    x_132 = 'b000111011;
    x_133 = 'b000110110;
    x_134 = 'b000100111;
    x_135 = 'b000100101;
    x_136 = 'b000111100;
    x_137 = 'b001001000;
    x_138 = 'b001001011;
    x_139 = 'b001001001;
    x_140 = 'b001000111;
    x_141 = 'b000101101;
    x_142 = 'b000111011;
    x_143 = 'b001000110;
    x_144 = 'b001001010;
    x_145 = 'b001001101;
    x_146 = 'b001001111;
    x_147 = 'b001001110;
    x_148 = 'b000110111;
    x_149 = 'b000010001;
    x_150 = 'b000010100;
    x_151 = 'b000010111;
    x_152 = 'b000001100;
    x_153 = 'b000001110;
    x_154 = 'b000101001;
    x_155 = 'b000011100;
    x_156 = 'b000011110;
    x_157 = 'b000001100;
    x_158 = 'b000011000;
    x_159 = 'b000110010;
    x_160 = 'b000111110;
    x_161 = 'b000111110;
    x_162 = 'b000111000;
    x_163 = 'b000101111;
    x_164 = 'b000101000;
    x_165 = 'b000010100;
    x_166 = 'b000010111;
    x_167 = 'b000100100;
    x_168 = 'b000101010;
    x_169 = 'b000110100;
    x_170 = 'b000100000;
    x_171 = 'b000011011;
    x_172 = 'b000110001;
    x_173 = 'b000010111;
    x_174 = 'b000111011;
    x_175 = 'b001000011;
    x_176 = 'b000111111;
    x_177 = 'b001000110;
    x_178 = 'b001010001;
    x_179 = 'b001010101;
    x_180 = 'b001010001;
    x_181 = 'b001000110;
    x_182 = 'b000110111;
    x_183 = 'b000110111;
    x_184 = 'b001000011;
    x_185 = 'b001000110;
    x_186 = 'b001001001;
    x_187 = 'b000101111;
    x_188 = 'b000110000;
    x_189 = 'b000110011;
    x_190 = 'b000100101;
    x_191 = 'b000110000;
    x_192 = 'b000100100;
    x_193 = 'b000110111;
    x_194 = 'b001000001;
    x_195 = 'b001001001;
    x_196 = 'b000111011;
    x_197 = 'b000110110;
    x_198 = 'b000100111;
    x_199 = 'b000100101;
    x_200 = 'b000111100;
    x_201 = 'b001001000;
    x_202 = 'b001001011;
    x_203 = 'b001001001;
    x_204 = 'b001000111;
    x_205 = 'b000101101;
    x_206 = 'b000111011;
    x_207 = 'b001000110;
    x_208 = 'b001001010;
    x_209 = 'b001001101;
    x_210 = 'b001001111;
    x_211 = 'b001001110;
    x_212 = 'b000110111;
    x_213 = 'b000010001;
    x_214 = 'b000010100;
    x_215 = 'b000010111;
    x_216 = 'b000001100;
    x_217 = 'b000001110;
    x_218 = 'b000101001;
    x_219 = 'b000011100;
    x_220 = 'b000011110;
    x_221 = 'b000001100;
    x_222 = 'b000011000;
    x_223 = 'b000110010;
    x_224 = 'b000111110;
    x_225 = 'b000111110;
    x_226 = 'b000111000;
    x_227 = 'b000101111;
    x_228 = 'b000101000;
    x_229 = 'b000010100;
    x_230 = 'b000010111;
    x_231 = 'b000100100;
    x_232 = 'b000101010;
    x_233 = 'b000110100;
    x_234 = 'b000100000;
    x_235 = 'b000011011;
    x_236 = 'b000110001;
    x_237 = 'b000010111;
    x_238 = 'b000111011;
    x_239 = 'b001000011;
    x_240 = 'b000111111;
    x_241 = 'b001000110;
    x_242 = 'b001010001;
    x_243 = 'b001010101;
    x_244 = 'b001010001;
    x_245 = 'b001000110;
    x_246 = 'b000110111;
    x_247 = 'b000110111;
    x_248 = 'b001000011;
    x_249 = 'b001000110;
    x_250 = 'b001001001;
    x_251 = 'b000101111;
    x_252 = 'b000110000;
    x_253 = 'b000110011;
    x_254 = 'b000100101;
    x_255 = 'b000110000;

    h_0 = 'b000100100;
    h_1 = 'b000110111;
    h_2 = 'b001000001;
    h_3 = 'b001001001;
    h_4 = 'b000111011;
    h_5 = 'b000110110;
    h_6 = 'b000100111;
    h_7 = 'b000100101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000101110;
    x_1 = 'b001001001;
    x_2 = 'b001010010;
    x_3 = 'b001010101;
    x_4 = 'b001001111;
    x_5 = 'b001001100;
    x_6 = 'b000111111;
    x_7 = 'b000110111;
    x_8 = 'b001010001;
    x_9 = 'b001011010;
    x_10 = 'b001011011;
    x_11 = 'b001011111;
    x_12 = 'b001011010;
    x_13 = 'b001000000;
    x_14 = 'b001001101;
    x_15 = 'b001010111;
    x_16 = 'b001011000;
    x_17 = 'b001011101;
    x_18 = 'b001011110;
    x_19 = 'b001011101;
    x_20 = 'b001000011;
    x_21 = 'b000010011;
    x_22 = 'b000010100;
    x_23 = 'b000010110;
    x_24 = 'b000011000;
    x_25 = 'b000011010;
    x_26 = 'b000101101;
    x_27 = 'b000100001;
    x_28 = 'b000011010;
    x_29 = 'b000100011;
    x_30 = 'b000101010;
    x_31 = 'b000111000;
    x_32 = 'b001000010;
    x_33 = 'b001000000;
    x_34 = 'b000111010;
    x_35 = 'b000110101;
    x_36 = 'b000101001;
    x_37 = 'b000011001;
    x_38 = 'b000110101;
    x_39 = 'b000010110;
    x_40 = 'b001000010;
    x_41 = 'b111111101;
    x_42 = 'b000111010;
    x_43 = 'b000100101;
    x_44 = 'b001001000;
    x_45 = 'b000000101;
    x_46 = 'b001001001;
    x_47 = 'b001001001;
    x_48 = 'b001000000;
    x_49 = 'b001000001;
    x_50 = 'b001001110;
    x_51 = 'b001010010;
    x_52 = 'b001001001;
    x_53 = 'b000111100;
    x_54 = 'b000101010;
    x_55 = 'b000110101;
    x_56 = 'b000111110;
    x_57 = 'b000111110;
    x_58 = 'b001000010;
    x_59 = 'b000101001;
    x_60 = 'b000101110;
    x_61 = 'b000110100;
    x_62 = 'b000100110;
    x_63 = 'b000101101;
    x_64 = 'b000101110;
    x_65 = 'b001001001;
    x_66 = 'b001010010;
    x_67 = 'b001010101;
    x_68 = 'b001001111;
    x_69 = 'b001001100;
    x_70 = 'b000111111;
    x_71 = 'b000110111;
    x_72 = 'b001010001;
    x_73 = 'b001011010;
    x_74 = 'b001011011;
    x_75 = 'b001011111;
    x_76 = 'b001011010;
    x_77 = 'b001000000;
    x_78 = 'b001001101;
    x_79 = 'b001010111;
    x_80 = 'b001011000;
    x_81 = 'b001011101;
    x_82 = 'b001011110;
    x_83 = 'b001011101;
    x_84 = 'b001000011;
    x_85 = 'b000010011;
    x_86 = 'b000010100;
    x_87 = 'b000010110;
    x_88 = 'b000011000;
    x_89 = 'b000011010;
    x_90 = 'b000101101;
    x_91 = 'b000100001;
    x_92 = 'b000011010;
    x_93 = 'b000100011;
    x_94 = 'b000101010;
    x_95 = 'b000111000;
    x_96 = 'b001000010;
    x_97 = 'b001000000;
    x_98 = 'b000111010;
    x_99 = 'b000110101;
    x_100 = 'b000101001;
    x_101 = 'b000011001;
    x_102 = 'b000110101;
    x_103 = 'b000010110;
    x_104 = 'b001000010;
    x_105 = 'b111111101;
    x_106 = 'b000111010;
    x_107 = 'b000100101;
    x_108 = 'b001001000;
    x_109 = 'b000000101;
    x_110 = 'b001001001;
    x_111 = 'b001001001;
    x_112 = 'b001000000;
    x_113 = 'b001000001;
    x_114 = 'b001001110;
    x_115 = 'b001010010;
    x_116 = 'b001001001;
    x_117 = 'b000111100;
    x_118 = 'b000101010;
    x_119 = 'b000110101;
    x_120 = 'b000111110;
    x_121 = 'b000111110;
    x_122 = 'b001000010;
    x_123 = 'b000101001;
    x_124 = 'b000101110;
    x_125 = 'b000110100;
    x_126 = 'b000100110;
    x_127 = 'b000101101;
    x_128 = 'b000101110;
    x_129 = 'b001001001;
    x_130 = 'b001010010;
    x_131 = 'b001010101;
    x_132 = 'b001001111;
    x_133 = 'b001001100;
    x_134 = 'b000111111;
    x_135 = 'b000110111;
    x_136 = 'b001010001;
    x_137 = 'b001011010;
    x_138 = 'b001011011;
    x_139 = 'b001011111;
    x_140 = 'b001011010;
    x_141 = 'b001000000;
    x_142 = 'b001001101;
    x_143 = 'b001010111;
    x_144 = 'b001011000;
    x_145 = 'b001011101;
    x_146 = 'b001011110;
    x_147 = 'b001011101;
    x_148 = 'b001000011;
    x_149 = 'b000010011;
    x_150 = 'b000010100;
    x_151 = 'b000010110;
    x_152 = 'b000011000;
    x_153 = 'b000011010;
    x_154 = 'b000101101;
    x_155 = 'b000100001;
    x_156 = 'b000011010;
    x_157 = 'b000100011;
    x_158 = 'b000101010;
    x_159 = 'b000111000;
    x_160 = 'b001000010;
    x_161 = 'b001000000;
    x_162 = 'b000111010;
    x_163 = 'b000110101;
    x_164 = 'b000101001;
    x_165 = 'b000011001;
    x_166 = 'b000110101;
    x_167 = 'b000010110;
    x_168 = 'b001000010;
    x_169 = 'b111111101;
    x_170 = 'b000111010;
    x_171 = 'b000100101;
    x_172 = 'b001001000;
    x_173 = 'b000000101;
    x_174 = 'b001001001;
    x_175 = 'b001001001;
    x_176 = 'b001000000;
    x_177 = 'b001000001;
    x_178 = 'b001001110;
    x_179 = 'b001010010;
    x_180 = 'b001001001;
    x_181 = 'b000111100;
    x_182 = 'b000101010;
    x_183 = 'b000110101;
    x_184 = 'b000111110;
    x_185 = 'b000111110;
    x_186 = 'b001000010;
    x_187 = 'b000101001;
    x_188 = 'b000101110;
    x_189 = 'b000110100;
    x_190 = 'b000100110;
    x_191 = 'b000101101;
    x_192 = 'b000101110;
    x_193 = 'b001001001;
    x_194 = 'b001010010;
    x_195 = 'b001010101;
    x_196 = 'b001001111;
    x_197 = 'b001001100;
    x_198 = 'b000111111;
    x_199 = 'b000110111;
    x_200 = 'b001010001;
    x_201 = 'b001011010;
    x_202 = 'b001011011;
    x_203 = 'b001011111;
    x_204 = 'b001011010;
    x_205 = 'b001000000;
    x_206 = 'b001001101;
    x_207 = 'b001010111;
    x_208 = 'b001011000;
    x_209 = 'b001011101;
    x_210 = 'b001011110;
    x_211 = 'b001011101;
    x_212 = 'b001000011;
    x_213 = 'b000010011;
    x_214 = 'b000010100;
    x_215 = 'b000010110;
    x_216 = 'b000011000;
    x_217 = 'b000011010;
    x_218 = 'b000101101;
    x_219 = 'b000100001;
    x_220 = 'b000011010;
    x_221 = 'b000100011;
    x_222 = 'b000101010;
    x_223 = 'b000111000;
    x_224 = 'b001000010;
    x_225 = 'b001000000;
    x_226 = 'b000111010;
    x_227 = 'b000110101;
    x_228 = 'b000101001;
    x_229 = 'b000011001;
    x_230 = 'b000110101;
    x_231 = 'b000010110;
    x_232 = 'b001000010;
    x_233 = 'b111111101;
    x_234 = 'b000111010;
    x_235 = 'b000100101;
    x_236 = 'b001001000;
    x_237 = 'b000000101;
    x_238 = 'b001001001;
    x_239 = 'b001001001;
    x_240 = 'b001000000;
    x_241 = 'b001000001;
    x_242 = 'b001001110;
    x_243 = 'b001010010;
    x_244 = 'b001001001;
    x_245 = 'b000111100;
    x_246 = 'b000101010;
    x_247 = 'b000110101;
    x_248 = 'b000111110;
    x_249 = 'b000111110;
    x_250 = 'b001000010;
    x_251 = 'b000101001;
    x_252 = 'b000101110;
    x_253 = 'b000110100;
    x_254 = 'b000100110;
    x_255 = 'b000101101;

    h_0 = 'b000101110;
    h_1 = 'b001001001;
    h_2 = 'b001010010;
    h_3 = 'b001010101;
    h_4 = 'b001001111;
    h_5 = 'b001001100;
    h_6 = 'b000111111;
    h_7 = 'b000110111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000111111;
    x_1 = 'b001000011;
    x_2 = 'b001000001;
    x_3 = 'b001000000;
    x_4 = 'b000110111;
    x_5 = 'b000101101;
    x_6 = 'b000011110;
    x_7 = 'b000110010;
    x_8 = 'b001000010;
    x_9 = 'b001000001;
    x_10 = 'b001000000;
    x_11 = 'b001000011;
    x_12 = 'b000110100;
    x_13 = 'b000001110;
    x_14 = 'b001000001;
    x_15 = 'b001000010;
    x_16 = 'b001000001;
    x_17 = 'b001000011;
    x_18 = 'b001000001;
    x_19 = 'b000111100;
    x_20 = 'b000011101;
    x_21 = 'b000100001;
    x_22 = 'b000011010;
    x_23 = 'b000010111;
    x_24 = 'b000101100;
    x_25 = 'b000101101;
    x_26 = 'b000100100;
    x_27 = 'b000011100;
    x_28 = 'b000011000;
    x_29 = 'b000111011;
    x_30 = 'b000101011;
    x_31 = 'b000101001;
    x_32 = 'b000110011;
    x_33 = 'b000101110;
    x_34 = 'b000100111;
    x_35 = 'b000100010;
    x_36 = 'b000011001;
    x_37 = 'b000010010;
    x_38 = 'b000110100;
    x_39 = 'b000000010;
    x_40 = 'b000111000;
    x_41 = 'b000000001;
    x_42 = 'b000110110;
    x_43 = 'b000100010;
    x_44 = 'b000111100;
    x_45 = 'b000000100;
    x_46 = 'b000111010;
    x_47 = 'b000110111;
    x_48 = 'b000101011;
    x_49 = 'b000101100;
    x_50 = 'b000111000;
    x_51 = 'b000111011;
    x_52 = 'b000110011;
    x_53 = 'b000101011;
    x_54 = 'b000100010;
    x_55 = 'b000100101;
    x_56 = 'b000110000;
    x_57 = 'b000101110;
    x_58 = 'b000110101;
    x_59 = 'b000100101;
    x_60 = 'b000100110;
    x_61 = 'b000101110;
    x_62 = 'b000100010;
    x_63 = 'b000101110;
    x_64 = 'b000111111;
    x_65 = 'b001000011;
    x_66 = 'b001000001;
    x_67 = 'b001000000;
    x_68 = 'b000110111;
    x_69 = 'b000101101;
    x_70 = 'b000011110;
    x_71 = 'b000110010;
    x_72 = 'b001000010;
    x_73 = 'b001000001;
    x_74 = 'b001000000;
    x_75 = 'b001000011;
    x_76 = 'b000110100;
    x_77 = 'b000001110;
    x_78 = 'b001000001;
    x_79 = 'b001000010;
    x_80 = 'b001000001;
    x_81 = 'b001000011;
    x_82 = 'b001000001;
    x_83 = 'b000111100;
    x_84 = 'b000011101;
    x_85 = 'b000100001;
    x_86 = 'b000011010;
    x_87 = 'b000010111;
    x_88 = 'b000101100;
    x_89 = 'b000101101;
    x_90 = 'b000100100;
    x_91 = 'b000011100;
    x_92 = 'b000011000;
    x_93 = 'b000111011;
    x_94 = 'b000101011;
    x_95 = 'b000101001;
    x_96 = 'b000110011;
    x_97 = 'b000101110;
    x_98 = 'b000100111;
    x_99 = 'b000100010;
    x_100 = 'b000011001;
    x_101 = 'b000010010;
    x_102 = 'b000110100;
    x_103 = 'b000000010;
    x_104 = 'b000111000;
    x_105 = 'b000000001;
    x_106 = 'b000110110;
    x_107 = 'b000100010;
    x_108 = 'b000111100;
    x_109 = 'b000000100;
    x_110 = 'b000111010;
    x_111 = 'b000110111;
    x_112 = 'b000101011;
    x_113 = 'b000101100;
    x_114 = 'b000111000;
    x_115 = 'b000111011;
    x_116 = 'b000110011;
    x_117 = 'b000101011;
    x_118 = 'b000100010;
    x_119 = 'b000100101;
    x_120 = 'b000110000;
    x_121 = 'b000101110;
    x_122 = 'b000110101;
    x_123 = 'b000100101;
    x_124 = 'b000100110;
    x_125 = 'b000101110;
    x_126 = 'b000100010;
    x_127 = 'b000101110;
    x_128 = 'b000111111;
    x_129 = 'b001000011;
    x_130 = 'b001000001;
    x_131 = 'b001000000;
    x_132 = 'b000110111;
    x_133 = 'b000101101;
    x_134 = 'b000011110;
    x_135 = 'b000110010;
    x_136 = 'b001000010;
    x_137 = 'b001000001;
    x_138 = 'b001000000;
    x_139 = 'b001000011;
    x_140 = 'b000110100;
    x_141 = 'b000001110;
    x_142 = 'b001000001;
    x_143 = 'b001000010;
    x_144 = 'b001000001;
    x_145 = 'b001000011;
    x_146 = 'b001000001;
    x_147 = 'b000111100;
    x_148 = 'b000011101;
    x_149 = 'b000100001;
    x_150 = 'b000011010;
    x_151 = 'b000010111;
    x_152 = 'b000101100;
    x_153 = 'b000101101;
    x_154 = 'b000100100;
    x_155 = 'b000011100;
    x_156 = 'b000011000;
    x_157 = 'b000111011;
    x_158 = 'b000101011;
    x_159 = 'b000101001;
    x_160 = 'b000110011;
    x_161 = 'b000101110;
    x_162 = 'b000100111;
    x_163 = 'b000100010;
    x_164 = 'b000011001;
    x_165 = 'b000010010;
    x_166 = 'b000110100;
    x_167 = 'b000000010;
    x_168 = 'b000111000;
    x_169 = 'b000000001;
    x_170 = 'b000110110;
    x_171 = 'b000100010;
    x_172 = 'b000111100;
    x_173 = 'b000000100;
    x_174 = 'b000111010;
    x_175 = 'b000110111;
    x_176 = 'b000101011;
    x_177 = 'b000101100;
    x_178 = 'b000111000;
    x_179 = 'b000111011;
    x_180 = 'b000110011;
    x_181 = 'b000101011;
    x_182 = 'b000100010;
    x_183 = 'b000100101;
    x_184 = 'b000110000;
    x_185 = 'b000101110;
    x_186 = 'b000110101;
    x_187 = 'b000100101;
    x_188 = 'b000100110;
    x_189 = 'b000101110;
    x_190 = 'b000100010;
    x_191 = 'b000101110;
    x_192 = 'b000111111;
    x_193 = 'b001000011;
    x_194 = 'b001000001;
    x_195 = 'b001000000;
    x_196 = 'b000110111;
    x_197 = 'b000101101;
    x_198 = 'b000011110;
    x_199 = 'b000110010;
    x_200 = 'b001000010;
    x_201 = 'b001000001;
    x_202 = 'b001000000;
    x_203 = 'b001000011;
    x_204 = 'b000110100;
    x_205 = 'b000001110;
    x_206 = 'b001000001;
    x_207 = 'b001000010;
    x_208 = 'b001000001;
    x_209 = 'b001000011;
    x_210 = 'b001000001;
    x_211 = 'b000111100;
    x_212 = 'b000011101;
    x_213 = 'b000100001;
    x_214 = 'b000011010;
    x_215 = 'b000010111;
    x_216 = 'b000101100;
    x_217 = 'b000101101;
    x_218 = 'b000100100;
    x_219 = 'b000011100;
    x_220 = 'b000011000;
    x_221 = 'b000111011;
    x_222 = 'b000101011;
    x_223 = 'b000101001;
    x_224 = 'b000110011;
    x_225 = 'b000101110;
    x_226 = 'b000100111;
    x_227 = 'b000100010;
    x_228 = 'b000011001;
    x_229 = 'b000010010;
    x_230 = 'b000110100;
    x_231 = 'b000000010;
    x_232 = 'b000111000;
    x_233 = 'b000000001;
    x_234 = 'b000110110;
    x_235 = 'b000100010;
    x_236 = 'b000111100;
    x_237 = 'b000000100;
    x_238 = 'b000111010;
    x_239 = 'b000110111;
    x_240 = 'b000101011;
    x_241 = 'b000101100;
    x_242 = 'b000111000;
    x_243 = 'b000111011;
    x_244 = 'b000110011;
    x_245 = 'b000101011;
    x_246 = 'b000100010;
    x_247 = 'b000100101;
    x_248 = 'b000110000;
    x_249 = 'b000101110;
    x_250 = 'b000110101;
    x_251 = 'b000100101;
    x_252 = 'b000100110;
    x_253 = 'b000101110;
    x_254 = 'b000100010;
    x_255 = 'b000101110;

    h_0 = 'b000111111;
    h_1 = 'b001000011;
    h_2 = 'b001000001;
    h_3 = 'b001000000;
    h_4 = 'b000110111;
    h_5 = 'b000101101;
    h_6 = 'b000011110;
    h_7 = 'b000110010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000101101;
    x_1 = 'b000101111;
    x_2 = 'b000110100;
    x_3 = 'b000111010;
    x_4 = 'b000110001;
    x_5 = 'b000100100;
    x_6 = 'b000011100;
    x_7 = 'b000011111;
    x_8 = 'b000110001;
    x_9 = 'b000110101;
    x_10 = 'b000111000;
    x_11 = 'b000111100;
    x_12 = 'b000101011;
    x_13 = 'b000010001;
    x_14 = 'b000101110;
    x_15 = 'b000110110;
    x_16 = 'b000110101;
    x_17 = 'b000110110;
    x_18 = 'b000110111;
    x_19 = 'b000110010;
    x_20 = 'b000011100;
    x_21 = 'b000011011;
    x_22 = 'b000011001;
    x_23 = 'b000011111;
    x_24 = 'b000100000;
    x_25 = 'b000100010;
    x_26 = 'b000100110;
    x_27 = 'b000100010;
    x_28 = 'b000100100;
    x_29 = 'b000100001;
    x_30 = 'b000011111;
    x_31 = 'b000101000;
    x_32 = 'b000110001;
    x_33 = 'b000110000;
    x_34 = 'b000101100;
    x_35 = 'b000100101;
    x_36 = 'b000100011;
    x_37 = 'b000011011;
    x_38 = 'b000011100;
    x_39 = 'b000011100;
    x_40 = 'b000110001;
    x_41 = 'b000101101;
    x_42 = 'b000100001;
    x_43 = 'b000001101;
    x_44 = 'b000100010;
    x_45 = 'b000001111;
    x_46 = 'b000100011;
    x_47 = 'b000101001;
    x_48 = 'b000100011;
    x_49 = 'b000100100;
    x_50 = 'b000101100;
    x_51 = 'b000101110;
    x_52 = 'b000100111;
    x_53 = 'b000100100;
    x_54 = 'b000011111;
    x_55 = 'b000011101;
    x_56 = 'b000100111;
    x_57 = 'b000100111;
    x_58 = 'b000101100;
    x_59 = 'b000100001;
    x_60 = 'b000011101;
    x_61 = 'b000100111;
    x_62 = 'b000011010;
    x_63 = 'b000101110;
    x_64 = 'b000101101;
    x_65 = 'b000101111;
    x_66 = 'b000110100;
    x_67 = 'b000111010;
    x_68 = 'b000110001;
    x_69 = 'b000100100;
    x_70 = 'b000011100;
    x_71 = 'b000011111;
    x_72 = 'b000110001;
    x_73 = 'b000110101;
    x_74 = 'b000111000;
    x_75 = 'b000111100;
    x_76 = 'b000101011;
    x_77 = 'b000010001;
    x_78 = 'b000101110;
    x_79 = 'b000110110;
    x_80 = 'b000110101;
    x_81 = 'b000110110;
    x_82 = 'b000110111;
    x_83 = 'b000110010;
    x_84 = 'b000011100;
    x_85 = 'b000011011;
    x_86 = 'b000011001;
    x_87 = 'b000011111;
    x_88 = 'b000100000;
    x_89 = 'b000100010;
    x_90 = 'b000100110;
    x_91 = 'b000100010;
    x_92 = 'b000100100;
    x_93 = 'b000100001;
    x_94 = 'b000011111;
    x_95 = 'b000101000;
    x_96 = 'b000110001;
    x_97 = 'b000110000;
    x_98 = 'b000101100;
    x_99 = 'b000100101;
    x_100 = 'b000100011;
    x_101 = 'b000011011;
    x_102 = 'b000011100;
    x_103 = 'b000011100;
    x_104 = 'b000110001;
    x_105 = 'b000101101;
    x_106 = 'b000100001;
    x_107 = 'b000001101;
    x_108 = 'b000100010;
    x_109 = 'b000001111;
    x_110 = 'b000100011;
    x_111 = 'b000101001;
    x_112 = 'b000100011;
    x_113 = 'b000100100;
    x_114 = 'b000101100;
    x_115 = 'b000101110;
    x_116 = 'b000100111;
    x_117 = 'b000100100;
    x_118 = 'b000011111;
    x_119 = 'b000011101;
    x_120 = 'b000100111;
    x_121 = 'b000100111;
    x_122 = 'b000101100;
    x_123 = 'b000100001;
    x_124 = 'b000011101;
    x_125 = 'b000100111;
    x_126 = 'b000011010;
    x_127 = 'b000101110;
    x_128 = 'b000101101;
    x_129 = 'b000101111;
    x_130 = 'b000110100;
    x_131 = 'b000111010;
    x_132 = 'b000110001;
    x_133 = 'b000100100;
    x_134 = 'b000011100;
    x_135 = 'b000011111;
    x_136 = 'b000110001;
    x_137 = 'b000110101;
    x_138 = 'b000111000;
    x_139 = 'b000111100;
    x_140 = 'b000101011;
    x_141 = 'b000010001;
    x_142 = 'b000101110;
    x_143 = 'b000110110;
    x_144 = 'b000110101;
    x_145 = 'b000110110;
    x_146 = 'b000110111;
    x_147 = 'b000110010;
    x_148 = 'b000011100;
    x_149 = 'b000011011;
    x_150 = 'b000011001;
    x_151 = 'b000011111;
    x_152 = 'b000100000;
    x_153 = 'b000100010;
    x_154 = 'b000100110;
    x_155 = 'b000100010;
    x_156 = 'b000100100;
    x_157 = 'b000100001;
    x_158 = 'b000011111;
    x_159 = 'b000101000;
    x_160 = 'b000110001;
    x_161 = 'b000110000;
    x_162 = 'b000101100;
    x_163 = 'b000100101;
    x_164 = 'b000100011;
    x_165 = 'b000011011;
    x_166 = 'b000011100;
    x_167 = 'b000011100;
    x_168 = 'b000110001;
    x_169 = 'b000101101;
    x_170 = 'b000100001;
    x_171 = 'b000001101;
    x_172 = 'b000100010;
    x_173 = 'b000001111;
    x_174 = 'b000100011;
    x_175 = 'b000101001;
    x_176 = 'b000100011;
    x_177 = 'b000100100;
    x_178 = 'b000101100;
    x_179 = 'b000101110;
    x_180 = 'b000100111;
    x_181 = 'b000100100;
    x_182 = 'b000011111;
    x_183 = 'b000011101;
    x_184 = 'b000100111;
    x_185 = 'b000100111;
    x_186 = 'b000101100;
    x_187 = 'b000100001;
    x_188 = 'b000011101;
    x_189 = 'b000100111;
    x_190 = 'b000011010;
    x_191 = 'b000101110;
    x_192 = 'b000101101;
    x_193 = 'b000101111;
    x_194 = 'b000110100;
    x_195 = 'b000111010;
    x_196 = 'b000110001;
    x_197 = 'b000100100;
    x_198 = 'b000011100;
    x_199 = 'b000011111;
    x_200 = 'b000110001;
    x_201 = 'b000110101;
    x_202 = 'b000111000;
    x_203 = 'b000111100;
    x_204 = 'b000101011;
    x_205 = 'b000010001;
    x_206 = 'b000101110;
    x_207 = 'b000110110;
    x_208 = 'b000110101;
    x_209 = 'b000110110;
    x_210 = 'b000110111;
    x_211 = 'b000110010;
    x_212 = 'b000011100;
    x_213 = 'b000011011;
    x_214 = 'b000011001;
    x_215 = 'b000011111;
    x_216 = 'b000100000;
    x_217 = 'b000100010;
    x_218 = 'b000100110;
    x_219 = 'b000100010;
    x_220 = 'b000100100;
    x_221 = 'b000100001;
    x_222 = 'b000011111;
    x_223 = 'b000101000;
    x_224 = 'b000110001;
    x_225 = 'b000110000;
    x_226 = 'b000101100;
    x_227 = 'b000100101;
    x_228 = 'b000100011;
    x_229 = 'b000011011;
    x_230 = 'b000011100;
    x_231 = 'b000011100;
    x_232 = 'b000110001;
    x_233 = 'b000101101;
    x_234 = 'b000100001;
    x_235 = 'b000001101;
    x_236 = 'b000100010;
    x_237 = 'b000001111;
    x_238 = 'b000100011;
    x_239 = 'b000101001;
    x_240 = 'b000100011;
    x_241 = 'b000100100;
    x_242 = 'b000101100;
    x_243 = 'b000101110;
    x_244 = 'b000100111;
    x_245 = 'b000100100;
    x_246 = 'b000011111;
    x_247 = 'b000011101;
    x_248 = 'b000100111;
    x_249 = 'b000100111;
    x_250 = 'b000101100;
    x_251 = 'b000100001;
    x_252 = 'b000011101;
    x_253 = 'b000100111;
    x_254 = 'b000011010;
    x_255 = 'b000101110;

    h_0 = 'b000101101;
    h_1 = 'b000101111;
    h_2 = 'b000110100;
    h_3 = 'b000111010;
    h_4 = 'b000110001;
    h_5 = 'b000100100;
    h_6 = 'b000011100;
    h_7 = 'b000011111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000011100;
    x_1 = 'b000100110;
    x_2 = 'b000101001;
    x_3 = 'b000110001;
    x_4 = 'b000101100;
    x_5 = 'b000100000;
    x_6 = 'b000011101;
    x_7 = 'b000010100;
    x_8 = 'b000100001;
    x_9 = 'b000100111;
    x_10 = 'b000101010;
    x_11 = 'b000110000;
    x_12 = 'b000100001;
    x_13 = 'b000010000;
    x_14 = 'b000100010;
    x_15 = 'b000101000;
    x_16 = 'b000101000;
    x_17 = 'b000101000;
    x_18 = 'b000100111;
    x_19 = 'b000100010;
    x_20 = 'b000010010;
    x_21 = 'b000011111;
    x_22 = 'b000010101;
    x_23 = 'b000011011;
    x_24 = 'b000010110;
    x_25 = 'b000010111;
    x_26 = 'b000100000;
    x_27 = 'b000011101;
    x_28 = 'b000011111;
    x_29 = 'b000001110;
    x_30 = 'b000011001;
    x_31 = 'b000100001;
    x_32 = 'b000101000;
    x_33 = 'b000100110;
    x_34 = 'b000100101;
    x_35 = 'b000011011;
    x_36 = 'b000011010;
    x_37 = 'b000010100;
    x_38 = 'b000001100;
    x_39 = 'b000001110;
    x_40 = 'b000000110;
    x_41 = 'b000001100;
    x_42 = 'b000000100;
    x_43 = 'b111111011;
    x_44 = 'b000010001;
    x_45 = 'b000000100;
    x_46 = 'b000011101;
    x_47 = 'b000100100;
    x_48 = 'b000011101;
    x_49 = 'b000011111;
    x_50 = 'b000100101;
    x_51 = 'b000100101;
    x_52 = 'b000011101;
    x_53 = 'b000011010;
    x_54 = 'b000010011;
    x_55 = 'b000011010;
    x_56 = 'b000100100;
    x_57 = 'b000100011;
    x_58 = 'b000100101;
    x_59 = 'b000011010;
    x_60 = 'b000011000;
    x_61 = 'b000100001;
    x_62 = 'b000010010;
    x_63 = 'b000101010;
    x_64 = 'b000011100;
    x_65 = 'b000100110;
    x_66 = 'b000101001;
    x_67 = 'b000110001;
    x_68 = 'b000101100;
    x_69 = 'b000100000;
    x_70 = 'b000011101;
    x_71 = 'b000010100;
    x_72 = 'b000100001;
    x_73 = 'b000100111;
    x_74 = 'b000101010;
    x_75 = 'b000110000;
    x_76 = 'b000100001;
    x_77 = 'b000010000;
    x_78 = 'b000100010;
    x_79 = 'b000101000;
    x_80 = 'b000101000;
    x_81 = 'b000101000;
    x_82 = 'b000100111;
    x_83 = 'b000100010;
    x_84 = 'b000010010;
    x_85 = 'b000011111;
    x_86 = 'b000010101;
    x_87 = 'b000011011;
    x_88 = 'b000010110;
    x_89 = 'b000010111;
    x_90 = 'b000100000;
    x_91 = 'b000011101;
    x_92 = 'b000011111;
    x_93 = 'b000001110;
    x_94 = 'b000011001;
    x_95 = 'b000100001;
    x_96 = 'b000101000;
    x_97 = 'b000100110;
    x_98 = 'b000100101;
    x_99 = 'b000011011;
    x_100 = 'b000011010;
    x_101 = 'b000010100;
    x_102 = 'b000001100;
    x_103 = 'b000001110;
    x_104 = 'b000000110;
    x_105 = 'b000001100;
    x_106 = 'b000000100;
    x_107 = 'b111111011;
    x_108 = 'b000010001;
    x_109 = 'b000000100;
    x_110 = 'b000011101;
    x_111 = 'b000100100;
    x_112 = 'b000011101;
    x_113 = 'b000011111;
    x_114 = 'b000100101;
    x_115 = 'b000100101;
    x_116 = 'b000011101;
    x_117 = 'b000011010;
    x_118 = 'b000010011;
    x_119 = 'b000011010;
    x_120 = 'b000100100;
    x_121 = 'b000100011;
    x_122 = 'b000100101;
    x_123 = 'b000011010;
    x_124 = 'b000011000;
    x_125 = 'b000100001;
    x_126 = 'b000010010;
    x_127 = 'b000101010;
    x_128 = 'b000011100;
    x_129 = 'b000100110;
    x_130 = 'b000101001;
    x_131 = 'b000110001;
    x_132 = 'b000101100;
    x_133 = 'b000100000;
    x_134 = 'b000011101;
    x_135 = 'b000010100;
    x_136 = 'b000100001;
    x_137 = 'b000100111;
    x_138 = 'b000101010;
    x_139 = 'b000110000;
    x_140 = 'b000100001;
    x_141 = 'b000010000;
    x_142 = 'b000100010;
    x_143 = 'b000101000;
    x_144 = 'b000101000;
    x_145 = 'b000101000;
    x_146 = 'b000100111;
    x_147 = 'b000100010;
    x_148 = 'b000010010;
    x_149 = 'b000011111;
    x_150 = 'b000010101;
    x_151 = 'b000011011;
    x_152 = 'b000010110;
    x_153 = 'b000010111;
    x_154 = 'b000100000;
    x_155 = 'b000011101;
    x_156 = 'b000011111;
    x_157 = 'b000001110;
    x_158 = 'b000011001;
    x_159 = 'b000100001;
    x_160 = 'b000101000;
    x_161 = 'b000100110;
    x_162 = 'b000100101;
    x_163 = 'b000011011;
    x_164 = 'b000011010;
    x_165 = 'b000010100;
    x_166 = 'b000001100;
    x_167 = 'b000001110;
    x_168 = 'b000000110;
    x_169 = 'b000001100;
    x_170 = 'b000000100;
    x_171 = 'b111111011;
    x_172 = 'b000010001;
    x_173 = 'b000000100;
    x_174 = 'b000011101;
    x_175 = 'b000100100;
    x_176 = 'b000011101;
    x_177 = 'b000011111;
    x_178 = 'b000100101;
    x_179 = 'b000100101;
    x_180 = 'b000011101;
    x_181 = 'b000011010;
    x_182 = 'b000010011;
    x_183 = 'b000011010;
    x_184 = 'b000100100;
    x_185 = 'b000100011;
    x_186 = 'b000100101;
    x_187 = 'b000011010;
    x_188 = 'b000011000;
    x_189 = 'b000100001;
    x_190 = 'b000010010;
    x_191 = 'b000101010;
    x_192 = 'b000011100;
    x_193 = 'b000100110;
    x_194 = 'b000101001;
    x_195 = 'b000110001;
    x_196 = 'b000101100;
    x_197 = 'b000100000;
    x_198 = 'b000011101;
    x_199 = 'b000010100;
    x_200 = 'b000100001;
    x_201 = 'b000100111;
    x_202 = 'b000101010;
    x_203 = 'b000110000;
    x_204 = 'b000100001;
    x_205 = 'b000010000;
    x_206 = 'b000100010;
    x_207 = 'b000101000;
    x_208 = 'b000101000;
    x_209 = 'b000101000;
    x_210 = 'b000100111;
    x_211 = 'b000100010;
    x_212 = 'b000010010;
    x_213 = 'b000011111;
    x_214 = 'b000010101;
    x_215 = 'b000011011;
    x_216 = 'b000010110;
    x_217 = 'b000010111;
    x_218 = 'b000100000;
    x_219 = 'b000011101;
    x_220 = 'b000011111;
    x_221 = 'b000001110;
    x_222 = 'b000011001;
    x_223 = 'b000100001;
    x_224 = 'b000101000;
    x_225 = 'b000100110;
    x_226 = 'b000100101;
    x_227 = 'b000011011;
    x_228 = 'b000011010;
    x_229 = 'b000010100;
    x_230 = 'b000001100;
    x_231 = 'b000001110;
    x_232 = 'b000000110;
    x_233 = 'b000001100;
    x_234 = 'b000000100;
    x_235 = 'b111111011;
    x_236 = 'b000010001;
    x_237 = 'b000000100;
    x_238 = 'b000011101;
    x_239 = 'b000100100;
    x_240 = 'b000011101;
    x_241 = 'b000011111;
    x_242 = 'b000100101;
    x_243 = 'b000100101;
    x_244 = 'b000011101;
    x_245 = 'b000011010;
    x_246 = 'b000010011;
    x_247 = 'b000011010;
    x_248 = 'b000100100;
    x_249 = 'b000100011;
    x_250 = 'b000100101;
    x_251 = 'b000011010;
    x_252 = 'b000011000;
    x_253 = 'b000100001;
    x_254 = 'b000010010;
    x_255 = 'b000101010;

    h_0 = 'b000011100;
    h_1 = 'b000100110;
    h_2 = 'b000101001;
    h_3 = 'b000110001;
    h_4 = 'b000101100;
    h_5 = 'b000100000;
    h_6 = 'b000011101;
    h_7 = 'b000010100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000010011;
    x_1 = 'b000011111;
    x_2 = 'b000100100;
    x_3 = 'b000101100;
    x_4 = 'b000100101;
    x_5 = 'b000010111;
    x_6 = 'b000010101;
    x_7 = 'b000001011;
    x_8 = 'b000011101;
    x_9 = 'b000100101;
    x_10 = 'b000101000;
    x_11 = 'b000101111;
    x_12 = 'b000011110;
    x_13 = 'b000001101;
    x_14 = 'b000100000;
    x_15 = 'b000100111;
    x_16 = 'b000100111;
    x_17 = 'b000101001;
    x_18 = 'b000100111;
    x_19 = 'b000100100;
    x_20 = 'b000010101;
    x_21 = 'b000010011;
    x_22 = 'b000010000;
    x_23 = 'b000010010;
    x_24 = 'b000010010;
    x_25 = 'b000010011;
    x_26 = 'b000011010;
    x_27 = 'b000010011;
    x_28 = 'b000010011;
    x_29 = 'b000001100;
    x_30 = 'b000011101;
    x_31 = 'b000011110;
    x_32 = 'b000101000;
    x_33 = 'b000100101;
    x_34 = 'b000100001;
    x_35 = 'b000011010;
    x_36 = 'b000010100;
    x_37 = 'b000001101;
    x_38 = 'b000001011;
    x_39 = 'b000001001;
    x_40 = 'b000010001;
    x_41 = 'b000000101;
    x_42 = 'b000010101;
    x_43 = 'b000011011;
    x_44 = 'b000011010;
    x_45 = 'b000001010;
    x_46 = 'b000011001;
    x_47 = 'b000011101;
    x_48 = 'b000010101;
    x_49 = 'b000011100;
    x_50 = 'b000100101;
    x_51 = 'b000101001;
    x_52 = 'b000100100;
    x_53 = 'b000100101;
    x_54 = 'b000011011;
    x_55 = 'b000010001;
    x_56 = 'b000011100;
    x_57 = 'b000011111;
    x_58 = 'b000100111;
    x_59 = 'b000011001;
    x_60 = 'b000010100;
    x_61 = 'b000011011;
    x_62 = 'b000001011;
    x_63 = 'b000100011;
    x_64 = 'b000010011;
    x_65 = 'b000011111;
    x_66 = 'b000100100;
    x_67 = 'b000101100;
    x_68 = 'b000100101;
    x_69 = 'b000010111;
    x_70 = 'b000010101;
    x_71 = 'b000001011;
    x_72 = 'b000011101;
    x_73 = 'b000100101;
    x_74 = 'b000101000;
    x_75 = 'b000101111;
    x_76 = 'b000011110;
    x_77 = 'b000001101;
    x_78 = 'b000100000;
    x_79 = 'b000100111;
    x_80 = 'b000100111;
    x_81 = 'b000101001;
    x_82 = 'b000100111;
    x_83 = 'b000100100;
    x_84 = 'b000010101;
    x_85 = 'b000010011;
    x_86 = 'b000010000;
    x_87 = 'b000010010;
    x_88 = 'b000010010;
    x_89 = 'b000010011;
    x_90 = 'b000011010;
    x_91 = 'b000010011;
    x_92 = 'b000010011;
    x_93 = 'b000001100;
    x_94 = 'b000011101;
    x_95 = 'b000011110;
    x_96 = 'b000101000;
    x_97 = 'b000100101;
    x_98 = 'b000100001;
    x_99 = 'b000011010;
    x_100 = 'b000010100;
    x_101 = 'b000001101;
    x_102 = 'b000001011;
    x_103 = 'b000001001;
    x_104 = 'b000010001;
    x_105 = 'b000000101;
    x_106 = 'b000010101;
    x_107 = 'b000011011;
    x_108 = 'b000011010;
    x_109 = 'b000001010;
    x_110 = 'b000011001;
    x_111 = 'b000011101;
    x_112 = 'b000010101;
    x_113 = 'b000011100;
    x_114 = 'b000100101;
    x_115 = 'b000101001;
    x_116 = 'b000100100;
    x_117 = 'b000100101;
    x_118 = 'b000011011;
    x_119 = 'b000010001;
    x_120 = 'b000011100;
    x_121 = 'b000011111;
    x_122 = 'b000100111;
    x_123 = 'b000011001;
    x_124 = 'b000010100;
    x_125 = 'b000011011;
    x_126 = 'b000001011;
    x_127 = 'b000100011;
    x_128 = 'b000010011;
    x_129 = 'b000011111;
    x_130 = 'b000100100;
    x_131 = 'b000101100;
    x_132 = 'b000100101;
    x_133 = 'b000010111;
    x_134 = 'b000010101;
    x_135 = 'b000001011;
    x_136 = 'b000011101;
    x_137 = 'b000100101;
    x_138 = 'b000101000;
    x_139 = 'b000101111;
    x_140 = 'b000011110;
    x_141 = 'b000001101;
    x_142 = 'b000100000;
    x_143 = 'b000100111;
    x_144 = 'b000100111;
    x_145 = 'b000101001;
    x_146 = 'b000100111;
    x_147 = 'b000100100;
    x_148 = 'b000010101;
    x_149 = 'b000010011;
    x_150 = 'b000010000;
    x_151 = 'b000010010;
    x_152 = 'b000010010;
    x_153 = 'b000010011;
    x_154 = 'b000011010;
    x_155 = 'b000010011;
    x_156 = 'b000010011;
    x_157 = 'b000001100;
    x_158 = 'b000011101;
    x_159 = 'b000011110;
    x_160 = 'b000101000;
    x_161 = 'b000100101;
    x_162 = 'b000100001;
    x_163 = 'b000011010;
    x_164 = 'b000010100;
    x_165 = 'b000001101;
    x_166 = 'b000001011;
    x_167 = 'b000001001;
    x_168 = 'b000010001;
    x_169 = 'b000000101;
    x_170 = 'b000010101;
    x_171 = 'b000011011;
    x_172 = 'b000011010;
    x_173 = 'b000001010;
    x_174 = 'b000011001;
    x_175 = 'b000011101;
    x_176 = 'b000010101;
    x_177 = 'b000011100;
    x_178 = 'b000100101;
    x_179 = 'b000101001;
    x_180 = 'b000100100;
    x_181 = 'b000100101;
    x_182 = 'b000011011;
    x_183 = 'b000010001;
    x_184 = 'b000011100;
    x_185 = 'b000011111;
    x_186 = 'b000100111;
    x_187 = 'b000011001;
    x_188 = 'b000010100;
    x_189 = 'b000011011;
    x_190 = 'b000001011;
    x_191 = 'b000100011;
    x_192 = 'b000010011;
    x_193 = 'b000011111;
    x_194 = 'b000100100;
    x_195 = 'b000101100;
    x_196 = 'b000100101;
    x_197 = 'b000010111;
    x_198 = 'b000010101;
    x_199 = 'b000001011;
    x_200 = 'b000011101;
    x_201 = 'b000100101;
    x_202 = 'b000101000;
    x_203 = 'b000101111;
    x_204 = 'b000011110;
    x_205 = 'b000001101;
    x_206 = 'b000100000;
    x_207 = 'b000100111;
    x_208 = 'b000100111;
    x_209 = 'b000101001;
    x_210 = 'b000100111;
    x_211 = 'b000100100;
    x_212 = 'b000010101;
    x_213 = 'b000010011;
    x_214 = 'b000010000;
    x_215 = 'b000010010;
    x_216 = 'b000010010;
    x_217 = 'b000010011;
    x_218 = 'b000011010;
    x_219 = 'b000010011;
    x_220 = 'b000010011;
    x_221 = 'b000001100;
    x_222 = 'b000011101;
    x_223 = 'b000011110;
    x_224 = 'b000101000;
    x_225 = 'b000100101;
    x_226 = 'b000100001;
    x_227 = 'b000011010;
    x_228 = 'b000010100;
    x_229 = 'b000001101;
    x_230 = 'b000001011;
    x_231 = 'b000001001;
    x_232 = 'b000010001;
    x_233 = 'b000000101;
    x_234 = 'b000010101;
    x_235 = 'b000011011;
    x_236 = 'b000011010;
    x_237 = 'b000001010;
    x_238 = 'b000011001;
    x_239 = 'b000011101;
    x_240 = 'b000010101;
    x_241 = 'b000011100;
    x_242 = 'b000100101;
    x_243 = 'b000101001;
    x_244 = 'b000100100;
    x_245 = 'b000100101;
    x_246 = 'b000011011;
    x_247 = 'b000010001;
    x_248 = 'b000011100;
    x_249 = 'b000011111;
    x_250 = 'b000100111;
    x_251 = 'b000011001;
    x_252 = 'b000010100;
    x_253 = 'b000011011;
    x_254 = 'b000001011;
    x_255 = 'b000100011;

    h_0 = 'b000010011;
    h_1 = 'b000011111;
    h_2 = 'b000100100;
    h_3 = 'b000101100;
    h_4 = 'b000100101;
    h_5 = 'b000010111;
    h_6 = 'b000010101;
    h_7 = 'b000001011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000011001;
    x_1 = 'b000100101;
    x_2 = 'b000101100;
    x_3 = 'b000110101;
    x_4 = 'b000101111;
    x_5 = 'b000100010;
    x_6 = 'b000011100;
    x_7 = 'b000000110;
    x_8 = 'b000100000;
    x_9 = 'b000101011;
    x_10 = 'b000110001;
    x_11 = 'b000111010;
    x_12 = 'b000101111;
    x_13 = 'b000011100;
    x_14 = 'b000010011;
    x_15 = 'b000100101;
    x_16 = 'b000101000;
    x_17 = 'b000101010;
    x_18 = 'b000101110;
    x_19 = 'b000110010;
    x_20 = 'b000101001;
    x_21 = 'b000010001;
    x_22 = 'b000001111;
    x_23 = 'b000001111;
    x_24 = 'b000010110;
    x_25 = 'b000010111;
    x_26 = 'b000011101;
    x_27 = 'b000010110;
    x_28 = 'b000010010;
    x_29 = 'b000010001;
    x_30 = 'b000100100;
    x_31 = 'b000100011;
    x_32 = 'b000101010;
    x_33 = 'b000101010;
    x_34 = 'b000100110;
    x_35 = 'b000100000;
    x_36 = 'b000011101;
    x_37 = 'b000010100;
    x_38 = 'b000010011;
    x_39 = 'b000010011;
    x_40 = 'b000100000;
    x_41 = 'b000010011;
    x_42 = 'b000010101;
    x_43 = 'b001001010;
    x_44 = 'b000011001;
    x_45 = 'b000100001;
    x_46 = 'b000010011;
    x_47 = 'b000010101;
    x_48 = 'b000001101;
    x_49 = 'b000010100;
    x_50 = 'b000100011;
    x_51 = 'b000101101;
    x_52 = 'b000101111;
    x_53 = 'b000110011;
    x_54 = 'b000101111;
    x_55 = 'b000001001;
    x_56 = 'b000010101;
    x_57 = 'b000011011;
    x_58 = 'b000101101;
    x_59 = 'b000100000;
    x_60 = 'b000001110;
    x_61 = 'b000010100;
    x_62 = 'b000000111;
    x_63 = 'b000011000;
    x_64 = 'b000011001;
    x_65 = 'b000100101;
    x_66 = 'b000101100;
    x_67 = 'b000110101;
    x_68 = 'b000101111;
    x_69 = 'b000100010;
    x_70 = 'b000011100;
    x_71 = 'b000000110;
    x_72 = 'b000100000;
    x_73 = 'b000101011;
    x_74 = 'b000110001;
    x_75 = 'b000111010;
    x_76 = 'b000101111;
    x_77 = 'b000011100;
    x_78 = 'b000010011;
    x_79 = 'b000100101;
    x_80 = 'b000101000;
    x_81 = 'b000101010;
    x_82 = 'b000101110;
    x_83 = 'b000110010;
    x_84 = 'b000101001;
    x_85 = 'b000010001;
    x_86 = 'b000001111;
    x_87 = 'b000001111;
    x_88 = 'b000010110;
    x_89 = 'b000010111;
    x_90 = 'b000011101;
    x_91 = 'b000010110;
    x_92 = 'b000010010;
    x_93 = 'b000010001;
    x_94 = 'b000100100;
    x_95 = 'b000100011;
    x_96 = 'b000101010;
    x_97 = 'b000101010;
    x_98 = 'b000100110;
    x_99 = 'b000100000;
    x_100 = 'b000011101;
    x_101 = 'b000010100;
    x_102 = 'b000010011;
    x_103 = 'b000010011;
    x_104 = 'b000100000;
    x_105 = 'b000010011;
    x_106 = 'b000010101;
    x_107 = 'b001001010;
    x_108 = 'b000011001;
    x_109 = 'b000100001;
    x_110 = 'b000010011;
    x_111 = 'b000010101;
    x_112 = 'b000001101;
    x_113 = 'b000010100;
    x_114 = 'b000100011;
    x_115 = 'b000101101;
    x_116 = 'b000101111;
    x_117 = 'b000110011;
    x_118 = 'b000101111;
    x_119 = 'b000001001;
    x_120 = 'b000010101;
    x_121 = 'b000011011;
    x_122 = 'b000101101;
    x_123 = 'b000100000;
    x_124 = 'b000001110;
    x_125 = 'b000010100;
    x_126 = 'b000000111;
    x_127 = 'b000011000;
    x_128 = 'b000011001;
    x_129 = 'b000100101;
    x_130 = 'b000101100;
    x_131 = 'b000110101;
    x_132 = 'b000101111;
    x_133 = 'b000100010;
    x_134 = 'b000011100;
    x_135 = 'b000000110;
    x_136 = 'b000100000;
    x_137 = 'b000101011;
    x_138 = 'b000110001;
    x_139 = 'b000111010;
    x_140 = 'b000101111;
    x_141 = 'b000011100;
    x_142 = 'b000010011;
    x_143 = 'b000100101;
    x_144 = 'b000101000;
    x_145 = 'b000101010;
    x_146 = 'b000101110;
    x_147 = 'b000110010;
    x_148 = 'b000101001;
    x_149 = 'b000010001;
    x_150 = 'b000001111;
    x_151 = 'b000001111;
    x_152 = 'b000010110;
    x_153 = 'b000010111;
    x_154 = 'b000011101;
    x_155 = 'b000010110;
    x_156 = 'b000010010;
    x_157 = 'b000010001;
    x_158 = 'b000100100;
    x_159 = 'b000100011;
    x_160 = 'b000101010;
    x_161 = 'b000101010;
    x_162 = 'b000100110;
    x_163 = 'b000100000;
    x_164 = 'b000011101;
    x_165 = 'b000010100;
    x_166 = 'b000010011;
    x_167 = 'b000010011;
    x_168 = 'b000100000;
    x_169 = 'b000010011;
    x_170 = 'b000010101;
    x_171 = 'b001001010;
    x_172 = 'b000011001;
    x_173 = 'b000100001;
    x_174 = 'b000010011;
    x_175 = 'b000010101;
    x_176 = 'b000001101;
    x_177 = 'b000010100;
    x_178 = 'b000100011;
    x_179 = 'b000101101;
    x_180 = 'b000101111;
    x_181 = 'b000110011;
    x_182 = 'b000101111;
    x_183 = 'b000001001;
    x_184 = 'b000010101;
    x_185 = 'b000011011;
    x_186 = 'b000101101;
    x_187 = 'b000100000;
    x_188 = 'b000001110;
    x_189 = 'b000010100;
    x_190 = 'b000000111;
    x_191 = 'b000011000;
    x_192 = 'b000011001;
    x_193 = 'b000100101;
    x_194 = 'b000101100;
    x_195 = 'b000110101;
    x_196 = 'b000101111;
    x_197 = 'b000100010;
    x_198 = 'b000011100;
    x_199 = 'b000000110;
    x_200 = 'b000100000;
    x_201 = 'b000101011;
    x_202 = 'b000110001;
    x_203 = 'b000111010;
    x_204 = 'b000101111;
    x_205 = 'b000011100;
    x_206 = 'b000010011;
    x_207 = 'b000100101;
    x_208 = 'b000101000;
    x_209 = 'b000101010;
    x_210 = 'b000101110;
    x_211 = 'b000110010;
    x_212 = 'b000101001;
    x_213 = 'b000010001;
    x_214 = 'b000001111;
    x_215 = 'b000001111;
    x_216 = 'b000010110;
    x_217 = 'b000010111;
    x_218 = 'b000011101;
    x_219 = 'b000010110;
    x_220 = 'b000010010;
    x_221 = 'b000010001;
    x_222 = 'b000100100;
    x_223 = 'b000100011;
    x_224 = 'b000101010;
    x_225 = 'b000101010;
    x_226 = 'b000100110;
    x_227 = 'b000100000;
    x_228 = 'b000011101;
    x_229 = 'b000010100;
    x_230 = 'b000010011;
    x_231 = 'b000010011;
    x_232 = 'b000100000;
    x_233 = 'b000010011;
    x_234 = 'b000010101;
    x_235 = 'b001001010;
    x_236 = 'b000011001;
    x_237 = 'b000100001;
    x_238 = 'b000010011;
    x_239 = 'b000010101;
    x_240 = 'b000001101;
    x_241 = 'b000010100;
    x_242 = 'b000100011;
    x_243 = 'b000101101;
    x_244 = 'b000101111;
    x_245 = 'b000110011;
    x_246 = 'b000101111;
    x_247 = 'b000001001;
    x_248 = 'b000010101;
    x_249 = 'b000011011;
    x_250 = 'b000101101;
    x_251 = 'b000100000;
    x_252 = 'b000001110;
    x_253 = 'b000010100;
    x_254 = 'b000000111;
    x_255 = 'b000011000;

    h_0 = 'b000011001;
    h_1 = 'b000100101;
    h_2 = 'b000101100;
    h_3 = 'b000110101;
    h_4 = 'b000101111;
    h_5 = 'b000100010;
    h_6 = 'b000011100;
    h_7 = 'b000000110;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000011001;
    x_1 = 'b000100011;
    x_2 = 'b000101001;
    x_3 = 'b000110101;
    x_4 = 'b000110001;
    x_5 = 'b000100111;
    x_6 = 'b000100110;
    x_7 = 'b000001001;
    x_8 = 'b000011100;
    x_9 = 'b000100101;
    x_10 = 'b000101110;
    x_11 = 'b000111010;
    x_12 = 'b000110011;
    x_13 = 'b000100111;
    x_14 = 'b000010011;
    x_15 = 'b000100000;
    x_16 = 'b000100010;
    x_17 = 'b000100110;
    x_18 = 'b000101110;
    x_19 = 'b000110100;
    x_20 = 'b000110000;
    x_21 = 'b000010110;
    x_22 = 'b000010010;
    x_23 = 'b000010101;
    x_24 = 'b000010110;
    x_25 = 'b000011000;
    x_26 = 'b000100001;
    x_27 = 'b000011011;
    x_28 = 'b000011000;
    x_29 = 'b000010001;
    x_30 = 'b000100001;
    x_31 = 'b000100110;
    x_32 = 'b000101011;
    x_33 = 'b000101001;
    x_34 = 'b000100111;
    x_35 = 'b000100001;
    x_36 = 'b000100011;
    x_37 = 'b000011100;
    x_38 = 'b000001101;
    x_39 = 'b000011000;
    x_40 = 'b000011000;
    x_41 = 'b000011001;
    x_42 = 'b000001110;
    x_43 = 'b000101010;
    x_44 = 'b000001110;
    x_45 = 'b000100100;
    x_46 = 'b000001101;
    x_47 = 'b000010010;
    x_48 = 'b000001011;
    x_49 = 'b000010011;
    x_50 = 'b000100001;
    x_51 = 'b000101100;
    x_52 = 'b000101011;
    x_53 = 'b000110001;
    x_54 = 'b000101010;
    x_55 = 'b000001001;
    x_56 = 'b000010100;
    x_57 = 'b000011010;
    x_58 = 'b000101000;
    x_59 = 'b000010111;
    x_60 = 'b000001001;
    x_61 = 'b000001110;
    x_62 = 'b000000011;
    x_63 = 'b000001100;
    x_64 = 'b000011001;
    x_65 = 'b000100011;
    x_66 = 'b000101001;
    x_67 = 'b000110101;
    x_68 = 'b000110001;
    x_69 = 'b000100111;
    x_70 = 'b000100110;
    x_71 = 'b000001001;
    x_72 = 'b000011100;
    x_73 = 'b000100101;
    x_74 = 'b000101110;
    x_75 = 'b000111010;
    x_76 = 'b000110011;
    x_77 = 'b000100111;
    x_78 = 'b000010011;
    x_79 = 'b000100000;
    x_80 = 'b000100010;
    x_81 = 'b000100110;
    x_82 = 'b000101110;
    x_83 = 'b000110100;
    x_84 = 'b000110000;
    x_85 = 'b000010110;
    x_86 = 'b000010010;
    x_87 = 'b000010101;
    x_88 = 'b000010110;
    x_89 = 'b000011000;
    x_90 = 'b000100001;
    x_91 = 'b000011011;
    x_92 = 'b000011000;
    x_93 = 'b000010001;
    x_94 = 'b000100001;
    x_95 = 'b000100110;
    x_96 = 'b000101011;
    x_97 = 'b000101001;
    x_98 = 'b000100111;
    x_99 = 'b000100001;
    x_100 = 'b000100011;
    x_101 = 'b000011100;
    x_102 = 'b000001101;
    x_103 = 'b000011000;
    x_104 = 'b000011000;
    x_105 = 'b000011001;
    x_106 = 'b000001110;
    x_107 = 'b000101010;
    x_108 = 'b000001110;
    x_109 = 'b000100100;
    x_110 = 'b000001101;
    x_111 = 'b000010010;
    x_112 = 'b000001011;
    x_113 = 'b000010011;
    x_114 = 'b000100001;
    x_115 = 'b000101100;
    x_116 = 'b000101011;
    x_117 = 'b000110001;
    x_118 = 'b000101010;
    x_119 = 'b000001001;
    x_120 = 'b000010100;
    x_121 = 'b000011010;
    x_122 = 'b000101000;
    x_123 = 'b000010111;
    x_124 = 'b000001001;
    x_125 = 'b000001110;
    x_126 = 'b000000011;
    x_127 = 'b000001100;
    x_128 = 'b000011001;
    x_129 = 'b000100011;
    x_130 = 'b000101001;
    x_131 = 'b000110101;
    x_132 = 'b000110001;
    x_133 = 'b000100111;
    x_134 = 'b000100110;
    x_135 = 'b000001001;
    x_136 = 'b000011100;
    x_137 = 'b000100101;
    x_138 = 'b000101110;
    x_139 = 'b000111010;
    x_140 = 'b000110011;
    x_141 = 'b000100111;
    x_142 = 'b000010011;
    x_143 = 'b000100000;
    x_144 = 'b000100010;
    x_145 = 'b000100110;
    x_146 = 'b000101110;
    x_147 = 'b000110100;
    x_148 = 'b000110000;
    x_149 = 'b000010110;
    x_150 = 'b000010010;
    x_151 = 'b000010101;
    x_152 = 'b000010110;
    x_153 = 'b000011000;
    x_154 = 'b000100001;
    x_155 = 'b000011011;
    x_156 = 'b000011000;
    x_157 = 'b000010001;
    x_158 = 'b000100001;
    x_159 = 'b000100110;
    x_160 = 'b000101011;
    x_161 = 'b000101001;
    x_162 = 'b000100111;
    x_163 = 'b000100001;
    x_164 = 'b000100011;
    x_165 = 'b000011100;
    x_166 = 'b000001101;
    x_167 = 'b000011000;
    x_168 = 'b000011000;
    x_169 = 'b000011001;
    x_170 = 'b000001110;
    x_171 = 'b000101010;
    x_172 = 'b000001110;
    x_173 = 'b000100100;
    x_174 = 'b000001101;
    x_175 = 'b000010010;
    x_176 = 'b000001011;
    x_177 = 'b000010011;
    x_178 = 'b000100001;
    x_179 = 'b000101100;
    x_180 = 'b000101011;
    x_181 = 'b000110001;
    x_182 = 'b000101010;
    x_183 = 'b000001001;
    x_184 = 'b000010100;
    x_185 = 'b000011010;
    x_186 = 'b000101000;
    x_187 = 'b000010111;
    x_188 = 'b000001001;
    x_189 = 'b000001110;
    x_190 = 'b000000011;
    x_191 = 'b000001100;
    x_192 = 'b000011001;
    x_193 = 'b000100011;
    x_194 = 'b000101001;
    x_195 = 'b000110101;
    x_196 = 'b000110001;
    x_197 = 'b000100111;
    x_198 = 'b000100110;
    x_199 = 'b000001001;
    x_200 = 'b000011100;
    x_201 = 'b000100101;
    x_202 = 'b000101110;
    x_203 = 'b000111010;
    x_204 = 'b000110011;
    x_205 = 'b000100111;
    x_206 = 'b000010011;
    x_207 = 'b000100000;
    x_208 = 'b000100010;
    x_209 = 'b000100110;
    x_210 = 'b000101110;
    x_211 = 'b000110100;
    x_212 = 'b000110000;
    x_213 = 'b000010110;
    x_214 = 'b000010010;
    x_215 = 'b000010101;
    x_216 = 'b000010110;
    x_217 = 'b000011000;
    x_218 = 'b000100001;
    x_219 = 'b000011011;
    x_220 = 'b000011000;
    x_221 = 'b000010001;
    x_222 = 'b000100001;
    x_223 = 'b000100110;
    x_224 = 'b000101011;
    x_225 = 'b000101001;
    x_226 = 'b000100111;
    x_227 = 'b000100001;
    x_228 = 'b000100011;
    x_229 = 'b000011100;
    x_230 = 'b000001101;
    x_231 = 'b000011000;
    x_232 = 'b000011000;
    x_233 = 'b000011001;
    x_234 = 'b000001110;
    x_235 = 'b000101010;
    x_236 = 'b000001110;
    x_237 = 'b000100100;
    x_238 = 'b000001101;
    x_239 = 'b000010010;
    x_240 = 'b000001011;
    x_241 = 'b000010011;
    x_242 = 'b000100001;
    x_243 = 'b000101100;
    x_244 = 'b000101011;
    x_245 = 'b000110001;
    x_246 = 'b000101010;
    x_247 = 'b000001001;
    x_248 = 'b000010100;
    x_249 = 'b000011010;
    x_250 = 'b000101000;
    x_251 = 'b000010111;
    x_252 = 'b000001001;
    x_253 = 'b000001110;
    x_254 = 'b000000011;
    x_255 = 'b000001100;

    h_0 = 'b000011001;
    h_1 = 'b000100011;
    h_2 = 'b000101001;
    h_3 = 'b000110101;
    h_4 = 'b000110001;
    h_5 = 'b000100111;
    h_6 = 'b000100110;
    h_7 = 'b000001001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000010111;
    x_1 = 'b000011110;
    x_2 = 'b000100110;
    x_3 = 'b000101111;
    x_4 = 'b000101011;
    x_5 = 'b000100100;
    x_6 = 'b000100110;
    x_7 = 'b000000110;
    x_8 = 'b000010101;
    x_9 = 'b000011101;
    x_10 = 'b000100101;
    x_11 = 'b000110100;
    x_12 = 'b000101100;
    x_13 = 'b000101001;
    x_14 = 'b000001110;
    x_15 = 'b000011000;
    x_16 = 'b000011011;
    x_17 = 'b000100001;
    x_18 = 'b000100111;
    x_19 = 'b000101100;
    x_20 = 'b000101000;
    x_21 = 'b000011011;
    x_22 = 'b000010011;
    x_23 = 'b000010110;
    x_24 = 'b000011001;
    x_25 = 'b000011011;
    x_26 = 'b000100001;
    x_27 = 'b000011010;
    x_28 = 'b000010010;
    x_29 = 'b000010011;
    x_30 = 'b000100001;
    x_31 = 'b000100010;
    x_32 = 'b000101001;
    x_33 = 'b000100110;
    x_34 = 'b000100011;
    x_35 = 'b000011111;
    x_36 = 'b000011001;
    x_37 = 'b000010111;
    x_38 = 'b000010000;
    x_39 = 'b000001110;
    x_40 = 'b000010111;
    x_41 = 'b000001101;
    x_42 = 'b000001110;
    x_43 = 'b000100101;
    x_44 = 'b000000011;
    x_45 = 'b000010000;
    x_46 = 'b000010010;
    x_47 = 'b000010110;
    x_48 = 'b000001100;
    x_49 = 'b000010101;
    x_50 = 'b000011110;
    x_51 = 'b000100110;
    x_52 = 'b000100010;
    x_53 = 'b000100011;
    x_54 = 'b000011111;
    x_55 = 'b000010101;
    x_56 = 'b000011101;
    x_57 = 'b000011110;
    x_58 = 'b000100011;
    x_59 = 'b000010010;
    x_60 = 'b000001101;
    x_61 = 'b000001110;
    x_62 = 'b000000001;
    x_63 = 'b000001011;
    x_64 = 'b000010111;
    x_65 = 'b000011110;
    x_66 = 'b000100110;
    x_67 = 'b000101111;
    x_68 = 'b000101011;
    x_69 = 'b000100100;
    x_70 = 'b000100110;
    x_71 = 'b000000110;
    x_72 = 'b000010101;
    x_73 = 'b000011101;
    x_74 = 'b000100101;
    x_75 = 'b000110100;
    x_76 = 'b000101100;
    x_77 = 'b000101001;
    x_78 = 'b000001110;
    x_79 = 'b000011000;
    x_80 = 'b000011011;
    x_81 = 'b000100001;
    x_82 = 'b000100111;
    x_83 = 'b000101100;
    x_84 = 'b000101000;
    x_85 = 'b000011011;
    x_86 = 'b000010011;
    x_87 = 'b000010110;
    x_88 = 'b000011001;
    x_89 = 'b000011011;
    x_90 = 'b000100001;
    x_91 = 'b000011010;
    x_92 = 'b000010010;
    x_93 = 'b000010011;
    x_94 = 'b000100001;
    x_95 = 'b000100010;
    x_96 = 'b000101001;
    x_97 = 'b000100110;
    x_98 = 'b000100011;
    x_99 = 'b000011111;
    x_100 = 'b000011001;
    x_101 = 'b000010111;
    x_102 = 'b000010000;
    x_103 = 'b000001110;
    x_104 = 'b000010111;
    x_105 = 'b000001101;
    x_106 = 'b000001110;
    x_107 = 'b000100101;
    x_108 = 'b000000011;
    x_109 = 'b000010000;
    x_110 = 'b000010010;
    x_111 = 'b000010110;
    x_112 = 'b000001100;
    x_113 = 'b000010101;
    x_114 = 'b000011110;
    x_115 = 'b000100110;
    x_116 = 'b000100010;
    x_117 = 'b000100011;
    x_118 = 'b000011111;
    x_119 = 'b000010101;
    x_120 = 'b000011101;
    x_121 = 'b000011110;
    x_122 = 'b000100011;
    x_123 = 'b000010010;
    x_124 = 'b000001101;
    x_125 = 'b000001110;
    x_126 = 'b000000001;
    x_127 = 'b000001011;
    x_128 = 'b000010111;
    x_129 = 'b000011110;
    x_130 = 'b000100110;
    x_131 = 'b000101111;
    x_132 = 'b000101011;
    x_133 = 'b000100100;
    x_134 = 'b000100110;
    x_135 = 'b000000110;
    x_136 = 'b000010101;
    x_137 = 'b000011101;
    x_138 = 'b000100101;
    x_139 = 'b000110100;
    x_140 = 'b000101100;
    x_141 = 'b000101001;
    x_142 = 'b000001110;
    x_143 = 'b000011000;
    x_144 = 'b000011011;
    x_145 = 'b000100001;
    x_146 = 'b000100111;
    x_147 = 'b000101100;
    x_148 = 'b000101000;
    x_149 = 'b000011011;
    x_150 = 'b000010011;
    x_151 = 'b000010110;
    x_152 = 'b000011001;
    x_153 = 'b000011011;
    x_154 = 'b000100001;
    x_155 = 'b000011010;
    x_156 = 'b000010010;
    x_157 = 'b000010011;
    x_158 = 'b000100001;
    x_159 = 'b000100010;
    x_160 = 'b000101001;
    x_161 = 'b000100110;
    x_162 = 'b000100011;
    x_163 = 'b000011111;
    x_164 = 'b000011001;
    x_165 = 'b000010111;
    x_166 = 'b000010000;
    x_167 = 'b000001110;
    x_168 = 'b000010111;
    x_169 = 'b000001101;
    x_170 = 'b000001110;
    x_171 = 'b000100101;
    x_172 = 'b000000011;
    x_173 = 'b000010000;
    x_174 = 'b000010010;
    x_175 = 'b000010110;
    x_176 = 'b000001100;
    x_177 = 'b000010101;
    x_178 = 'b000011110;
    x_179 = 'b000100110;
    x_180 = 'b000100010;
    x_181 = 'b000100011;
    x_182 = 'b000011111;
    x_183 = 'b000010101;
    x_184 = 'b000011101;
    x_185 = 'b000011110;
    x_186 = 'b000100011;
    x_187 = 'b000010010;
    x_188 = 'b000001101;
    x_189 = 'b000001110;
    x_190 = 'b000000001;
    x_191 = 'b000001011;
    x_192 = 'b000010111;
    x_193 = 'b000011110;
    x_194 = 'b000100110;
    x_195 = 'b000101111;
    x_196 = 'b000101011;
    x_197 = 'b000100100;
    x_198 = 'b000100110;
    x_199 = 'b000000110;
    x_200 = 'b000010101;
    x_201 = 'b000011101;
    x_202 = 'b000100101;
    x_203 = 'b000110100;
    x_204 = 'b000101100;
    x_205 = 'b000101001;
    x_206 = 'b000001110;
    x_207 = 'b000011000;
    x_208 = 'b000011011;
    x_209 = 'b000100001;
    x_210 = 'b000100111;
    x_211 = 'b000101100;
    x_212 = 'b000101000;
    x_213 = 'b000011011;
    x_214 = 'b000010011;
    x_215 = 'b000010110;
    x_216 = 'b000011001;
    x_217 = 'b000011011;
    x_218 = 'b000100001;
    x_219 = 'b000011010;
    x_220 = 'b000010010;
    x_221 = 'b000010011;
    x_222 = 'b000100001;
    x_223 = 'b000100010;
    x_224 = 'b000101001;
    x_225 = 'b000100110;
    x_226 = 'b000100011;
    x_227 = 'b000011111;
    x_228 = 'b000011001;
    x_229 = 'b000010111;
    x_230 = 'b000010000;
    x_231 = 'b000001110;
    x_232 = 'b000010111;
    x_233 = 'b000001101;
    x_234 = 'b000001110;
    x_235 = 'b000100101;
    x_236 = 'b000000011;
    x_237 = 'b000010000;
    x_238 = 'b000010010;
    x_239 = 'b000010110;
    x_240 = 'b000001100;
    x_241 = 'b000010101;
    x_242 = 'b000011110;
    x_243 = 'b000100110;
    x_244 = 'b000100010;
    x_245 = 'b000100011;
    x_246 = 'b000011111;
    x_247 = 'b000010101;
    x_248 = 'b000011101;
    x_249 = 'b000011110;
    x_250 = 'b000100011;
    x_251 = 'b000010010;
    x_252 = 'b000001101;
    x_253 = 'b000001110;
    x_254 = 'b000000001;
    x_255 = 'b000001011;

    h_0 = 'b000010111;
    h_1 = 'b000011110;
    h_2 = 'b000100110;
    h_3 = 'b000101111;
    h_4 = 'b000101011;
    h_5 = 'b000100100;
    h_6 = 'b000100110;
    h_7 = 'b000000110;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000010001;
    x_1 = 'b000010011;
    x_2 = 'b000011010;
    x_3 = 'b000100010;
    x_4 = 'b000011111;
    x_5 = 'b000010011;
    x_6 = 'b000001110;
    x_7 = 'b000001000;
    x_8 = 'b000010000;
    x_9 = 'b000010100;
    x_10 = 'b000011010;
    x_11 = 'b000100101;
    x_12 = 'b000011010;
    x_13 = 'b000001001;
    x_14 = 'b000010011;
    x_15 = 'b000011010;
    x_16 = 'b000011001;
    x_17 = 'b000011010;
    x_18 = 'b000011011;
    x_19 = 'b000011100;
    x_20 = 'b000010011;
    x_21 = 'b000010100;
    x_22 = 'b000001100;
    x_23 = 'b000001111;
    x_24 = 'b000001101;
    x_25 = 'b000001111;
    x_26 = 'b000010011;
    x_27 = 'b000001101;
    x_28 = 'b000010001;
    x_29 = 'b000000111;
    x_30 = 'b000010011;
    x_31 = 'b000001111;
    x_32 = 'b000010110;
    x_33 = 'b000010011;
    x_34 = 'b000010000;
    x_35 = 'b000001001;
    x_36 = 'b000000010;
    x_37 = 'b000001001;
    x_38 = 'b000000111;
    x_39 = 'b111111010;
    x_40 = 'b000001001;
    x_41 = 'b111111101;
    x_42 = 'b000001100;
    x_43 = 'b000100011;
    x_44 = 'b000011000;
    x_45 = 'b000010011;
    x_46 = 'b000101010;
    x_47 = 'b000100010;
    x_48 = 'b000010011;
    x_49 = 'b000011011;
    x_50 = 'b000011101;
    x_51 = 'b000011111;
    x_52 = 'b000011001;
    x_53 = 'b000011100;
    x_54 = 'b000011100;
    x_55 = 'b000100011;
    x_56 = 'b000101010;
    x_57 = 'b000100010;
    x_58 = 'b000100001;
    x_59 = 'b000010101;
    x_60 = 'b000011000;
    x_61 = 'b000011001;
    x_62 = 'b000000110;
    x_63 = 'b000011001;
    x_64 = 'b000010001;
    x_65 = 'b000010011;
    x_66 = 'b000011010;
    x_67 = 'b000100010;
    x_68 = 'b000011111;
    x_69 = 'b000010011;
    x_70 = 'b000001110;
    x_71 = 'b000001000;
    x_72 = 'b000010000;
    x_73 = 'b000010100;
    x_74 = 'b000011010;
    x_75 = 'b000100101;
    x_76 = 'b000011010;
    x_77 = 'b000001001;
    x_78 = 'b000010011;
    x_79 = 'b000011010;
    x_80 = 'b000011001;
    x_81 = 'b000011010;
    x_82 = 'b000011011;
    x_83 = 'b000011100;
    x_84 = 'b000010011;
    x_85 = 'b000010100;
    x_86 = 'b000001100;
    x_87 = 'b000001111;
    x_88 = 'b000001101;
    x_89 = 'b000001111;
    x_90 = 'b000010011;
    x_91 = 'b000001101;
    x_92 = 'b000010001;
    x_93 = 'b000000111;
    x_94 = 'b000010011;
    x_95 = 'b000001111;
    x_96 = 'b000010110;
    x_97 = 'b000010011;
    x_98 = 'b000010000;
    x_99 = 'b000001001;
    x_100 = 'b000000010;
    x_101 = 'b000001001;
    x_102 = 'b000000111;
    x_103 = 'b111111010;
    x_104 = 'b000001001;
    x_105 = 'b111111101;
    x_106 = 'b000001100;
    x_107 = 'b000100011;
    x_108 = 'b000011000;
    x_109 = 'b000010011;
    x_110 = 'b000101010;
    x_111 = 'b000100010;
    x_112 = 'b000010011;
    x_113 = 'b000011011;
    x_114 = 'b000011101;
    x_115 = 'b000011111;
    x_116 = 'b000011001;
    x_117 = 'b000011100;
    x_118 = 'b000011100;
    x_119 = 'b000100011;
    x_120 = 'b000101010;
    x_121 = 'b000100010;
    x_122 = 'b000100001;
    x_123 = 'b000010101;
    x_124 = 'b000011000;
    x_125 = 'b000011001;
    x_126 = 'b000000110;
    x_127 = 'b000011001;
    x_128 = 'b000010001;
    x_129 = 'b000010011;
    x_130 = 'b000011010;
    x_131 = 'b000100010;
    x_132 = 'b000011111;
    x_133 = 'b000010011;
    x_134 = 'b000001110;
    x_135 = 'b000001000;
    x_136 = 'b000010000;
    x_137 = 'b000010100;
    x_138 = 'b000011010;
    x_139 = 'b000100101;
    x_140 = 'b000011010;
    x_141 = 'b000001001;
    x_142 = 'b000010011;
    x_143 = 'b000011010;
    x_144 = 'b000011001;
    x_145 = 'b000011010;
    x_146 = 'b000011011;
    x_147 = 'b000011100;
    x_148 = 'b000010011;
    x_149 = 'b000010100;
    x_150 = 'b000001100;
    x_151 = 'b000001111;
    x_152 = 'b000001101;
    x_153 = 'b000001111;
    x_154 = 'b000010011;
    x_155 = 'b000001101;
    x_156 = 'b000010001;
    x_157 = 'b000000111;
    x_158 = 'b000010011;
    x_159 = 'b000001111;
    x_160 = 'b000010110;
    x_161 = 'b000010011;
    x_162 = 'b000010000;
    x_163 = 'b000001001;
    x_164 = 'b000000010;
    x_165 = 'b000001001;
    x_166 = 'b000000111;
    x_167 = 'b111111010;
    x_168 = 'b000001001;
    x_169 = 'b111111101;
    x_170 = 'b000001100;
    x_171 = 'b000100011;
    x_172 = 'b000011000;
    x_173 = 'b000010011;
    x_174 = 'b000101010;
    x_175 = 'b000100010;
    x_176 = 'b000010011;
    x_177 = 'b000011011;
    x_178 = 'b000011101;
    x_179 = 'b000011111;
    x_180 = 'b000011001;
    x_181 = 'b000011100;
    x_182 = 'b000011100;
    x_183 = 'b000100011;
    x_184 = 'b000101010;
    x_185 = 'b000100010;
    x_186 = 'b000100001;
    x_187 = 'b000010101;
    x_188 = 'b000011000;
    x_189 = 'b000011001;
    x_190 = 'b000000110;
    x_191 = 'b000011001;
    x_192 = 'b000010001;
    x_193 = 'b000010011;
    x_194 = 'b000011010;
    x_195 = 'b000100010;
    x_196 = 'b000011111;
    x_197 = 'b000010011;
    x_198 = 'b000001110;
    x_199 = 'b000001000;
    x_200 = 'b000010000;
    x_201 = 'b000010100;
    x_202 = 'b000011010;
    x_203 = 'b000100101;
    x_204 = 'b000011010;
    x_205 = 'b000001001;
    x_206 = 'b000010011;
    x_207 = 'b000011010;
    x_208 = 'b000011001;
    x_209 = 'b000011010;
    x_210 = 'b000011011;
    x_211 = 'b000011100;
    x_212 = 'b000010011;
    x_213 = 'b000010100;
    x_214 = 'b000001100;
    x_215 = 'b000001111;
    x_216 = 'b000001101;
    x_217 = 'b000001111;
    x_218 = 'b000010011;
    x_219 = 'b000001101;
    x_220 = 'b000010001;
    x_221 = 'b000000111;
    x_222 = 'b000010011;
    x_223 = 'b000001111;
    x_224 = 'b000010110;
    x_225 = 'b000010011;
    x_226 = 'b000010000;
    x_227 = 'b000001001;
    x_228 = 'b000000010;
    x_229 = 'b000001001;
    x_230 = 'b000000111;
    x_231 = 'b111111010;
    x_232 = 'b000001001;
    x_233 = 'b111111101;
    x_234 = 'b000001100;
    x_235 = 'b000100011;
    x_236 = 'b000011000;
    x_237 = 'b000010011;
    x_238 = 'b000101010;
    x_239 = 'b000100010;
    x_240 = 'b000010011;
    x_241 = 'b000011011;
    x_242 = 'b000011101;
    x_243 = 'b000011111;
    x_244 = 'b000011001;
    x_245 = 'b000011100;
    x_246 = 'b000011100;
    x_247 = 'b000100011;
    x_248 = 'b000101010;
    x_249 = 'b000100010;
    x_250 = 'b000100001;
    x_251 = 'b000010101;
    x_252 = 'b000011000;
    x_253 = 'b000011001;
    x_254 = 'b000000110;
    x_255 = 'b000011001;

    h_0 = 'b000010001;
    h_1 = 'b000010011;
    h_2 = 'b000011010;
    h_3 = 'b000100010;
    h_4 = 'b000011111;
    h_5 = 'b000010011;
    h_6 = 'b000001110;
    h_7 = 'b000001000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000000110;
    x_1 = 'b000000111;
    x_2 = 'b000001011;
    x_3 = 'b000010001;
    x_4 = 'b000001101;
    x_5 = 'b000000000;
    x_6 = 'b111111100;
    x_7 = 'b111111111;
    x_8 = 'b000001100;
    x_9 = 'b000001111;
    x_10 = 'b000010001;
    x_11 = 'b000010010;
    x_12 = 'b000001011;
    x_13 = 'b111111100;
    x_14 = 'b000011000;
    x_15 = 'b000011100;
    x_16 = 'b000011000;
    x_17 = 'b000010111;
    x_18 = 'b000010001;
    x_19 = 'b000010001;
    x_20 = 'b000001011;
    x_21 = 'b000000111;
    x_22 = 'b000000010;
    x_23 = 'b000000110;
    x_24 = 'b000000111;
    x_25 = 'b000001000;
    x_26 = 'b000000100;
    x_27 = 'b111111110;
    x_28 = 'b000000111;
    x_29 = 'b000000011;
    x_30 = 'b000001111;
    x_31 = 'b000000110;
    x_32 = 'b000001101;
    x_33 = 'b000001000;
    x_34 = 'b000000011;
    x_35 = 'b111111110;
    x_36 = 'b111110110;
    x_37 = 'b000000000;
    x_38 = 'b000001110;
    x_39 = 'b111110011;
    x_40 = 'b000011110;
    x_41 = 'b000010010;
    x_42 = 'b000100001;
    x_43 = 'b000000110;
    x_44 = 'b000100111;
    x_45 = 'b000001111;
    x_46 = 'b000101101;
    x_47 = 'b000101001;
    x_48 = 'b000010111;
    x_49 = 'b000011111;
    x_50 = 'b000011100;
    x_51 = 'b000011011;
    x_52 = 'b000010100;
    x_53 = 'b000011000;
    x_54 = 'b000011010;
    x_55 = 'b000101011;
    x_56 = 'b000110000;
    x_57 = 'b000100110;
    x_58 = 'b000011110;
    x_59 = 'b000010110;
    x_60 = 'b000100110;
    x_61 = 'b000100101;
    x_62 = 'b000001100;
    x_63 = 'b000101010;
    x_64 = 'b000000110;
    x_65 = 'b000000111;
    x_66 = 'b000001011;
    x_67 = 'b000010001;
    x_68 = 'b000001101;
    x_69 = 'b000000000;
    x_70 = 'b111111100;
    x_71 = 'b111111111;
    x_72 = 'b000001100;
    x_73 = 'b000001111;
    x_74 = 'b000010001;
    x_75 = 'b000010010;
    x_76 = 'b000001011;
    x_77 = 'b111111100;
    x_78 = 'b000011000;
    x_79 = 'b000011100;
    x_80 = 'b000011000;
    x_81 = 'b000010111;
    x_82 = 'b000010001;
    x_83 = 'b000010001;
    x_84 = 'b000001011;
    x_85 = 'b000000111;
    x_86 = 'b000000010;
    x_87 = 'b000000110;
    x_88 = 'b000000111;
    x_89 = 'b000001000;
    x_90 = 'b000000100;
    x_91 = 'b111111110;
    x_92 = 'b000000111;
    x_93 = 'b000000011;
    x_94 = 'b000001111;
    x_95 = 'b000000110;
    x_96 = 'b000001101;
    x_97 = 'b000001000;
    x_98 = 'b000000011;
    x_99 = 'b111111110;
    x_100 = 'b111110110;
    x_101 = 'b000000000;
    x_102 = 'b000001110;
    x_103 = 'b111110011;
    x_104 = 'b000011110;
    x_105 = 'b000010010;
    x_106 = 'b000100001;
    x_107 = 'b000000110;
    x_108 = 'b000100111;
    x_109 = 'b000001111;
    x_110 = 'b000101101;
    x_111 = 'b000101001;
    x_112 = 'b000010111;
    x_113 = 'b000011111;
    x_114 = 'b000011100;
    x_115 = 'b000011011;
    x_116 = 'b000010100;
    x_117 = 'b000011000;
    x_118 = 'b000011010;
    x_119 = 'b000101011;
    x_120 = 'b000110000;
    x_121 = 'b000100110;
    x_122 = 'b000011110;
    x_123 = 'b000010110;
    x_124 = 'b000100110;
    x_125 = 'b000100101;
    x_126 = 'b000001100;
    x_127 = 'b000101010;
    x_128 = 'b000000110;
    x_129 = 'b000000111;
    x_130 = 'b000001011;
    x_131 = 'b000010001;
    x_132 = 'b000001101;
    x_133 = 'b000000000;
    x_134 = 'b111111100;
    x_135 = 'b111111111;
    x_136 = 'b000001100;
    x_137 = 'b000001111;
    x_138 = 'b000010001;
    x_139 = 'b000010010;
    x_140 = 'b000001011;
    x_141 = 'b111111100;
    x_142 = 'b000011000;
    x_143 = 'b000011100;
    x_144 = 'b000011000;
    x_145 = 'b000010111;
    x_146 = 'b000010001;
    x_147 = 'b000010001;
    x_148 = 'b000001011;
    x_149 = 'b000000111;
    x_150 = 'b000000010;
    x_151 = 'b000000110;
    x_152 = 'b000000111;
    x_153 = 'b000001000;
    x_154 = 'b000000100;
    x_155 = 'b111111110;
    x_156 = 'b000000111;
    x_157 = 'b000000011;
    x_158 = 'b000001111;
    x_159 = 'b000000110;
    x_160 = 'b000001101;
    x_161 = 'b000001000;
    x_162 = 'b000000011;
    x_163 = 'b111111110;
    x_164 = 'b111110110;
    x_165 = 'b000000000;
    x_166 = 'b000001110;
    x_167 = 'b111110011;
    x_168 = 'b000011110;
    x_169 = 'b000010010;
    x_170 = 'b000100001;
    x_171 = 'b000000110;
    x_172 = 'b000100111;
    x_173 = 'b000001111;
    x_174 = 'b000101101;
    x_175 = 'b000101001;
    x_176 = 'b000010111;
    x_177 = 'b000011111;
    x_178 = 'b000011100;
    x_179 = 'b000011011;
    x_180 = 'b000010100;
    x_181 = 'b000011000;
    x_182 = 'b000011010;
    x_183 = 'b000101011;
    x_184 = 'b000110000;
    x_185 = 'b000100110;
    x_186 = 'b000011110;
    x_187 = 'b000010110;
    x_188 = 'b000100110;
    x_189 = 'b000100101;
    x_190 = 'b000001100;
    x_191 = 'b000101010;
    x_192 = 'b000000110;
    x_193 = 'b000000111;
    x_194 = 'b000001011;
    x_195 = 'b000010001;
    x_196 = 'b000001101;
    x_197 = 'b000000000;
    x_198 = 'b111111100;
    x_199 = 'b111111111;
    x_200 = 'b000001100;
    x_201 = 'b000001111;
    x_202 = 'b000010001;
    x_203 = 'b000010010;
    x_204 = 'b000001011;
    x_205 = 'b111111100;
    x_206 = 'b000011000;
    x_207 = 'b000011100;
    x_208 = 'b000011000;
    x_209 = 'b000010111;
    x_210 = 'b000010001;
    x_211 = 'b000010001;
    x_212 = 'b000001011;
    x_213 = 'b000000111;
    x_214 = 'b000000010;
    x_215 = 'b000000110;
    x_216 = 'b000000111;
    x_217 = 'b000001000;
    x_218 = 'b000000100;
    x_219 = 'b111111110;
    x_220 = 'b000000111;
    x_221 = 'b000000011;
    x_222 = 'b000001111;
    x_223 = 'b000000110;
    x_224 = 'b000001101;
    x_225 = 'b000001000;
    x_226 = 'b000000011;
    x_227 = 'b111111110;
    x_228 = 'b111110110;
    x_229 = 'b000000000;
    x_230 = 'b000001110;
    x_231 = 'b111110011;
    x_232 = 'b000011110;
    x_233 = 'b000010010;
    x_234 = 'b000100001;
    x_235 = 'b000000110;
    x_236 = 'b000100111;
    x_237 = 'b000001111;
    x_238 = 'b000101101;
    x_239 = 'b000101001;
    x_240 = 'b000010111;
    x_241 = 'b000011111;
    x_242 = 'b000011100;
    x_243 = 'b000011011;
    x_244 = 'b000010100;
    x_245 = 'b000011000;
    x_246 = 'b000011010;
    x_247 = 'b000101011;
    x_248 = 'b000110000;
    x_249 = 'b000100110;
    x_250 = 'b000011110;
    x_251 = 'b000010110;
    x_252 = 'b000100110;
    x_253 = 'b000100101;
    x_254 = 'b000001100;
    x_255 = 'b000101010;

    h_0 = 'b000000110;
    h_1 = 'b000000111;
    h_2 = 'b000001011;
    h_3 = 'b000010001;
    h_4 = 'b000001101;
    h_5 = 'b000000000;
    h_6 = 'b111111100;
    h_7 = 'b111111111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000010101;
    x_1 = 'b000010000;
    x_2 = 'b000010000;
    x_3 = 'b000010001;
    x_4 = 'b000001101;
    x_5 = 'b111111101;
    x_6 = 'b111111011;
    x_7 = 'b000001101;
    x_8 = 'b000010100;
    x_9 = 'b000010001;
    x_10 = 'b000001110;
    x_11 = 'b000001111;
    x_12 = 'b000000110;
    x_13 = 'b111111011;
    x_14 = 'b000100000;
    x_15 = 'b000011111;
    x_16 = 'b000011000;
    x_17 = 'b000010001;
    x_18 = 'b000001011;
    x_19 = 'b000001100;
    x_20 = 'b000000110;
    x_21 = 'b000001011;
    x_22 = 'b000000100;
    x_23 = 'b000000100;
    x_24 = 'b000001100;
    x_25 = 'b000001101;
    x_26 = 'b000000110;
    x_27 = 'b111111111;
    x_28 = 'b000000100;
    x_29 = 'b000010000;
    x_30 = 'b000010001;
    x_31 = 'b000000111;
    x_32 = 'b000010010;
    x_33 = 'b000001110;
    x_34 = 'b000001000;
    x_35 = 'b000000011;
    x_36 = 'b111111000;
    x_37 = 'b000000010;
    x_38 = 'b000010011;
    x_39 = 'b111101110;
    x_40 = 'b000100110;
    x_41 = 'b111111000;
    x_42 = 'b000101101;
    x_43 = 'b111101010;
    x_44 = 'b000101000;
    x_45 = 'b000000000;
    x_46 = 'b000101010;
    x_47 = 'b000101001;
    x_48 = 'b000010111;
    x_49 = 'b000011011;
    x_50 = 'b000010110;
    x_51 = 'b000010100;
    x_52 = 'b000001011;
    x_53 = 'b000001110;
    x_54 = 'b000001100;
    x_55 = 'b000101010;
    x_56 = 'b000101110;
    x_57 = 'b000100011;
    x_58 = 'b000010110;
    x_59 = 'b000001010;
    x_60 = 'b000101011;
    x_61 = 'b000101000;
    x_62 = 'b000001100;
    x_63 = 'b000101111;
    x_64 = 'b000010101;
    x_65 = 'b000010000;
    x_66 = 'b000010000;
    x_67 = 'b000010001;
    x_68 = 'b000001101;
    x_69 = 'b111111101;
    x_70 = 'b111111011;
    x_71 = 'b000001101;
    x_72 = 'b000010100;
    x_73 = 'b000010001;
    x_74 = 'b000001110;
    x_75 = 'b000001111;
    x_76 = 'b000000110;
    x_77 = 'b111111011;
    x_78 = 'b000100000;
    x_79 = 'b000011111;
    x_80 = 'b000011000;
    x_81 = 'b000010001;
    x_82 = 'b000001011;
    x_83 = 'b000001100;
    x_84 = 'b000000110;
    x_85 = 'b000001011;
    x_86 = 'b000000100;
    x_87 = 'b000000100;
    x_88 = 'b000001100;
    x_89 = 'b000001101;
    x_90 = 'b000000110;
    x_91 = 'b111111111;
    x_92 = 'b000000100;
    x_93 = 'b000010000;
    x_94 = 'b000010001;
    x_95 = 'b000000111;
    x_96 = 'b000010010;
    x_97 = 'b000001110;
    x_98 = 'b000001000;
    x_99 = 'b000000011;
    x_100 = 'b111111000;
    x_101 = 'b000000010;
    x_102 = 'b000010011;
    x_103 = 'b111101110;
    x_104 = 'b000100110;
    x_105 = 'b111111000;
    x_106 = 'b000101101;
    x_107 = 'b111101010;
    x_108 = 'b000101000;
    x_109 = 'b000000000;
    x_110 = 'b000101010;
    x_111 = 'b000101001;
    x_112 = 'b000010111;
    x_113 = 'b000011011;
    x_114 = 'b000010110;
    x_115 = 'b000010100;
    x_116 = 'b000001011;
    x_117 = 'b000001110;
    x_118 = 'b000001100;
    x_119 = 'b000101010;
    x_120 = 'b000101110;
    x_121 = 'b000100011;
    x_122 = 'b000010110;
    x_123 = 'b000001010;
    x_124 = 'b000101011;
    x_125 = 'b000101000;
    x_126 = 'b000001100;
    x_127 = 'b000101111;
    x_128 = 'b000010101;
    x_129 = 'b000010000;
    x_130 = 'b000010000;
    x_131 = 'b000010001;
    x_132 = 'b000001101;
    x_133 = 'b111111101;
    x_134 = 'b111111011;
    x_135 = 'b000001101;
    x_136 = 'b000010100;
    x_137 = 'b000010001;
    x_138 = 'b000001110;
    x_139 = 'b000001111;
    x_140 = 'b000000110;
    x_141 = 'b111111011;
    x_142 = 'b000100000;
    x_143 = 'b000011111;
    x_144 = 'b000011000;
    x_145 = 'b000010001;
    x_146 = 'b000001011;
    x_147 = 'b000001100;
    x_148 = 'b000000110;
    x_149 = 'b000001011;
    x_150 = 'b000000100;
    x_151 = 'b000000100;
    x_152 = 'b000001100;
    x_153 = 'b000001101;
    x_154 = 'b000000110;
    x_155 = 'b111111111;
    x_156 = 'b000000100;
    x_157 = 'b000010000;
    x_158 = 'b000010001;
    x_159 = 'b000000111;
    x_160 = 'b000010010;
    x_161 = 'b000001110;
    x_162 = 'b000001000;
    x_163 = 'b000000011;
    x_164 = 'b111111000;
    x_165 = 'b000000010;
    x_166 = 'b000010011;
    x_167 = 'b111101110;
    x_168 = 'b000100110;
    x_169 = 'b111111000;
    x_170 = 'b000101101;
    x_171 = 'b111101010;
    x_172 = 'b000101000;
    x_173 = 'b000000000;
    x_174 = 'b000101010;
    x_175 = 'b000101001;
    x_176 = 'b000010111;
    x_177 = 'b000011011;
    x_178 = 'b000010110;
    x_179 = 'b000010100;
    x_180 = 'b000001011;
    x_181 = 'b000001110;
    x_182 = 'b000001100;
    x_183 = 'b000101010;
    x_184 = 'b000101110;
    x_185 = 'b000100011;
    x_186 = 'b000010110;
    x_187 = 'b000001010;
    x_188 = 'b000101011;
    x_189 = 'b000101000;
    x_190 = 'b000001100;
    x_191 = 'b000101111;
    x_192 = 'b000010101;
    x_193 = 'b000010000;
    x_194 = 'b000010000;
    x_195 = 'b000010001;
    x_196 = 'b000001101;
    x_197 = 'b111111101;
    x_198 = 'b111111011;
    x_199 = 'b000001101;
    x_200 = 'b000010100;
    x_201 = 'b000010001;
    x_202 = 'b000001110;
    x_203 = 'b000001111;
    x_204 = 'b000000110;
    x_205 = 'b111111011;
    x_206 = 'b000100000;
    x_207 = 'b000011111;
    x_208 = 'b000011000;
    x_209 = 'b000010001;
    x_210 = 'b000001011;
    x_211 = 'b000001100;
    x_212 = 'b000000110;
    x_213 = 'b000001011;
    x_214 = 'b000000100;
    x_215 = 'b000000100;
    x_216 = 'b000001100;
    x_217 = 'b000001101;
    x_218 = 'b000000110;
    x_219 = 'b111111111;
    x_220 = 'b000000100;
    x_221 = 'b000010000;
    x_222 = 'b000010001;
    x_223 = 'b000000111;
    x_224 = 'b000010010;
    x_225 = 'b000001110;
    x_226 = 'b000001000;
    x_227 = 'b000000011;
    x_228 = 'b111111000;
    x_229 = 'b000000010;
    x_230 = 'b000010011;
    x_231 = 'b111101110;
    x_232 = 'b000100110;
    x_233 = 'b111111000;
    x_234 = 'b000101101;
    x_235 = 'b111101010;
    x_236 = 'b000101000;
    x_237 = 'b000000000;
    x_238 = 'b000101010;
    x_239 = 'b000101001;
    x_240 = 'b000010111;
    x_241 = 'b000011011;
    x_242 = 'b000010110;
    x_243 = 'b000010100;
    x_244 = 'b000001011;
    x_245 = 'b000001110;
    x_246 = 'b000001100;
    x_247 = 'b000101010;
    x_248 = 'b000101110;
    x_249 = 'b000100011;
    x_250 = 'b000010110;
    x_251 = 'b000001010;
    x_252 = 'b000101011;
    x_253 = 'b000101000;
    x_254 = 'b000001100;
    x_255 = 'b000101111;

    h_0 = 'b000010101;
    h_1 = 'b000010000;
    h_2 = 'b000010000;
    h_3 = 'b000010001;
    h_4 = 'b000001101;
    h_5 = 'b111111101;
    h_6 = 'b111111011;
    h_7 = 'b000001101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000010101;
    x_1 = 'b000010010;
    x_2 = 'b000010001;
    x_3 = 'b000010010;
    x_4 = 'b000001010;
    x_5 = 'b111111001;
    x_6 = 'b111111000;
    x_7 = 'b000010000;
    x_8 = 'b000010010;
    x_9 = 'b000001110;
    x_10 = 'b000001101;
    x_11 = 'b000001101;
    x_12 = 'b000000000;
    x_13 = 'b111110010;
    x_14 = 'b000100000;
    x_15 = 'b000011100;
    x_16 = 'b000010100;
    x_17 = 'b000001100;
    x_18 = 'b000001001;
    x_19 = 'b000001001;
    x_20 = 'b000000000;
    x_21 = 'b000001100;
    x_22 = 'b000000001;
    x_23 = 'b000000010;
    x_24 = 'b000001111;
    x_25 = 'b000010000;
    x_26 = 'b000000100;
    x_27 = 'b111111110;
    x_28 = 'b000000100;
    x_29 = 'b000010110;
    x_30 = 'b000001011;
    x_31 = 'b000000110;
    x_32 = 'b000001111;
    x_33 = 'b000001001;
    x_34 = 'b000000011;
    x_35 = 'b111111100;
    x_36 = 'b111110111;
    x_37 = 'b000000010;
    x_38 = 'b000011000;
    x_39 = 'b111100111;
    x_40 = 'b000101011;
    x_41 = 'b111100010;
    x_42 = 'b000100110;
    x_43 = 'b000110000;
    x_44 = 'b000100111;
    x_45 = 'b111111101;
    x_46 = 'b000100101;
    x_47 = 'b000100010;
    x_48 = 'b000010010;
    x_49 = 'b000011000;
    x_50 = 'b000010101;
    x_51 = 'b000010011;
    x_52 = 'b000001010;
    x_53 = 'b000001011;
    x_54 = 'b000000100;
    x_55 = 'b000011101;
    x_56 = 'b000100100;
    x_57 = 'b000011100;
    x_58 = 'b000010000;
    x_59 = 'b000000010;
    x_60 = 'b000100100;
    x_61 = 'b000100001;
    x_62 = 'b000000100;
    x_63 = 'b000100000;
    x_64 = 'b000010101;
    x_65 = 'b000010010;
    x_66 = 'b000010001;
    x_67 = 'b000010010;
    x_68 = 'b000001010;
    x_69 = 'b111111001;
    x_70 = 'b111111000;
    x_71 = 'b000010000;
    x_72 = 'b000010010;
    x_73 = 'b000001110;
    x_74 = 'b000001101;
    x_75 = 'b000001101;
    x_76 = 'b000000000;
    x_77 = 'b111110010;
    x_78 = 'b000100000;
    x_79 = 'b000011100;
    x_80 = 'b000010100;
    x_81 = 'b000001100;
    x_82 = 'b000001001;
    x_83 = 'b000001001;
    x_84 = 'b000000000;
    x_85 = 'b000001100;
    x_86 = 'b000000001;
    x_87 = 'b000000010;
    x_88 = 'b000001111;
    x_89 = 'b000010000;
    x_90 = 'b000000100;
    x_91 = 'b111111110;
    x_92 = 'b000000100;
    x_93 = 'b000010110;
    x_94 = 'b000001011;
    x_95 = 'b000000110;
    x_96 = 'b000001111;
    x_97 = 'b000001001;
    x_98 = 'b000000011;
    x_99 = 'b111111100;
    x_100 = 'b111110111;
    x_101 = 'b000000010;
    x_102 = 'b000011000;
    x_103 = 'b111100111;
    x_104 = 'b000101011;
    x_105 = 'b111100010;
    x_106 = 'b000100110;
    x_107 = 'b000110000;
    x_108 = 'b000100111;
    x_109 = 'b111111101;
    x_110 = 'b000100101;
    x_111 = 'b000100010;
    x_112 = 'b000010010;
    x_113 = 'b000011000;
    x_114 = 'b000010101;
    x_115 = 'b000010011;
    x_116 = 'b000001010;
    x_117 = 'b000001011;
    x_118 = 'b000000100;
    x_119 = 'b000011101;
    x_120 = 'b000100100;
    x_121 = 'b000011100;
    x_122 = 'b000010000;
    x_123 = 'b000000010;
    x_124 = 'b000100100;
    x_125 = 'b000100001;
    x_126 = 'b000000100;
    x_127 = 'b000100000;
    x_128 = 'b000010101;
    x_129 = 'b000010010;
    x_130 = 'b000010001;
    x_131 = 'b000010010;
    x_132 = 'b000001010;
    x_133 = 'b111111001;
    x_134 = 'b111111000;
    x_135 = 'b000010000;
    x_136 = 'b000010010;
    x_137 = 'b000001110;
    x_138 = 'b000001101;
    x_139 = 'b000001101;
    x_140 = 'b000000000;
    x_141 = 'b111110010;
    x_142 = 'b000100000;
    x_143 = 'b000011100;
    x_144 = 'b000010100;
    x_145 = 'b000001100;
    x_146 = 'b000001001;
    x_147 = 'b000001001;
    x_148 = 'b000000000;
    x_149 = 'b000001100;
    x_150 = 'b000000001;
    x_151 = 'b000000010;
    x_152 = 'b000001111;
    x_153 = 'b000010000;
    x_154 = 'b000000100;
    x_155 = 'b111111110;
    x_156 = 'b000000100;
    x_157 = 'b000010110;
    x_158 = 'b000001011;
    x_159 = 'b000000110;
    x_160 = 'b000001111;
    x_161 = 'b000001001;
    x_162 = 'b000000011;
    x_163 = 'b111111100;
    x_164 = 'b111110111;
    x_165 = 'b000000010;
    x_166 = 'b000011000;
    x_167 = 'b111100111;
    x_168 = 'b000101011;
    x_169 = 'b111100010;
    x_170 = 'b000100110;
    x_171 = 'b000110000;
    x_172 = 'b000100111;
    x_173 = 'b111111101;
    x_174 = 'b000100101;
    x_175 = 'b000100010;
    x_176 = 'b000010010;
    x_177 = 'b000011000;
    x_178 = 'b000010101;
    x_179 = 'b000010011;
    x_180 = 'b000001010;
    x_181 = 'b000001011;
    x_182 = 'b000000100;
    x_183 = 'b000011101;
    x_184 = 'b000100100;
    x_185 = 'b000011100;
    x_186 = 'b000010000;
    x_187 = 'b000000010;
    x_188 = 'b000100100;
    x_189 = 'b000100001;
    x_190 = 'b000000100;
    x_191 = 'b000100000;
    x_192 = 'b000010101;
    x_193 = 'b000010010;
    x_194 = 'b000010001;
    x_195 = 'b000010010;
    x_196 = 'b000001010;
    x_197 = 'b111111001;
    x_198 = 'b111111000;
    x_199 = 'b000010000;
    x_200 = 'b000010010;
    x_201 = 'b000001110;
    x_202 = 'b000001101;
    x_203 = 'b000001101;
    x_204 = 'b000000000;
    x_205 = 'b111110010;
    x_206 = 'b000100000;
    x_207 = 'b000011100;
    x_208 = 'b000010100;
    x_209 = 'b000001100;
    x_210 = 'b000001001;
    x_211 = 'b000001001;
    x_212 = 'b000000000;
    x_213 = 'b000001100;
    x_214 = 'b000000001;
    x_215 = 'b000000010;
    x_216 = 'b000001111;
    x_217 = 'b000010000;
    x_218 = 'b000000100;
    x_219 = 'b111111110;
    x_220 = 'b000000100;
    x_221 = 'b000010110;
    x_222 = 'b000001011;
    x_223 = 'b000000110;
    x_224 = 'b000001111;
    x_225 = 'b000001001;
    x_226 = 'b000000011;
    x_227 = 'b111111100;
    x_228 = 'b111110111;
    x_229 = 'b000000010;
    x_230 = 'b000011000;
    x_231 = 'b111100111;
    x_232 = 'b000101011;
    x_233 = 'b111100010;
    x_234 = 'b000100110;
    x_235 = 'b000110000;
    x_236 = 'b000100111;
    x_237 = 'b111111101;
    x_238 = 'b000100101;
    x_239 = 'b000100010;
    x_240 = 'b000010010;
    x_241 = 'b000011000;
    x_242 = 'b000010101;
    x_243 = 'b000010011;
    x_244 = 'b000001010;
    x_245 = 'b000001011;
    x_246 = 'b000000100;
    x_247 = 'b000011101;
    x_248 = 'b000100100;
    x_249 = 'b000011100;
    x_250 = 'b000010000;
    x_251 = 'b000000010;
    x_252 = 'b000100100;
    x_253 = 'b000100001;
    x_254 = 'b000000100;
    x_255 = 'b000100000;

    h_0 = 'b000010101;
    h_1 = 'b000010010;
    h_2 = 'b000010001;
    h_3 = 'b000010010;
    h_4 = 'b000001010;
    h_5 = 'b111111001;
    h_6 = 'b111111000;
    h_7 = 'b000010000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000001111;
    x_1 = 'b000000110;
    x_2 = 'b000001000;
    x_3 = 'b000001101;
    x_4 = 'b111111110;
    x_5 = 'b111101101;
    x_6 = 'b111101110;
    x_7 = 'b000000001;
    x_8 = 'b000000111;
    x_9 = 'b000000110;
    x_10 = 'b000001000;
    x_11 = 'b000000100;
    x_12 = 'b111110101;
    x_13 = 'b111101100;
    x_14 = 'b000001111;
    x_15 = 'b000001111;
    x_16 = 'b000001001;
    x_17 = 'b000000101;
    x_18 = 'b000000010;
    x_19 = 'b000000001;
    x_20 = 'b111110111;
    x_21 = 'b000000111;
    x_22 = 'b111110101;
    x_23 = 'b111110111;
    x_24 = 'b000001011;
    x_25 = 'b000001100;
    x_26 = 'b111110100;
    x_27 = 'b111101110;
    x_28 = 'b111110111;
    x_29 = 'b000001110;
    x_30 = 'b000000101;
    x_31 = 'b111111001;
    x_32 = 'b000000100;
    x_33 = 'b111111001;
    x_34 = 'b111110010;
    x_35 = 'b111101111;
    x_36 = 'b111100101;
    x_37 = 'b111110101;
    x_38 = 'b000010110;
    x_39 = 'b111011010;
    x_40 = 'b000100100;
    x_41 = 'b111101001;
    x_42 = 'b000001100;
    x_43 = 'b000101011;
    x_44 = 'b000010000;
    x_45 = 'b111011001;
    x_46 = 'b000001110;
    x_47 = 'b000001111;
    x_48 = 'b000000010;
    x_49 = 'b000001001;
    x_50 = 'b000000111;
    x_51 = 'b000000101;
    x_52 = 'b111111011;
    x_53 = 'b111111000;
    x_54 = 'b111101011;
    x_55 = 'b000001100;
    x_56 = 'b000010011;
    x_57 = 'b000001111;
    x_58 = 'b000000010;
    x_59 = 'b111110110;
    x_60 = 'b000010101;
    x_61 = 'b000010000;
    x_62 = 'b111110100;
    x_63 = 'b000001000;
    x_64 = 'b000001111;
    x_65 = 'b000000110;
    x_66 = 'b000001000;
    x_67 = 'b000001101;
    x_68 = 'b111111110;
    x_69 = 'b111101101;
    x_70 = 'b111101110;
    x_71 = 'b000000001;
    x_72 = 'b000000111;
    x_73 = 'b000000110;
    x_74 = 'b000001000;
    x_75 = 'b000000100;
    x_76 = 'b111110101;
    x_77 = 'b111101100;
    x_78 = 'b000001111;
    x_79 = 'b000001111;
    x_80 = 'b000001001;
    x_81 = 'b000000101;
    x_82 = 'b000000010;
    x_83 = 'b000000001;
    x_84 = 'b111110111;
    x_85 = 'b000000111;
    x_86 = 'b111110101;
    x_87 = 'b111110111;
    x_88 = 'b000001011;
    x_89 = 'b000001100;
    x_90 = 'b111110100;
    x_91 = 'b111101110;
    x_92 = 'b111110111;
    x_93 = 'b000001110;
    x_94 = 'b000000101;
    x_95 = 'b111111001;
    x_96 = 'b000000100;
    x_97 = 'b111111001;
    x_98 = 'b111110010;
    x_99 = 'b111101111;
    x_100 = 'b111100101;
    x_101 = 'b111110101;
    x_102 = 'b000010110;
    x_103 = 'b111011010;
    x_104 = 'b000100100;
    x_105 = 'b111101001;
    x_106 = 'b000001100;
    x_107 = 'b000101011;
    x_108 = 'b000010000;
    x_109 = 'b111011001;
    x_110 = 'b000001110;
    x_111 = 'b000001111;
    x_112 = 'b000000010;
    x_113 = 'b000001001;
    x_114 = 'b000000111;
    x_115 = 'b000000101;
    x_116 = 'b111111011;
    x_117 = 'b111111000;
    x_118 = 'b111101011;
    x_119 = 'b000001100;
    x_120 = 'b000010011;
    x_121 = 'b000001111;
    x_122 = 'b000000010;
    x_123 = 'b111110110;
    x_124 = 'b000010101;
    x_125 = 'b000010000;
    x_126 = 'b111110100;
    x_127 = 'b000001000;
    x_128 = 'b000001111;
    x_129 = 'b000000110;
    x_130 = 'b000001000;
    x_131 = 'b000001101;
    x_132 = 'b111111110;
    x_133 = 'b111101101;
    x_134 = 'b111101110;
    x_135 = 'b000000001;
    x_136 = 'b000000111;
    x_137 = 'b000000110;
    x_138 = 'b000001000;
    x_139 = 'b000000100;
    x_140 = 'b111110101;
    x_141 = 'b111101100;
    x_142 = 'b000001111;
    x_143 = 'b000001111;
    x_144 = 'b000001001;
    x_145 = 'b000000101;
    x_146 = 'b000000010;
    x_147 = 'b000000001;
    x_148 = 'b111110111;
    x_149 = 'b000000111;
    x_150 = 'b111110101;
    x_151 = 'b111110111;
    x_152 = 'b000001011;
    x_153 = 'b000001100;
    x_154 = 'b111110100;
    x_155 = 'b111101110;
    x_156 = 'b111110111;
    x_157 = 'b000001110;
    x_158 = 'b000000101;
    x_159 = 'b111111001;
    x_160 = 'b000000100;
    x_161 = 'b111111001;
    x_162 = 'b111110010;
    x_163 = 'b111101111;
    x_164 = 'b111100101;
    x_165 = 'b111110101;
    x_166 = 'b000010110;
    x_167 = 'b111011010;
    x_168 = 'b000100100;
    x_169 = 'b111101001;
    x_170 = 'b000001100;
    x_171 = 'b000101011;
    x_172 = 'b000010000;
    x_173 = 'b111011001;
    x_174 = 'b000001110;
    x_175 = 'b000001111;
    x_176 = 'b000000010;
    x_177 = 'b000001001;
    x_178 = 'b000000111;
    x_179 = 'b000000101;
    x_180 = 'b111111011;
    x_181 = 'b111111000;
    x_182 = 'b111101011;
    x_183 = 'b000001100;
    x_184 = 'b000010011;
    x_185 = 'b000001111;
    x_186 = 'b000000010;
    x_187 = 'b111110110;
    x_188 = 'b000010101;
    x_189 = 'b000010000;
    x_190 = 'b111110100;
    x_191 = 'b000001000;
    x_192 = 'b000001111;
    x_193 = 'b000000110;
    x_194 = 'b000001000;
    x_195 = 'b000001101;
    x_196 = 'b111111110;
    x_197 = 'b111101101;
    x_198 = 'b111101110;
    x_199 = 'b000000001;
    x_200 = 'b000000111;
    x_201 = 'b000000110;
    x_202 = 'b000001000;
    x_203 = 'b000000100;
    x_204 = 'b111110101;
    x_205 = 'b111101100;
    x_206 = 'b000001111;
    x_207 = 'b000001111;
    x_208 = 'b000001001;
    x_209 = 'b000000101;
    x_210 = 'b000000010;
    x_211 = 'b000000001;
    x_212 = 'b111110111;
    x_213 = 'b000000111;
    x_214 = 'b111110101;
    x_215 = 'b111110111;
    x_216 = 'b000001011;
    x_217 = 'b000001100;
    x_218 = 'b111110100;
    x_219 = 'b111101110;
    x_220 = 'b111110111;
    x_221 = 'b000001110;
    x_222 = 'b000000101;
    x_223 = 'b111111001;
    x_224 = 'b000000100;
    x_225 = 'b111111001;
    x_226 = 'b111110010;
    x_227 = 'b111101111;
    x_228 = 'b111100101;
    x_229 = 'b111110101;
    x_230 = 'b000010110;
    x_231 = 'b111011010;
    x_232 = 'b000100100;
    x_233 = 'b111101001;
    x_234 = 'b000001100;
    x_235 = 'b000101011;
    x_236 = 'b000010000;
    x_237 = 'b111011001;
    x_238 = 'b000001110;
    x_239 = 'b000001111;
    x_240 = 'b000000010;
    x_241 = 'b000001001;
    x_242 = 'b000000111;
    x_243 = 'b000000101;
    x_244 = 'b111111011;
    x_245 = 'b111111000;
    x_246 = 'b111101011;
    x_247 = 'b000001100;
    x_248 = 'b000010011;
    x_249 = 'b000001111;
    x_250 = 'b000000010;
    x_251 = 'b111110110;
    x_252 = 'b000010101;
    x_253 = 'b000010000;
    x_254 = 'b111110100;
    x_255 = 'b000001000;

    h_0 = 'b000001111;
    h_1 = 'b000000110;
    h_2 = 'b000001000;
    h_3 = 'b000001101;
    h_4 = 'b111111110;
    h_5 = 'b111101101;
    h_6 = 'b111101110;
    h_7 = 'b000000001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000010100;
    x_1 = 'b000001011;
    x_2 = 'b000001011;
    x_3 = 'b000001110;
    x_4 = 'b000000001;
    x_5 = 'b111101110;
    x_6 = 'b111100111;
    x_7 = 'b000001101;
    x_8 = 'b000010000;
    x_9 = 'b000010001;
    x_10 = 'b000010011;
    x_11 = 'b000010001;
    x_12 = 'b111111101;
    x_13 = 'b111110000;
    x_14 = 'b000010101;
    x_15 = 'b000011001;
    x_16 = 'b000010011;
    x_17 = 'b000010001;
    x_18 = 'b000010000;
    x_19 = 'b000001110;
    x_20 = 'b111111111;
    x_21 = 'b000000011;
    x_22 = 'b111110111;
    x_23 = 'b111111011;
    x_24 = 'b000001001;
    x_25 = 'b000001011;
    x_26 = 'b111111101;
    x_27 = 'b111110011;
    x_28 = 'b111111011;
    x_29 = 'b000001111;
    x_30 = 'b000000111;
    x_31 = 'b000000100;
    x_32 = 'b000010010;
    x_33 = 'b000001011;
    x_34 = 'b000000010;
    x_35 = 'b111111110;
    x_36 = 'b111110010;
    x_37 = 'b000000110;
    x_38 = 'b000011100;
    x_39 = 'b111110000;
    x_40 = 'b000100000;
    x_41 = 'b000001100;
    x_42 = 'b000011001;
    x_43 = 'b000011011;
    x_44 = 'b000010111;
    x_45 = 'b000001100;
    x_46 = 'b000011001;
    x_47 = 'b000011101;
    x_48 = 'b000010001;
    x_49 = 'b000011010;
    x_50 = 'b000011011;
    x_51 = 'b000011001;
    x_52 = 'b000010001;
    x_53 = 'b000010000;
    x_54 = 'b000001101;
    x_55 = 'b000011000;
    x_56 = 'b000100001;
    x_57 = 'b000011101;
    x_58 = 'b000010010;
    x_59 = 'b000000101;
    x_60 = 'b000010001;
    x_61 = 'b000001111;
    x_62 = 'b111110011;
    x_63 = 'b000001000;
    x_64 = 'b000010100;
    x_65 = 'b000001011;
    x_66 = 'b000001011;
    x_67 = 'b000001110;
    x_68 = 'b000000001;
    x_69 = 'b111101110;
    x_70 = 'b111100111;
    x_71 = 'b000001101;
    x_72 = 'b000010000;
    x_73 = 'b000010001;
    x_74 = 'b000010011;
    x_75 = 'b000010001;
    x_76 = 'b111111101;
    x_77 = 'b111110000;
    x_78 = 'b000010101;
    x_79 = 'b000011001;
    x_80 = 'b000010011;
    x_81 = 'b000010001;
    x_82 = 'b000010000;
    x_83 = 'b000001110;
    x_84 = 'b111111111;
    x_85 = 'b000000011;
    x_86 = 'b111110111;
    x_87 = 'b111111011;
    x_88 = 'b000001001;
    x_89 = 'b000001011;
    x_90 = 'b111111101;
    x_91 = 'b111110011;
    x_92 = 'b111111011;
    x_93 = 'b000001111;
    x_94 = 'b000000111;
    x_95 = 'b000000100;
    x_96 = 'b000010010;
    x_97 = 'b000001011;
    x_98 = 'b000000010;
    x_99 = 'b111111110;
    x_100 = 'b111110010;
    x_101 = 'b000000110;
    x_102 = 'b000011100;
    x_103 = 'b111110000;
    x_104 = 'b000100000;
    x_105 = 'b000001100;
    x_106 = 'b000011001;
    x_107 = 'b000011011;
    x_108 = 'b000010111;
    x_109 = 'b000001100;
    x_110 = 'b000011001;
    x_111 = 'b000011101;
    x_112 = 'b000010001;
    x_113 = 'b000011010;
    x_114 = 'b000011011;
    x_115 = 'b000011001;
    x_116 = 'b000010001;
    x_117 = 'b000010000;
    x_118 = 'b000001101;
    x_119 = 'b000011000;
    x_120 = 'b000100001;
    x_121 = 'b000011101;
    x_122 = 'b000010010;
    x_123 = 'b000000101;
    x_124 = 'b000010001;
    x_125 = 'b000001111;
    x_126 = 'b111110011;
    x_127 = 'b000001000;
    x_128 = 'b000010100;
    x_129 = 'b000001011;
    x_130 = 'b000001011;
    x_131 = 'b000001110;
    x_132 = 'b000000001;
    x_133 = 'b111101110;
    x_134 = 'b111100111;
    x_135 = 'b000001101;
    x_136 = 'b000010000;
    x_137 = 'b000010001;
    x_138 = 'b000010011;
    x_139 = 'b000010001;
    x_140 = 'b111111101;
    x_141 = 'b111110000;
    x_142 = 'b000010101;
    x_143 = 'b000011001;
    x_144 = 'b000010011;
    x_145 = 'b000010001;
    x_146 = 'b000010000;
    x_147 = 'b000001110;
    x_148 = 'b111111111;
    x_149 = 'b000000011;
    x_150 = 'b111110111;
    x_151 = 'b111111011;
    x_152 = 'b000001001;
    x_153 = 'b000001011;
    x_154 = 'b111111101;
    x_155 = 'b111110011;
    x_156 = 'b111111011;
    x_157 = 'b000001111;
    x_158 = 'b000000111;
    x_159 = 'b000000100;
    x_160 = 'b000010010;
    x_161 = 'b000001011;
    x_162 = 'b000000010;
    x_163 = 'b111111110;
    x_164 = 'b111110010;
    x_165 = 'b000000110;
    x_166 = 'b000011100;
    x_167 = 'b111110000;
    x_168 = 'b000100000;
    x_169 = 'b000001100;
    x_170 = 'b000011001;
    x_171 = 'b000011011;
    x_172 = 'b000010111;
    x_173 = 'b000001100;
    x_174 = 'b000011001;
    x_175 = 'b000011101;
    x_176 = 'b000010001;
    x_177 = 'b000011010;
    x_178 = 'b000011011;
    x_179 = 'b000011001;
    x_180 = 'b000010001;
    x_181 = 'b000010000;
    x_182 = 'b000001101;
    x_183 = 'b000011000;
    x_184 = 'b000100001;
    x_185 = 'b000011101;
    x_186 = 'b000010010;
    x_187 = 'b000000101;
    x_188 = 'b000010001;
    x_189 = 'b000001111;
    x_190 = 'b111110011;
    x_191 = 'b000001000;
    x_192 = 'b000010100;
    x_193 = 'b000001011;
    x_194 = 'b000001011;
    x_195 = 'b000001110;
    x_196 = 'b000000001;
    x_197 = 'b111101110;
    x_198 = 'b111100111;
    x_199 = 'b000001101;
    x_200 = 'b000010000;
    x_201 = 'b000010001;
    x_202 = 'b000010011;
    x_203 = 'b000010001;
    x_204 = 'b111111101;
    x_205 = 'b111110000;
    x_206 = 'b000010101;
    x_207 = 'b000011001;
    x_208 = 'b000010011;
    x_209 = 'b000010001;
    x_210 = 'b000010000;
    x_211 = 'b000001110;
    x_212 = 'b111111111;
    x_213 = 'b000000011;
    x_214 = 'b111110111;
    x_215 = 'b111111011;
    x_216 = 'b000001001;
    x_217 = 'b000001011;
    x_218 = 'b111111101;
    x_219 = 'b111110011;
    x_220 = 'b111111011;
    x_221 = 'b000001111;
    x_222 = 'b000000111;
    x_223 = 'b000000100;
    x_224 = 'b000010010;
    x_225 = 'b000001011;
    x_226 = 'b000000010;
    x_227 = 'b111111110;
    x_228 = 'b111110010;
    x_229 = 'b000000110;
    x_230 = 'b000011100;
    x_231 = 'b111110000;
    x_232 = 'b000100000;
    x_233 = 'b000001100;
    x_234 = 'b000011001;
    x_235 = 'b000011011;
    x_236 = 'b000010111;
    x_237 = 'b000001100;
    x_238 = 'b000011001;
    x_239 = 'b000011101;
    x_240 = 'b000010001;
    x_241 = 'b000011010;
    x_242 = 'b000011011;
    x_243 = 'b000011001;
    x_244 = 'b000010001;
    x_245 = 'b000010000;
    x_246 = 'b000001101;
    x_247 = 'b000011000;
    x_248 = 'b000100001;
    x_249 = 'b000011101;
    x_250 = 'b000010010;
    x_251 = 'b000000101;
    x_252 = 'b000010001;
    x_253 = 'b000001111;
    x_254 = 'b111110011;
    x_255 = 'b000001000;

    h_0 = 'b000010100;
    h_1 = 'b000001011;
    h_2 = 'b000001011;
    h_3 = 'b000001110;
    h_4 = 'b000000001;
    h_5 = 'b111101110;
    h_6 = 'b111100111;
    h_7 = 'b000001101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000011010;
    x_1 = 'b000011001;
    x_2 = 'b000011100;
    x_3 = 'b000100000;
    x_4 = 'b000011001;
    x_5 = 'b000000101;
    x_6 = 'b111111101;
    x_7 = 'b000010111;
    x_8 = 'b000011101;
    x_9 = 'b000011110;
    x_10 = 'b000100011;
    x_11 = 'b000100100;
    x_12 = 'b000010111;
    x_13 = 'b000001001;
    x_14 = 'b000100101;
    x_15 = 'b000100100;
    x_16 = 'b000100011;
    x_17 = 'b000100001;
    x_18 = 'b000100001;
    x_19 = 'b000100000;
    x_20 = 'b000010011;
    x_21 = 'b000001000;
    x_22 = 'b000000001;
    x_23 = 'b000000010;
    x_24 = 'b000001001;
    x_25 = 'b000001100;
    x_26 = 'b000001000;
    x_27 = 'b111111100;
    x_28 = 'b000000000;
    x_29 = 'b000001110;
    x_30 = 'b000000111;
    x_31 = 'b000001011;
    x_32 = 'b000010110;
    x_33 = 'b000010000;
    x_34 = 'b000001010;
    x_35 = 'b000000010;
    x_36 = 'b111111000;
    x_37 = 'b000001011;
    x_38 = 'b000001101;
    x_39 = 'b111111000;
    x_40 = 'b000001111;
    x_41 = 'b000001100;
    x_42 = 'b000011001;
    x_43 = 'b000011110;
    x_44 = 'b000010101;
    x_45 = 'b000010101;
    x_46 = 'b000011111;
    x_47 = 'b000100010;
    x_48 = 'b000010010;
    x_49 = 'b000011110;
    x_50 = 'b000011110;
    x_51 = 'b000011101;
    x_52 = 'b000010111;
    x_53 = 'b000010011;
    x_54 = 'b000001010;
    x_55 = 'b000011101;
    x_56 = 'b000100101;
    x_57 = 'b000100000;
    x_58 = 'b000010110;
    x_59 = 'b000000110;
    x_60 = 'b000011001;
    x_61 = 'b000011001;
    x_62 = 'b111111111;
    x_63 = 'b000010101;
    x_64 = 'b000011010;
    x_65 = 'b000011001;
    x_66 = 'b000011100;
    x_67 = 'b000100000;
    x_68 = 'b000011001;
    x_69 = 'b000000101;
    x_70 = 'b111111101;
    x_71 = 'b000010111;
    x_72 = 'b000011101;
    x_73 = 'b000011110;
    x_74 = 'b000100011;
    x_75 = 'b000100100;
    x_76 = 'b000010111;
    x_77 = 'b000001001;
    x_78 = 'b000100101;
    x_79 = 'b000100100;
    x_80 = 'b000100011;
    x_81 = 'b000100001;
    x_82 = 'b000100001;
    x_83 = 'b000100000;
    x_84 = 'b000010011;
    x_85 = 'b000001000;
    x_86 = 'b000000001;
    x_87 = 'b000000010;
    x_88 = 'b000001001;
    x_89 = 'b000001100;
    x_90 = 'b000001000;
    x_91 = 'b111111100;
    x_92 = 'b000000000;
    x_93 = 'b000001110;
    x_94 = 'b000000111;
    x_95 = 'b000001011;
    x_96 = 'b000010110;
    x_97 = 'b000010000;
    x_98 = 'b000001010;
    x_99 = 'b000000010;
    x_100 = 'b111111000;
    x_101 = 'b000001011;
    x_102 = 'b000001101;
    x_103 = 'b111111000;
    x_104 = 'b000001111;
    x_105 = 'b000001100;
    x_106 = 'b000011001;
    x_107 = 'b000011110;
    x_108 = 'b000010101;
    x_109 = 'b000010101;
    x_110 = 'b000011111;
    x_111 = 'b000100010;
    x_112 = 'b000010010;
    x_113 = 'b000011110;
    x_114 = 'b000011110;
    x_115 = 'b000011101;
    x_116 = 'b000010111;
    x_117 = 'b000010011;
    x_118 = 'b000001010;
    x_119 = 'b000011101;
    x_120 = 'b000100101;
    x_121 = 'b000100000;
    x_122 = 'b000010110;
    x_123 = 'b000000110;
    x_124 = 'b000011001;
    x_125 = 'b000011001;
    x_126 = 'b111111111;
    x_127 = 'b000010101;
    x_128 = 'b000011010;
    x_129 = 'b000011001;
    x_130 = 'b000011100;
    x_131 = 'b000100000;
    x_132 = 'b000011001;
    x_133 = 'b000000101;
    x_134 = 'b111111101;
    x_135 = 'b000010111;
    x_136 = 'b000011101;
    x_137 = 'b000011110;
    x_138 = 'b000100011;
    x_139 = 'b000100100;
    x_140 = 'b000010111;
    x_141 = 'b000001001;
    x_142 = 'b000100101;
    x_143 = 'b000100100;
    x_144 = 'b000100011;
    x_145 = 'b000100001;
    x_146 = 'b000100001;
    x_147 = 'b000100000;
    x_148 = 'b000010011;
    x_149 = 'b000001000;
    x_150 = 'b000000001;
    x_151 = 'b000000010;
    x_152 = 'b000001001;
    x_153 = 'b000001100;
    x_154 = 'b000001000;
    x_155 = 'b111111100;
    x_156 = 'b000000000;
    x_157 = 'b000001110;
    x_158 = 'b000000111;
    x_159 = 'b000001011;
    x_160 = 'b000010110;
    x_161 = 'b000010000;
    x_162 = 'b000001010;
    x_163 = 'b000000010;
    x_164 = 'b111111000;
    x_165 = 'b000001011;
    x_166 = 'b000001101;
    x_167 = 'b111111000;
    x_168 = 'b000001111;
    x_169 = 'b000001100;
    x_170 = 'b000011001;
    x_171 = 'b000011110;
    x_172 = 'b000010101;
    x_173 = 'b000010101;
    x_174 = 'b000011111;
    x_175 = 'b000100010;
    x_176 = 'b000010010;
    x_177 = 'b000011110;
    x_178 = 'b000011110;
    x_179 = 'b000011101;
    x_180 = 'b000010111;
    x_181 = 'b000010011;
    x_182 = 'b000001010;
    x_183 = 'b000011101;
    x_184 = 'b000100101;
    x_185 = 'b000100000;
    x_186 = 'b000010110;
    x_187 = 'b000000110;
    x_188 = 'b000011001;
    x_189 = 'b000011001;
    x_190 = 'b111111111;
    x_191 = 'b000010101;
    x_192 = 'b000011010;
    x_193 = 'b000011001;
    x_194 = 'b000011100;
    x_195 = 'b000100000;
    x_196 = 'b000011001;
    x_197 = 'b000000101;
    x_198 = 'b111111101;
    x_199 = 'b000010111;
    x_200 = 'b000011101;
    x_201 = 'b000011110;
    x_202 = 'b000100011;
    x_203 = 'b000100100;
    x_204 = 'b000010111;
    x_205 = 'b000001001;
    x_206 = 'b000100101;
    x_207 = 'b000100100;
    x_208 = 'b000100011;
    x_209 = 'b000100001;
    x_210 = 'b000100001;
    x_211 = 'b000100000;
    x_212 = 'b000010011;
    x_213 = 'b000001000;
    x_214 = 'b000000001;
    x_215 = 'b000000010;
    x_216 = 'b000001001;
    x_217 = 'b000001100;
    x_218 = 'b000001000;
    x_219 = 'b111111100;
    x_220 = 'b000000000;
    x_221 = 'b000001110;
    x_222 = 'b000000111;
    x_223 = 'b000001011;
    x_224 = 'b000010110;
    x_225 = 'b000010000;
    x_226 = 'b000001010;
    x_227 = 'b000000010;
    x_228 = 'b111111000;
    x_229 = 'b000001011;
    x_230 = 'b000001101;
    x_231 = 'b111111000;
    x_232 = 'b000001111;
    x_233 = 'b000001100;
    x_234 = 'b000011001;
    x_235 = 'b000011110;
    x_236 = 'b000010101;
    x_237 = 'b000010101;
    x_238 = 'b000011111;
    x_239 = 'b000100010;
    x_240 = 'b000010010;
    x_241 = 'b000011110;
    x_242 = 'b000011110;
    x_243 = 'b000011101;
    x_244 = 'b000010111;
    x_245 = 'b000010011;
    x_246 = 'b000001010;
    x_247 = 'b000011101;
    x_248 = 'b000100101;
    x_249 = 'b000100000;
    x_250 = 'b000010110;
    x_251 = 'b000000110;
    x_252 = 'b000011001;
    x_253 = 'b000011001;
    x_254 = 'b111111111;
    x_255 = 'b000010101;

    h_0 = 'b000011010;
    h_1 = 'b000011001;
    h_2 = 'b000011100;
    h_3 = 'b000100000;
    h_4 = 'b000011001;
    h_5 = 'b000000101;
    h_6 = 'b111111101;
    h_7 = 'b000010111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000000101;
    x_1 = 'b000000111;
    x_2 = 'b111101000;
    x_3 = 'b111110000;
    x_4 = 'b111101101;
    x_5 = 'b111101001;
    x_6 = 'b111110100;
    x_7 = 'b000010001;
    x_8 = 'b000000001;
    x_9 = 'b111110100;
    x_10 = 'b111101100;
    x_11 = 'b111011111;
    x_12 = 'b111100010;
    x_13 = 'b111100110;
    x_14 = 'b000011000;
    x_15 = 'b000001001;
    x_16 = 'b111111000;
    x_17 = 'b111110000;
    x_18 = 'b111011111;
    x_19 = 'b111100000;
    x_20 = 'b111101010;
    x_21 = 'b111111111;
    x_22 = 'b000001000;
    x_23 = 'b000001010;
    x_24 = 'b000000110;
    x_25 = 'b000000101;
    x_26 = 'b111110001;
    x_27 = 'b111111000;
    x_28 = 'b000001111;
    x_29 = 'b000000011;
    x_30 = 'b000010010;
    x_31 = 'b111111110;
    x_32 = 'b111111001;
    x_33 = 'b111110101;
    x_34 = 'b111110011;
    x_35 = 'b111101110;
    x_36 = 'b111111110;
    x_37 = 'b111011001;
    x_38 = 'b000001001;
    x_39 = 'b000000100;
    x_40 = 'b000010001;
    x_41 = 'b000000111;
    x_42 = 'b000011000;
    x_43 = 'b111111110;
    x_44 = 'b000011100;
    x_45 = 'b000000000;
    x_46 = 'b000011011;
    x_47 = 'b000010110;
    x_48 = 'b000001110;
    x_49 = 'b000000101;
    x_50 = 'b111110101;
    x_51 = 'b111101111;
    x_52 = 'b111110001;
    x_53 = 'b111110111;
    x_54 = 'b000001010;
    x_55 = 'b000001110;
    x_56 = 'b000010101;
    x_57 = 'b111111010;
    x_58 = 'b111111001;
    x_59 = 'b000010101;
    x_60 = 'b000000011;
    x_61 = 'b111111010;
    x_62 = 'b111111101;
    x_63 = 'b000001000;
    x_64 = 'b000000101;
    x_65 = 'b000000111;
    x_66 = 'b111101000;
    x_67 = 'b111110000;
    x_68 = 'b111101101;
    x_69 = 'b111101001;
    x_70 = 'b111110100;
    x_71 = 'b000010001;
    x_72 = 'b000000001;
    x_73 = 'b111110100;
    x_74 = 'b111101100;
    x_75 = 'b111011111;
    x_76 = 'b111100010;
    x_77 = 'b111100110;
    x_78 = 'b000011000;
    x_79 = 'b000001001;
    x_80 = 'b111111000;
    x_81 = 'b111110000;
    x_82 = 'b111011111;
    x_83 = 'b111100000;
    x_84 = 'b111101010;
    x_85 = 'b111111111;
    x_86 = 'b000001000;
    x_87 = 'b000001010;
    x_88 = 'b000000110;
    x_89 = 'b000000101;
    x_90 = 'b111110001;
    x_91 = 'b111111000;
    x_92 = 'b000001111;
    x_93 = 'b000000011;
    x_94 = 'b000010010;
    x_95 = 'b111111110;
    x_96 = 'b111111001;
    x_97 = 'b111110101;
    x_98 = 'b111110011;
    x_99 = 'b111101110;
    x_100 = 'b111111110;
    x_101 = 'b111011001;
    x_102 = 'b000001001;
    x_103 = 'b000000100;
    x_104 = 'b000010001;
    x_105 = 'b000000111;
    x_106 = 'b000011000;
    x_107 = 'b111111110;
    x_108 = 'b000011100;
    x_109 = 'b000000000;
    x_110 = 'b000011011;
    x_111 = 'b000010110;
    x_112 = 'b000001110;
    x_113 = 'b000000101;
    x_114 = 'b111110101;
    x_115 = 'b111101111;
    x_116 = 'b111110001;
    x_117 = 'b111110111;
    x_118 = 'b000001010;
    x_119 = 'b000001110;
    x_120 = 'b000010101;
    x_121 = 'b111111010;
    x_122 = 'b111111001;
    x_123 = 'b000010101;
    x_124 = 'b000000011;
    x_125 = 'b111111010;
    x_126 = 'b111111101;
    x_127 = 'b000001000;
    x_128 = 'b000000101;
    x_129 = 'b000000111;
    x_130 = 'b111101000;
    x_131 = 'b111110000;
    x_132 = 'b111101101;
    x_133 = 'b111101001;
    x_134 = 'b111110100;
    x_135 = 'b000010001;
    x_136 = 'b000000001;
    x_137 = 'b111110100;
    x_138 = 'b111101100;
    x_139 = 'b111011111;
    x_140 = 'b111100010;
    x_141 = 'b111100110;
    x_142 = 'b000011000;
    x_143 = 'b000001001;
    x_144 = 'b111111000;
    x_145 = 'b111110000;
    x_146 = 'b111011111;
    x_147 = 'b111100000;
    x_148 = 'b111101010;
    x_149 = 'b111111111;
    x_150 = 'b000001000;
    x_151 = 'b000001010;
    x_152 = 'b000000110;
    x_153 = 'b000000101;
    x_154 = 'b111110001;
    x_155 = 'b111111000;
    x_156 = 'b000001111;
    x_157 = 'b000000011;
    x_158 = 'b000010010;
    x_159 = 'b111111110;
    x_160 = 'b111111001;
    x_161 = 'b111110101;
    x_162 = 'b111110011;
    x_163 = 'b111101110;
    x_164 = 'b111111110;
    x_165 = 'b111011001;
    x_166 = 'b000001001;
    x_167 = 'b000000100;
    x_168 = 'b000010001;
    x_169 = 'b000000111;
    x_170 = 'b000011000;
    x_171 = 'b111111110;
    x_172 = 'b000011100;
    x_173 = 'b000000000;
    x_174 = 'b000011011;
    x_175 = 'b000010110;
    x_176 = 'b000001110;
    x_177 = 'b000000101;
    x_178 = 'b111110101;
    x_179 = 'b111101111;
    x_180 = 'b111110001;
    x_181 = 'b111110111;
    x_182 = 'b000001010;
    x_183 = 'b000001110;
    x_184 = 'b000010101;
    x_185 = 'b111111010;
    x_186 = 'b111111001;
    x_187 = 'b000010101;
    x_188 = 'b000000011;
    x_189 = 'b111111010;
    x_190 = 'b111111101;
    x_191 = 'b000001000;
    x_192 = 'b000000101;
    x_193 = 'b000000111;
    x_194 = 'b111101000;
    x_195 = 'b111110000;
    x_196 = 'b111101101;
    x_197 = 'b111101001;
    x_198 = 'b111110100;
    x_199 = 'b000010001;
    x_200 = 'b000000001;
    x_201 = 'b111110100;
    x_202 = 'b111101100;
    x_203 = 'b111011111;
    x_204 = 'b111100010;
    x_205 = 'b111100110;
    x_206 = 'b000011000;
    x_207 = 'b000001001;
    x_208 = 'b111111000;
    x_209 = 'b111110000;
    x_210 = 'b111011111;
    x_211 = 'b111100000;
    x_212 = 'b111101010;
    x_213 = 'b111111111;
    x_214 = 'b000001000;
    x_215 = 'b000001010;
    x_216 = 'b000000110;
    x_217 = 'b000000101;
    x_218 = 'b111110001;
    x_219 = 'b111111000;
    x_220 = 'b000001111;
    x_221 = 'b000000011;
    x_222 = 'b000010010;
    x_223 = 'b111111110;
    x_224 = 'b111111001;
    x_225 = 'b111110101;
    x_226 = 'b111110011;
    x_227 = 'b111101110;
    x_228 = 'b111111110;
    x_229 = 'b111011001;
    x_230 = 'b000001001;
    x_231 = 'b000000100;
    x_232 = 'b000010001;
    x_233 = 'b000000111;
    x_234 = 'b000011000;
    x_235 = 'b111111110;
    x_236 = 'b000011100;
    x_237 = 'b000000000;
    x_238 = 'b000011011;
    x_239 = 'b000010110;
    x_240 = 'b000001110;
    x_241 = 'b000000101;
    x_242 = 'b111110101;
    x_243 = 'b111101111;
    x_244 = 'b111110001;
    x_245 = 'b111110111;
    x_246 = 'b000001010;
    x_247 = 'b000001110;
    x_248 = 'b000010101;
    x_249 = 'b111111010;
    x_250 = 'b111111001;
    x_251 = 'b000010101;
    x_252 = 'b000000011;
    x_253 = 'b111111010;
    x_254 = 'b111111101;
    x_255 = 'b000001000;

    h_0 = 'b000000101;
    h_1 = 'b000000111;
    h_2 = 'b111101000;
    h_3 = 'b111110000;
    h_4 = 'b111101101;
    h_5 = 'b111101001;
    h_6 = 'b111110100;
    h_7 = 'b000010001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000010101;
    x_1 = 'b000011000;
    x_2 = 'b000000000;
    x_3 = 'b000000101;
    x_4 = 'b111111101;
    x_5 = 'b111111001;
    x_6 = 'b111111110;
    x_7 = 'b000100110;
    x_8 = 'b000010010;
    x_9 = 'b000000111;
    x_10 = 'b000000000;
    x_11 = 'b111110110;
    x_12 = 'b111111000;
    x_13 = 'b111111011;
    x_14 = 'b000011000;
    x_15 = 'b000010100;
    x_16 = 'b000001000;
    x_17 = 'b000000110;
    x_18 = 'b111110110;
    x_19 = 'b111111010;
    x_20 = 'b000000000;
    x_21 = 'b000000001;
    x_22 = 'b000001010;
    x_23 = 'b000001101;
    x_24 = 'b000001011;
    x_25 = 'b000001011;
    x_26 = 'b111111100;
    x_27 = 'b111111111;
    x_28 = 'b000010000;
    x_29 = 'b000001111;
    x_30 = 'b000011110;
    x_31 = 'b000001000;
    x_32 = 'b000001001;
    x_33 = 'b000000010;
    x_34 = 'b111111101;
    x_35 = 'b111111011;
    x_36 = 'b000000010;
    x_37 = 'b111010101;
    x_38 = 'b000011101;
    x_39 = 'b000000110;
    x_40 = 'b000100111;
    x_41 = 'b111110011;
    x_42 = 'b000011001;
    x_43 = 'b000010100;
    x_44 = 'b000011100;
    x_45 = 'b000001010;
    x_46 = 'b000010000;
    x_47 = 'b000010011;
    x_48 = 'b000001110;
    x_49 = 'b000001001;
    x_50 = 'b000000010;
    x_51 = 'b000000001;
    x_52 = 'b000000010;
    x_53 = 'b000000100;
    x_54 = 'b000010010;
    x_55 = 'b000001001;
    x_56 = 'b000001111;
    x_57 = 'b000000000;
    x_58 = 'b000001010;
    x_59 = 'b000010110;
    x_60 = 'b111111100;
    x_61 = 'b111111101;
    x_62 = 'b000001001;
    x_63 = 'b111110111;
    x_64 = 'b000010101;
    x_65 = 'b000011000;
    x_66 = 'b000000000;
    x_67 = 'b000000101;
    x_68 = 'b111111101;
    x_69 = 'b111111001;
    x_70 = 'b111111110;
    x_71 = 'b000100110;
    x_72 = 'b000010010;
    x_73 = 'b000000111;
    x_74 = 'b000000000;
    x_75 = 'b111110110;
    x_76 = 'b111111000;
    x_77 = 'b111111011;
    x_78 = 'b000011000;
    x_79 = 'b000010100;
    x_80 = 'b000001000;
    x_81 = 'b000000110;
    x_82 = 'b111110110;
    x_83 = 'b111111010;
    x_84 = 'b000000000;
    x_85 = 'b000000001;
    x_86 = 'b000001010;
    x_87 = 'b000001101;
    x_88 = 'b000001011;
    x_89 = 'b000001011;
    x_90 = 'b111111100;
    x_91 = 'b111111111;
    x_92 = 'b000010000;
    x_93 = 'b000001111;
    x_94 = 'b000011110;
    x_95 = 'b000001000;
    x_96 = 'b000001001;
    x_97 = 'b000000010;
    x_98 = 'b111111101;
    x_99 = 'b111111011;
    x_100 = 'b000000010;
    x_101 = 'b111010101;
    x_102 = 'b000011101;
    x_103 = 'b000000110;
    x_104 = 'b000100111;
    x_105 = 'b111110011;
    x_106 = 'b000011001;
    x_107 = 'b000010100;
    x_108 = 'b000011100;
    x_109 = 'b000001010;
    x_110 = 'b000010000;
    x_111 = 'b000010011;
    x_112 = 'b000001110;
    x_113 = 'b000001001;
    x_114 = 'b000000010;
    x_115 = 'b000000001;
    x_116 = 'b000000010;
    x_117 = 'b000000100;
    x_118 = 'b000010010;
    x_119 = 'b000001001;
    x_120 = 'b000001111;
    x_121 = 'b000000000;
    x_122 = 'b000001010;
    x_123 = 'b000010110;
    x_124 = 'b111111100;
    x_125 = 'b111111101;
    x_126 = 'b000001001;
    x_127 = 'b111110111;
    x_128 = 'b000010101;
    x_129 = 'b000011000;
    x_130 = 'b000000000;
    x_131 = 'b000000101;
    x_132 = 'b111111101;
    x_133 = 'b111111001;
    x_134 = 'b111111110;
    x_135 = 'b000100110;
    x_136 = 'b000010010;
    x_137 = 'b000000111;
    x_138 = 'b000000000;
    x_139 = 'b111110110;
    x_140 = 'b111111000;
    x_141 = 'b111111011;
    x_142 = 'b000011000;
    x_143 = 'b000010100;
    x_144 = 'b000001000;
    x_145 = 'b000000110;
    x_146 = 'b111110110;
    x_147 = 'b111111010;
    x_148 = 'b000000000;
    x_149 = 'b000000001;
    x_150 = 'b000001010;
    x_151 = 'b000001101;
    x_152 = 'b000001011;
    x_153 = 'b000001011;
    x_154 = 'b111111100;
    x_155 = 'b111111111;
    x_156 = 'b000010000;
    x_157 = 'b000001111;
    x_158 = 'b000011110;
    x_159 = 'b000001000;
    x_160 = 'b000001001;
    x_161 = 'b000000010;
    x_162 = 'b111111101;
    x_163 = 'b111111011;
    x_164 = 'b000000010;
    x_165 = 'b111010101;
    x_166 = 'b000011101;
    x_167 = 'b000000110;
    x_168 = 'b000100111;
    x_169 = 'b111110011;
    x_170 = 'b000011001;
    x_171 = 'b000010100;
    x_172 = 'b000011100;
    x_173 = 'b000001010;
    x_174 = 'b000010000;
    x_175 = 'b000010011;
    x_176 = 'b000001110;
    x_177 = 'b000001001;
    x_178 = 'b000000010;
    x_179 = 'b000000001;
    x_180 = 'b000000010;
    x_181 = 'b000000100;
    x_182 = 'b000010010;
    x_183 = 'b000001001;
    x_184 = 'b000001111;
    x_185 = 'b000000000;
    x_186 = 'b000001010;
    x_187 = 'b000010110;
    x_188 = 'b111111100;
    x_189 = 'b111111101;
    x_190 = 'b000001001;
    x_191 = 'b111110111;
    x_192 = 'b000010101;
    x_193 = 'b000011000;
    x_194 = 'b000000000;
    x_195 = 'b000000101;
    x_196 = 'b111111101;
    x_197 = 'b111111001;
    x_198 = 'b111111110;
    x_199 = 'b000100110;
    x_200 = 'b000010010;
    x_201 = 'b000000111;
    x_202 = 'b000000000;
    x_203 = 'b111110110;
    x_204 = 'b111111000;
    x_205 = 'b111111011;
    x_206 = 'b000011000;
    x_207 = 'b000010100;
    x_208 = 'b000001000;
    x_209 = 'b000000110;
    x_210 = 'b111110110;
    x_211 = 'b111111010;
    x_212 = 'b000000000;
    x_213 = 'b000000001;
    x_214 = 'b000001010;
    x_215 = 'b000001101;
    x_216 = 'b000001011;
    x_217 = 'b000001011;
    x_218 = 'b111111100;
    x_219 = 'b111111111;
    x_220 = 'b000010000;
    x_221 = 'b000001111;
    x_222 = 'b000011110;
    x_223 = 'b000001000;
    x_224 = 'b000001001;
    x_225 = 'b000000010;
    x_226 = 'b111111101;
    x_227 = 'b111111011;
    x_228 = 'b000000010;
    x_229 = 'b111010101;
    x_230 = 'b000011101;
    x_231 = 'b000000110;
    x_232 = 'b000100111;
    x_233 = 'b111110011;
    x_234 = 'b000011001;
    x_235 = 'b000010100;
    x_236 = 'b000011100;
    x_237 = 'b000001010;
    x_238 = 'b000010000;
    x_239 = 'b000010011;
    x_240 = 'b000001110;
    x_241 = 'b000001001;
    x_242 = 'b000000010;
    x_243 = 'b000000001;
    x_244 = 'b000000010;
    x_245 = 'b000000100;
    x_246 = 'b000010010;
    x_247 = 'b000001001;
    x_248 = 'b000001111;
    x_249 = 'b000000000;
    x_250 = 'b000001010;
    x_251 = 'b000010110;
    x_252 = 'b111111100;
    x_253 = 'b111111101;
    x_254 = 'b000001001;
    x_255 = 'b111110111;

    h_0 = 'b000010101;
    h_1 = 'b000011000;
    h_2 = 'b000000000;
    h_3 = 'b000000101;
    h_4 = 'b111111101;
    h_5 = 'b111111001;
    h_6 = 'b111111110;
    h_7 = 'b000100110;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000100101;
    x_1 = 'b000100001;
    x_2 = 'b000001010;
    x_3 = 'b000001011;
    x_4 = 'b000000001;
    x_5 = 'b111111101;
    x_6 = 'b111111101;
    x_7 = 'b000101010;
    x_8 = 'b000010100;
    x_9 = 'b000001100;
    x_10 = 'b000000100;
    x_11 = 'b000000001;
    x_12 = 'b000000010;
    x_13 = 'b111111011;
    x_14 = 'b000011100;
    x_15 = 'b000010110;
    x_16 = 'b000001011;
    x_17 = 'b000001101;
    x_18 = 'b000000101;
    x_19 = 'b000001011;
    x_20 = 'b000001110;
    x_21 = 'b000010100;
    x_22 = 'b000011001;
    x_23 = 'b000010110;
    x_24 = 'b000100100;
    x_25 = 'b000100010;
    x_26 = 'b000001000;
    x_27 = 'b000000110;
    x_28 = 'b000010011;
    x_29 = 'b000101000;
    x_30 = 'b000110111;
    x_31 = 'b000010101;
    x_32 = 'b000011000;
    x_33 = 'b000001111;
    x_34 = 'b000001001;
    x_35 = 'b000000110;
    x_36 = 'b000000011;
    x_37 = 'b111001110;
    x_38 = 'b000111001;
    x_39 = 'b111111110;
    x_40 = 'b000110111;
    x_41 = 'b111100001;
    x_42 = 'b000101110;
    x_43 = 'b000000001;
    x_44 = 'b000101001;
    x_45 = 'b000101010;
    x_46 = 'b000011110;
    x_47 = 'b000100000;
    x_48 = 'b000100000;
    x_49 = 'b000011011;
    x_50 = 'b000011100;
    x_51 = 'b000100011;
    x_52 = 'b000101000;
    x_53 = 'b000101001;
    x_54 = 'b000110000;
    x_55 = 'b000010111;
    x_56 = 'b000011101;
    x_57 = 'b000011100;
    x_58 = 'b000110000;
    x_59 = 'b000101110;
    x_60 = 'b111111100;
    x_61 = 'b000000100;
    x_62 = 'b000010000;
    x_63 = 'b111101000;
    x_64 = 'b000100101;
    x_65 = 'b000100001;
    x_66 = 'b000001010;
    x_67 = 'b000001011;
    x_68 = 'b000000001;
    x_69 = 'b111111101;
    x_70 = 'b111111101;
    x_71 = 'b000101010;
    x_72 = 'b000010100;
    x_73 = 'b000001100;
    x_74 = 'b000000100;
    x_75 = 'b000000001;
    x_76 = 'b000000010;
    x_77 = 'b111111011;
    x_78 = 'b000011100;
    x_79 = 'b000010110;
    x_80 = 'b000001011;
    x_81 = 'b000001101;
    x_82 = 'b000000101;
    x_83 = 'b000001011;
    x_84 = 'b000001110;
    x_85 = 'b000010100;
    x_86 = 'b000011001;
    x_87 = 'b000010110;
    x_88 = 'b000100100;
    x_89 = 'b000100010;
    x_90 = 'b000001000;
    x_91 = 'b000000110;
    x_92 = 'b000010011;
    x_93 = 'b000101000;
    x_94 = 'b000110111;
    x_95 = 'b000010101;
    x_96 = 'b000011000;
    x_97 = 'b000001111;
    x_98 = 'b000001001;
    x_99 = 'b000000110;
    x_100 = 'b000000011;
    x_101 = 'b111001110;
    x_102 = 'b000111001;
    x_103 = 'b111111110;
    x_104 = 'b000110111;
    x_105 = 'b111100001;
    x_106 = 'b000101110;
    x_107 = 'b000000001;
    x_108 = 'b000101001;
    x_109 = 'b000101010;
    x_110 = 'b000011110;
    x_111 = 'b000100000;
    x_112 = 'b000100000;
    x_113 = 'b000011011;
    x_114 = 'b000011100;
    x_115 = 'b000100011;
    x_116 = 'b000101000;
    x_117 = 'b000101001;
    x_118 = 'b000110000;
    x_119 = 'b000010111;
    x_120 = 'b000011101;
    x_121 = 'b000011100;
    x_122 = 'b000110000;
    x_123 = 'b000101110;
    x_124 = 'b111111100;
    x_125 = 'b000000100;
    x_126 = 'b000010000;
    x_127 = 'b111101000;
    x_128 = 'b000100101;
    x_129 = 'b000100001;
    x_130 = 'b000001010;
    x_131 = 'b000001011;
    x_132 = 'b000000001;
    x_133 = 'b111111101;
    x_134 = 'b111111101;
    x_135 = 'b000101010;
    x_136 = 'b000010100;
    x_137 = 'b000001100;
    x_138 = 'b000000100;
    x_139 = 'b000000001;
    x_140 = 'b000000010;
    x_141 = 'b111111011;
    x_142 = 'b000011100;
    x_143 = 'b000010110;
    x_144 = 'b000001011;
    x_145 = 'b000001101;
    x_146 = 'b000000101;
    x_147 = 'b000001011;
    x_148 = 'b000001110;
    x_149 = 'b000010100;
    x_150 = 'b000011001;
    x_151 = 'b000010110;
    x_152 = 'b000100100;
    x_153 = 'b000100010;
    x_154 = 'b000001000;
    x_155 = 'b000000110;
    x_156 = 'b000010011;
    x_157 = 'b000101000;
    x_158 = 'b000110111;
    x_159 = 'b000010101;
    x_160 = 'b000011000;
    x_161 = 'b000001111;
    x_162 = 'b000001001;
    x_163 = 'b000000110;
    x_164 = 'b000000011;
    x_165 = 'b111001110;
    x_166 = 'b000111001;
    x_167 = 'b111111110;
    x_168 = 'b000110111;
    x_169 = 'b111100001;
    x_170 = 'b000101110;
    x_171 = 'b000000001;
    x_172 = 'b000101001;
    x_173 = 'b000101010;
    x_174 = 'b000011110;
    x_175 = 'b000100000;
    x_176 = 'b000100000;
    x_177 = 'b000011011;
    x_178 = 'b000011100;
    x_179 = 'b000100011;
    x_180 = 'b000101000;
    x_181 = 'b000101001;
    x_182 = 'b000110000;
    x_183 = 'b000010111;
    x_184 = 'b000011101;
    x_185 = 'b000011100;
    x_186 = 'b000110000;
    x_187 = 'b000101110;
    x_188 = 'b111111100;
    x_189 = 'b000000100;
    x_190 = 'b000010000;
    x_191 = 'b111101000;
    x_192 = 'b000100101;
    x_193 = 'b000100001;
    x_194 = 'b000001010;
    x_195 = 'b000001011;
    x_196 = 'b000000001;
    x_197 = 'b111111101;
    x_198 = 'b111111101;
    x_199 = 'b000101010;
    x_200 = 'b000010100;
    x_201 = 'b000001100;
    x_202 = 'b000000100;
    x_203 = 'b000000001;
    x_204 = 'b000000010;
    x_205 = 'b111111011;
    x_206 = 'b000011100;
    x_207 = 'b000010110;
    x_208 = 'b000001011;
    x_209 = 'b000001101;
    x_210 = 'b000000101;
    x_211 = 'b000001011;
    x_212 = 'b000001110;
    x_213 = 'b000010100;
    x_214 = 'b000011001;
    x_215 = 'b000010110;
    x_216 = 'b000100100;
    x_217 = 'b000100010;
    x_218 = 'b000001000;
    x_219 = 'b000000110;
    x_220 = 'b000010011;
    x_221 = 'b000101000;
    x_222 = 'b000110111;
    x_223 = 'b000010101;
    x_224 = 'b000011000;
    x_225 = 'b000001111;
    x_226 = 'b000001001;
    x_227 = 'b000000110;
    x_228 = 'b000000011;
    x_229 = 'b111001110;
    x_230 = 'b000111001;
    x_231 = 'b111111110;
    x_232 = 'b000110111;
    x_233 = 'b111100001;
    x_234 = 'b000101110;
    x_235 = 'b000000001;
    x_236 = 'b000101001;
    x_237 = 'b000101010;
    x_238 = 'b000011110;
    x_239 = 'b000100000;
    x_240 = 'b000100000;
    x_241 = 'b000011011;
    x_242 = 'b000011100;
    x_243 = 'b000100011;
    x_244 = 'b000101000;
    x_245 = 'b000101001;
    x_246 = 'b000110000;
    x_247 = 'b000010111;
    x_248 = 'b000011101;
    x_249 = 'b000011100;
    x_250 = 'b000110000;
    x_251 = 'b000101110;
    x_252 = 'b111111100;
    x_253 = 'b000000100;
    x_254 = 'b000010000;
    x_255 = 'b111101000;

    h_0 = 'b000100101;
    h_1 = 'b000100001;
    h_2 = 'b000001010;
    h_3 = 'b000001011;
    h_4 = 'b000000001;
    h_5 = 'b111111101;
    h_6 = 'b111111101;
    h_7 = 'b000101010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000111001;
    x_1 = 'b000110110;
    x_2 = 'b000011111;
    x_3 = 'b000011100;
    x_4 = 'b000010111;
    x_5 = 'b000010110;
    x_6 = 'b000010000;
    x_7 = 'b000111011;
    x_8 = 'b000101010;
    x_9 = 'b000100101;
    x_10 = 'b000100001;
    x_11 = 'b000011101;
    x_12 = 'b000100110;
    x_13 = 'b000100000;
    x_14 = 'b000110001;
    x_15 = 'b000101111;
    x_16 = 'b000100101;
    x_17 = 'b000100111;
    x_18 = 'b000101010;
    x_19 = 'b000110011;
    x_20 = 'b000111001;
    x_21 = 'b000011000;
    x_22 = 'b000011001;
    x_23 = 'b000010110;
    x_24 = 'b000100011;
    x_25 = 'b000100011;
    x_26 = 'b000010000;
    x_27 = 'b000001011;
    x_28 = 'b000010100;
    x_29 = 'b000011111;
    x_30 = 'b000111000;
    x_31 = 'b000011001;
    x_32 = 'b000011010;
    x_33 = 'b000010100;
    x_34 = 'b000001111;
    x_35 = 'b000001011;
    x_36 = 'b000001011;
    x_37 = 'b111010110;
    x_38 = 'b000101101;
    x_39 = 'b000010011;
    x_40 = 'b000101101;
    x_41 = 'b000001110;
    x_42 = 'b000101001;
    x_43 = 'b111111110;
    x_44 = 'b000101100;
    x_45 = 'b001000011;
    x_46 = 'b000100110;
    x_47 = 'b000100100;
    x_48 = 'b000100011;
    x_49 = 'b000100011;
    x_50 = 'b000100110;
    x_51 = 'b000111000;
    x_52 = 'b000111101;
    x_53 = 'b000111110;
    x_54 = 'b001000000;
    x_55 = 'b000011001;
    x_56 = 'b000011100;
    x_57 = 'b000100111;
    x_58 = 'b001000100;
    x_59 = 'b000111010;
    x_60 = 'b000000100;
    x_61 = 'b000010101;
    x_62 = 'b000100001;
    x_63 = 'b111110100;
    x_64 = 'b000111001;
    x_65 = 'b000110110;
    x_66 = 'b000011111;
    x_67 = 'b000011100;
    x_68 = 'b000010111;
    x_69 = 'b000010110;
    x_70 = 'b000010000;
    x_71 = 'b000111011;
    x_72 = 'b000101010;
    x_73 = 'b000100101;
    x_74 = 'b000100001;
    x_75 = 'b000011101;
    x_76 = 'b000100110;
    x_77 = 'b000100000;
    x_78 = 'b000110001;
    x_79 = 'b000101111;
    x_80 = 'b000100101;
    x_81 = 'b000100111;
    x_82 = 'b000101010;
    x_83 = 'b000110011;
    x_84 = 'b000111001;
    x_85 = 'b000011000;
    x_86 = 'b000011001;
    x_87 = 'b000010110;
    x_88 = 'b000100011;
    x_89 = 'b000100011;
    x_90 = 'b000010000;
    x_91 = 'b000001011;
    x_92 = 'b000010100;
    x_93 = 'b000011111;
    x_94 = 'b000111000;
    x_95 = 'b000011001;
    x_96 = 'b000011010;
    x_97 = 'b000010100;
    x_98 = 'b000001111;
    x_99 = 'b000001011;
    x_100 = 'b000001011;
    x_101 = 'b111010110;
    x_102 = 'b000101101;
    x_103 = 'b000010011;
    x_104 = 'b000101101;
    x_105 = 'b000001110;
    x_106 = 'b000101001;
    x_107 = 'b111111110;
    x_108 = 'b000101100;
    x_109 = 'b001000011;
    x_110 = 'b000100110;
    x_111 = 'b000100100;
    x_112 = 'b000100011;
    x_113 = 'b000100011;
    x_114 = 'b000100110;
    x_115 = 'b000111000;
    x_116 = 'b000111101;
    x_117 = 'b000111110;
    x_118 = 'b001000000;
    x_119 = 'b000011001;
    x_120 = 'b000011100;
    x_121 = 'b000100111;
    x_122 = 'b001000100;
    x_123 = 'b000111010;
    x_124 = 'b000000100;
    x_125 = 'b000010101;
    x_126 = 'b000100001;
    x_127 = 'b111110100;
    x_128 = 'b000111001;
    x_129 = 'b000110110;
    x_130 = 'b000011111;
    x_131 = 'b000011100;
    x_132 = 'b000010111;
    x_133 = 'b000010110;
    x_134 = 'b000010000;
    x_135 = 'b000111011;
    x_136 = 'b000101010;
    x_137 = 'b000100101;
    x_138 = 'b000100001;
    x_139 = 'b000011101;
    x_140 = 'b000100110;
    x_141 = 'b000100000;
    x_142 = 'b000110001;
    x_143 = 'b000101111;
    x_144 = 'b000100101;
    x_145 = 'b000100111;
    x_146 = 'b000101010;
    x_147 = 'b000110011;
    x_148 = 'b000111001;
    x_149 = 'b000011000;
    x_150 = 'b000011001;
    x_151 = 'b000010110;
    x_152 = 'b000100011;
    x_153 = 'b000100011;
    x_154 = 'b000010000;
    x_155 = 'b000001011;
    x_156 = 'b000010100;
    x_157 = 'b000011111;
    x_158 = 'b000111000;
    x_159 = 'b000011001;
    x_160 = 'b000011010;
    x_161 = 'b000010100;
    x_162 = 'b000001111;
    x_163 = 'b000001011;
    x_164 = 'b000001011;
    x_165 = 'b111010110;
    x_166 = 'b000101101;
    x_167 = 'b000010011;
    x_168 = 'b000101101;
    x_169 = 'b000001110;
    x_170 = 'b000101001;
    x_171 = 'b111111110;
    x_172 = 'b000101100;
    x_173 = 'b001000011;
    x_174 = 'b000100110;
    x_175 = 'b000100100;
    x_176 = 'b000100011;
    x_177 = 'b000100011;
    x_178 = 'b000100110;
    x_179 = 'b000111000;
    x_180 = 'b000111101;
    x_181 = 'b000111110;
    x_182 = 'b001000000;
    x_183 = 'b000011001;
    x_184 = 'b000011100;
    x_185 = 'b000100111;
    x_186 = 'b001000100;
    x_187 = 'b000111010;
    x_188 = 'b000000100;
    x_189 = 'b000010101;
    x_190 = 'b000100001;
    x_191 = 'b111110100;
    x_192 = 'b000111001;
    x_193 = 'b000110110;
    x_194 = 'b000011111;
    x_195 = 'b000011100;
    x_196 = 'b000010111;
    x_197 = 'b000010110;
    x_198 = 'b000010000;
    x_199 = 'b000111011;
    x_200 = 'b000101010;
    x_201 = 'b000100101;
    x_202 = 'b000100001;
    x_203 = 'b000011101;
    x_204 = 'b000100110;
    x_205 = 'b000100000;
    x_206 = 'b000110001;
    x_207 = 'b000101111;
    x_208 = 'b000100101;
    x_209 = 'b000100111;
    x_210 = 'b000101010;
    x_211 = 'b000110011;
    x_212 = 'b000111001;
    x_213 = 'b000011000;
    x_214 = 'b000011001;
    x_215 = 'b000010110;
    x_216 = 'b000100011;
    x_217 = 'b000100011;
    x_218 = 'b000010000;
    x_219 = 'b000001011;
    x_220 = 'b000010100;
    x_221 = 'b000011111;
    x_222 = 'b000111000;
    x_223 = 'b000011001;
    x_224 = 'b000011010;
    x_225 = 'b000010100;
    x_226 = 'b000001111;
    x_227 = 'b000001011;
    x_228 = 'b000001011;
    x_229 = 'b111010110;
    x_230 = 'b000101101;
    x_231 = 'b000010011;
    x_232 = 'b000101101;
    x_233 = 'b000001110;
    x_234 = 'b000101001;
    x_235 = 'b111111110;
    x_236 = 'b000101100;
    x_237 = 'b001000011;
    x_238 = 'b000100110;
    x_239 = 'b000100100;
    x_240 = 'b000100011;
    x_241 = 'b000100011;
    x_242 = 'b000100110;
    x_243 = 'b000111000;
    x_244 = 'b000111101;
    x_245 = 'b000111110;
    x_246 = 'b001000000;
    x_247 = 'b000011001;
    x_248 = 'b000011100;
    x_249 = 'b000100111;
    x_250 = 'b001000100;
    x_251 = 'b000111010;
    x_252 = 'b000000100;
    x_253 = 'b000010101;
    x_254 = 'b000100001;
    x_255 = 'b111110100;

    h_0 = 'b000111001;
    h_1 = 'b000110110;
    h_2 = 'b000011111;
    h_3 = 'b000011100;
    h_4 = 'b000010111;
    h_5 = 'b000010110;
    h_6 = 'b000010000;
    h_7 = 'b000111011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000010111;
    x_1 = 'b000011001;
    x_2 = 'b000001000;
    x_3 = 'b000001001;
    x_4 = 'b000001101;
    x_5 = 'b000010000;
    x_6 = 'b000010101;
    x_7 = 'b000011010;
    x_8 = 'b000010000;
    x_9 = 'b000001110;
    x_10 = 'b000001110;
    x_11 = 'b000010000;
    x_12 = 'b000100100;
    x_13 = 'b000100110;
    x_14 = 'b000011000;
    x_15 = 'b000010111;
    x_16 = 'b000010010;
    x_17 = 'b000010111;
    x_18 = 'b000011101;
    x_19 = 'b000101011;
    x_20 = 'b000110110;
    x_21 = 'b111110111;
    x_22 = 'b000000001;
    x_23 = 'b000001011;
    x_24 = 'b111111010;
    x_25 = 'b111111010;
    x_26 = 'b111111001;
    x_27 = 'b000000001;
    x_28 = 'b000001101;
    x_29 = 'b111110110;
    x_30 = 'b000001001;
    x_31 = 'b000000111;
    x_32 = 'b111111011;
    x_33 = 'b111111011;
    x_34 = 'b111111110;
    x_35 = 'b111110111;
    x_36 = 'b000001011;
    x_37 = 'b111011100;
    x_38 = 'b111111101;
    x_39 = 'b000011000;
    x_40 = 'b000010011;
    x_41 = 'b000010111;
    x_42 = 'b000000100;
    x_43 = 'b000100111;
    x_44 = 'b000010001;
    x_45 = 'b000110001;
    x_46 = 'b000010010;
    x_47 = 'b000010010;
    x_48 = 'b000010001;
    x_49 = 'b000010011;
    x_50 = 'b000011011;
    x_51 = 'b000101101;
    x_52 = 'b000110000;
    x_53 = 'b000110001;
    x_54 = 'b000101010;
    x_55 = 'b000001111;
    x_56 = 'b000010011;
    x_57 = 'b000100001;
    x_58 = 'b000111001;
    x_59 = 'b000101110;
    x_60 = 'b000000111;
    x_61 = 'b000100010;
    x_62 = 'b000101101;
    x_63 = 'b000000011;
    x_64 = 'b000010111;
    x_65 = 'b000011001;
    x_66 = 'b000001000;
    x_67 = 'b000001001;
    x_68 = 'b000001101;
    x_69 = 'b000010000;
    x_70 = 'b000010101;
    x_71 = 'b000011010;
    x_72 = 'b000010000;
    x_73 = 'b000001110;
    x_74 = 'b000001110;
    x_75 = 'b000010000;
    x_76 = 'b000100100;
    x_77 = 'b000100110;
    x_78 = 'b000011000;
    x_79 = 'b000010111;
    x_80 = 'b000010010;
    x_81 = 'b000010111;
    x_82 = 'b000011101;
    x_83 = 'b000101011;
    x_84 = 'b000110110;
    x_85 = 'b111110111;
    x_86 = 'b000000001;
    x_87 = 'b000001011;
    x_88 = 'b111111010;
    x_89 = 'b111111010;
    x_90 = 'b111111001;
    x_91 = 'b000000001;
    x_92 = 'b000001101;
    x_93 = 'b111110110;
    x_94 = 'b000001001;
    x_95 = 'b000000111;
    x_96 = 'b111111011;
    x_97 = 'b111111011;
    x_98 = 'b111111110;
    x_99 = 'b111110111;
    x_100 = 'b000001011;
    x_101 = 'b111011100;
    x_102 = 'b111111101;
    x_103 = 'b000011000;
    x_104 = 'b000010011;
    x_105 = 'b000010111;
    x_106 = 'b000000100;
    x_107 = 'b000100111;
    x_108 = 'b000010001;
    x_109 = 'b000110001;
    x_110 = 'b000010010;
    x_111 = 'b000010010;
    x_112 = 'b000010001;
    x_113 = 'b000010011;
    x_114 = 'b000011011;
    x_115 = 'b000101101;
    x_116 = 'b000110000;
    x_117 = 'b000110001;
    x_118 = 'b000101010;
    x_119 = 'b000001111;
    x_120 = 'b000010011;
    x_121 = 'b000100001;
    x_122 = 'b000111001;
    x_123 = 'b000101110;
    x_124 = 'b000000111;
    x_125 = 'b000100010;
    x_126 = 'b000101101;
    x_127 = 'b000000011;
    x_128 = 'b000010111;
    x_129 = 'b000011001;
    x_130 = 'b000001000;
    x_131 = 'b000001001;
    x_132 = 'b000001101;
    x_133 = 'b000010000;
    x_134 = 'b000010101;
    x_135 = 'b000011010;
    x_136 = 'b000010000;
    x_137 = 'b000001110;
    x_138 = 'b000001110;
    x_139 = 'b000010000;
    x_140 = 'b000100100;
    x_141 = 'b000100110;
    x_142 = 'b000011000;
    x_143 = 'b000010111;
    x_144 = 'b000010010;
    x_145 = 'b000010111;
    x_146 = 'b000011101;
    x_147 = 'b000101011;
    x_148 = 'b000110110;
    x_149 = 'b111110111;
    x_150 = 'b000000001;
    x_151 = 'b000001011;
    x_152 = 'b111111010;
    x_153 = 'b111111010;
    x_154 = 'b111111001;
    x_155 = 'b000000001;
    x_156 = 'b000001101;
    x_157 = 'b111110110;
    x_158 = 'b000001001;
    x_159 = 'b000000111;
    x_160 = 'b111111011;
    x_161 = 'b111111011;
    x_162 = 'b111111110;
    x_163 = 'b111110111;
    x_164 = 'b000001011;
    x_165 = 'b111011100;
    x_166 = 'b111111101;
    x_167 = 'b000011000;
    x_168 = 'b000010011;
    x_169 = 'b000010111;
    x_170 = 'b000000100;
    x_171 = 'b000100111;
    x_172 = 'b000010001;
    x_173 = 'b000110001;
    x_174 = 'b000010010;
    x_175 = 'b000010010;
    x_176 = 'b000010001;
    x_177 = 'b000010011;
    x_178 = 'b000011011;
    x_179 = 'b000101101;
    x_180 = 'b000110000;
    x_181 = 'b000110001;
    x_182 = 'b000101010;
    x_183 = 'b000001111;
    x_184 = 'b000010011;
    x_185 = 'b000100001;
    x_186 = 'b000111001;
    x_187 = 'b000101110;
    x_188 = 'b000000111;
    x_189 = 'b000100010;
    x_190 = 'b000101101;
    x_191 = 'b000000011;
    x_192 = 'b000010111;
    x_193 = 'b000011001;
    x_194 = 'b000001000;
    x_195 = 'b000001001;
    x_196 = 'b000001101;
    x_197 = 'b000010000;
    x_198 = 'b000010101;
    x_199 = 'b000011010;
    x_200 = 'b000010000;
    x_201 = 'b000001110;
    x_202 = 'b000001110;
    x_203 = 'b000010000;
    x_204 = 'b000100100;
    x_205 = 'b000100110;
    x_206 = 'b000011000;
    x_207 = 'b000010111;
    x_208 = 'b000010010;
    x_209 = 'b000010111;
    x_210 = 'b000011101;
    x_211 = 'b000101011;
    x_212 = 'b000110110;
    x_213 = 'b111110111;
    x_214 = 'b000000001;
    x_215 = 'b000001011;
    x_216 = 'b111111010;
    x_217 = 'b111111010;
    x_218 = 'b111111001;
    x_219 = 'b000000001;
    x_220 = 'b000001101;
    x_221 = 'b111110110;
    x_222 = 'b000001001;
    x_223 = 'b000000111;
    x_224 = 'b111111011;
    x_225 = 'b111111011;
    x_226 = 'b111111110;
    x_227 = 'b111110111;
    x_228 = 'b000001011;
    x_229 = 'b111011100;
    x_230 = 'b111111101;
    x_231 = 'b000011000;
    x_232 = 'b000010011;
    x_233 = 'b000010111;
    x_234 = 'b000000100;
    x_235 = 'b000100111;
    x_236 = 'b000010001;
    x_237 = 'b000110001;
    x_238 = 'b000010010;
    x_239 = 'b000010010;
    x_240 = 'b000010001;
    x_241 = 'b000010011;
    x_242 = 'b000011011;
    x_243 = 'b000101101;
    x_244 = 'b000110000;
    x_245 = 'b000110001;
    x_246 = 'b000101010;
    x_247 = 'b000001111;
    x_248 = 'b000010011;
    x_249 = 'b000100001;
    x_250 = 'b000111001;
    x_251 = 'b000101110;
    x_252 = 'b000000111;
    x_253 = 'b000100010;
    x_254 = 'b000101101;
    x_255 = 'b000000011;

    h_0 = 'b000010111;
    h_1 = 'b000011001;
    h_2 = 'b000001000;
    h_3 = 'b000001001;
    h_4 = 'b000001101;
    h_5 = 'b000010000;
    h_6 = 'b000010101;
    h_7 = 'b000011010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000000110;
    x_1 = 'b000001011;
    x_2 = 'b111111101;
    x_3 = 'b000000010;
    x_4 = 'b000001001;
    x_5 = 'b000001110;
    x_6 = 'b000010101;
    x_7 = 'b000010110;
    x_8 = 'b000000111;
    x_9 = 'b000001000;
    x_10 = 'b000001011;
    x_11 = 'b000010000;
    x_12 = 'b000011111;
    x_13 = 'b000100111;
    x_14 = 'b000010110;
    x_15 = 'b000010011;
    x_16 = 'b000001110;
    x_17 = 'b000010101;
    x_18 = 'b000011001;
    x_19 = 'b000100100;
    x_20 = 'b000110001;
    x_21 = 'b000000011;
    x_22 = 'b000001010;
    x_23 = 'b000001110;
    x_24 = 'b000001101;
    x_25 = 'b000001011;
    x_26 = 'b111111110;
    x_27 = 'b000000100;
    x_28 = 'b000010001;
    x_29 = 'b000010000;
    x_30 = 'b000011111;
    x_31 = 'b000001110;
    x_32 = 'b000000101;
    x_33 = 'b000000100;
    x_34 = 'b000000011;
    x_35 = 'b000000000;
    x_36 = 'b000001101;
    x_37 = 'b111010100;
    x_38 = 'b000100001;
    x_39 = 'b000010000;
    x_40 = 'b000011100;
    x_41 = 'b000010000;
    x_42 = 'b000101111;
    x_43 = 'b111111110;
    x_44 = 'b000011110;
    x_45 = 'b000100011;
    x_46 = 'b000100100;
    x_47 = 'b000100100;
    x_48 = 'b000011111;
    x_49 = 'b000011111;
    x_50 = 'b000100010;
    x_51 = 'b000101111;
    x_52 = 'b000110000;
    x_53 = 'b000101101;
    x_54 = 'b000100111;
    x_55 = 'b000100101;
    x_56 = 'b000100111;
    x_57 = 'b000101011;
    x_58 = 'b000111010;
    x_59 = 'b000101110;
    x_60 = 'b000010001;
    x_61 = 'b000101100;
    x_62 = 'b000110010;
    x_63 = 'b000011010;
    x_64 = 'b000000110;
    x_65 = 'b000001011;
    x_66 = 'b111111101;
    x_67 = 'b000000010;
    x_68 = 'b000001001;
    x_69 = 'b000001110;
    x_70 = 'b000010101;
    x_71 = 'b000010110;
    x_72 = 'b000000111;
    x_73 = 'b000001000;
    x_74 = 'b000001011;
    x_75 = 'b000010000;
    x_76 = 'b000011111;
    x_77 = 'b000100111;
    x_78 = 'b000010110;
    x_79 = 'b000010011;
    x_80 = 'b000001110;
    x_81 = 'b000010101;
    x_82 = 'b000011001;
    x_83 = 'b000100100;
    x_84 = 'b000110001;
    x_85 = 'b000000011;
    x_86 = 'b000001010;
    x_87 = 'b000001110;
    x_88 = 'b000001101;
    x_89 = 'b000001011;
    x_90 = 'b111111110;
    x_91 = 'b000000100;
    x_92 = 'b000010001;
    x_93 = 'b000010000;
    x_94 = 'b000011111;
    x_95 = 'b000001110;
    x_96 = 'b000000101;
    x_97 = 'b000000100;
    x_98 = 'b000000011;
    x_99 = 'b000000000;
    x_100 = 'b000001101;
    x_101 = 'b111010100;
    x_102 = 'b000100001;
    x_103 = 'b000010000;
    x_104 = 'b000011100;
    x_105 = 'b000010000;
    x_106 = 'b000101111;
    x_107 = 'b111111110;
    x_108 = 'b000011110;
    x_109 = 'b000100011;
    x_110 = 'b000100100;
    x_111 = 'b000100100;
    x_112 = 'b000011111;
    x_113 = 'b000011111;
    x_114 = 'b000100010;
    x_115 = 'b000101111;
    x_116 = 'b000110000;
    x_117 = 'b000101101;
    x_118 = 'b000100111;
    x_119 = 'b000100101;
    x_120 = 'b000100111;
    x_121 = 'b000101011;
    x_122 = 'b000111010;
    x_123 = 'b000101110;
    x_124 = 'b000010001;
    x_125 = 'b000101100;
    x_126 = 'b000110010;
    x_127 = 'b000011010;
    x_128 = 'b000000110;
    x_129 = 'b000001011;
    x_130 = 'b111111101;
    x_131 = 'b000000010;
    x_132 = 'b000001001;
    x_133 = 'b000001110;
    x_134 = 'b000010101;
    x_135 = 'b000010110;
    x_136 = 'b000000111;
    x_137 = 'b000001000;
    x_138 = 'b000001011;
    x_139 = 'b000010000;
    x_140 = 'b000011111;
    x_141 = 'b000100111;
    x_142 = 'b000010110;
    x_143 = 'b000010011;
    x_144 = 'b000001110;
    x_145 = 'b000010101;
    x_146 = 'b000011001;
    x_147 = 'b000100100;
    x_148 = 'b000110001;
    x_149 = 'b000000011;
    x_150 = 'b000001010;
    x_151 = 'b000001110;
    x_152 = 'b000001101;
    x_153 = 'b000001011;
    x_154 = 'b111111110;
    x_155 = 'b000000100;
    x_156 = 'b000010001;
    x_157 = 'b000010000;
    x_158 = 'b000011111;
    x_159 = 'b000001110;
    x_160 = 'b000000101;
    x_161 = 'b000000100;
    x_162 = 'b000000011;
    x_163 = 'b000000000;
    x_164 = 'b000001101;
    x_165 = 'b111010100;
    x_166 = 'b000100001;
    x_167 = 'b000010000;
    x_168 = 'b000011100;
    x_169 = 'b000010000;
    x_170 = 'b000101111;
    x_171 = 'b111111110;
    x_172 = 'b000011110;
    x_173 = 'b000100011;
    x_174 = 'b000100100;
    x_175 = 'b000100100;
    x_176 = 'b000011111;
    x_177 = 'b000011111;
    x_178 = 'b000100010;
    x_179 = 'b000101111;
    x_180 = 'b000110000;
    x_181 = 'b000101101;
    x_182 = 'b000100111;
    x_183 = 'b000100101;
    x_184 = 'b000100111;
    x_185 = 'b000101011;
    x_186 = 'b000111010;
    x_187 = 'b000101110;
    x_188 = 'b000010001;
    x_189 = 'b000101100;
    x_190 = 'b000110010;
    x_191 = 'b000011010;
    x_192 = 'b000000110;
    x_193 = 'b000001011;
    x_194 = 'b111111101;
    x_195 = 'b000000010;
    x_196 = 'b000001001;
    x_197 = 'b000001110;
    x_198 = 'b000010101;
    x_199 = 'b000010110;
    x_200 = 'b000000111;
    x_201 = 'b000001000;
    x_202 = 'b000001011;
    x_203 = 'b000010000;
    x_204 = 'b000011111;
    x_205 = 'b000100111;
    x_206 = 'b000010110;
    x_207 = 'b000010011;
    x_208 = 'b000001110;
    x_209 = 'b000010101;
    x_210 = 'b000011001;
    x_211 = 'b000100100;
    x_212 = 'b000110001;
    x_213 = 'b000000011;
    x_214 = 'b000001010;
    x_215 = 'b000001110;
    x_216 = 'b000001101;
    x_217 = 'b000001011;
    x_218 = 'b111111110;
    x_219 = 'b000000100;
    x_220 = 'b000010001;
    x_221 = 'b000010000;
    x_222 = 'b000011111;
    x_223 = 'b000001110;
    x_224 = 'b000000101;
    x_225 = 'b000000100;
    x_226 = 'b000000011;
    x_227 = 'b000000000;
    x_228 = 'b000001101;
    x_229 = 'b111010100;
    x_230 = 'b000100001;
    x_231 = 'b000010000;
    x_232 = 'b000011100;
    x_233 = 'b000010000;
    x_234 = 'b000101111;
    x_235 = 'b111111110;
    x_236 = 'b000011110;
    x_237 = 'b000100011;
    x_238 = 'b000100100;
    x_239 = 'b000100100;
    x_240 = 'b000011111;
    x_241 = 'b000011111;
    x_242 = 'b000100010;
    x_243 = 'b000101111;
    x_244 = 'b000110000;
    x_245 = 'b000101101;
    x_246 = 'b000100111;
    x_247 = 'b000100101;
    x_248 = 'b000100111;
    x_249 = 'b000101011;
    x_250 = 'b000111010;
    x_251 = 'b000101110;
    x_252 = 'b000010001;
    x_253 = 'b000101100;
    x_254 = 'b000110010;
    x_255 = 'b000011010;

    h_0 = 'b000000110;
    h_1 = 'b000001011;
    h_2 = 'b111111101;
    h_3 = 'b000000010;
    h_4 = 'b000001001;
    h_5 = 'b000001110;
    h_6 = 'b000010101;
    h_7 = 'b000010110;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000100110;
    x_1 = 'b000100001;
    x_2 = 'b000001011;
    x_3 = 'b000010001;
    x_4 = 'b000001101;
    x_5 = 'b000001110;
    x_6 = 'b000010100;
    x_7 = 'b000110110;
    x_8 = 'b000011101;
    x_9 = 'b000010110;
    x_10 = 'b000010101;
    x_11 = 'b000010011;
    x_12 = 'b000011001;
    x_13 = 'b000011100;
    x_14 = 'b000110001;
    x_15 = 'b000100100;
    x_16 = 'b000011100;
    x_17 = 'b000011101;
    x_18 = 'b000011011;
    x_19 = 'b000100010;
    x_20 = 'b000101001;
    x_21 = 'b000001110;
    x_22 = 'b000010101;
    x_23 = 'b000010111;
    x_24 = 'b000010111;
    x_25 = 'b000010111;
    x_26 = 'b000000011;
    x_27 = 'b000001010;
    x_28 = 'b000011110;
    x_29 = 'b000011010;
    x_30 = 'b000100111;
    x_31 = 'b000001100;
    x_32 = 'b000001001;
    x_33 = 'b000000110;
    x_34 = 'b000000011;
    x_35 = 'b111111111;
    x_36 = 'b000001100;
    x_37 = 'b111011111;
    x_38 = 'b000100001;
    x_39 = 'b000010010;
    x_40 = 'b000100111;
    x_41 = 'b000000110;
    x_42 = 'b000101110;
    x_43 = 'b000001100;
    x_44 = 'b000110110;
    x_45 = 'b000011010;
    x_46 = 'b000110100;
    x_47 = 'b000101011;
    x_48 = 'b000100010;
    x_49 = 'b000011111;
    x_50 = 'b000011111;
    x_51 = 'b000101001;
    x_52 = 'b000100111;
    x_53 = 'b000100101;
    x_54 = 'b000100101;
    x_55 = 'b000100111;
    x_56 = 'b000100101;
    x_57 = 'b000100101;
    x_58 = 'b000110100;
    x_59 = 'b000101100;
    x_60 = 'b000011011;
    x_61 = 'b000110011;
    x_62 = 'b000110010;
    x_63 = 'b000101010;
    x_64 = 'b000100110;
    x_65 = 'b000100001;
    x_66 = 'b000001011;
    x_67 = 'b000010001;
    x_68 = 'b000001101;
    x_69 = 'b000001110;
    x_70 = 'b000010100;
    x_71 = 'b000110110;
    x_72 = 'b000011101;
    x_73 = 'b000010110;
    x_74 = 'b000010101;
    x_75 = 'b000010011;
    x_76 = 'b000011001;
    x_77 = 'b000011100;
    x_78 = 'b000110001;
    x_79 = 'b000100100;
    x_80 = 'b000011100;
    x_81 = 'b000011101;
    x_82 = 'b000011011;
    x_83 = 'b000100010;
    x_84 = 'b000101001;
    x_85 = 'b000001110;
    x_86 = 'b000010101;
    x_87 = 'b000010111;
    x_88 = 'b000010111;
    x_89 = 'b000010111;
    x_90 = 'b000000011;
    x_91 = 'b000001010;
    x_92 = 'b000011110;
    x_93 = 'b000011010;
    x_94 = 'b000100111;
    x_95 = 'b000001100;
    x_96 = 'b000001001;
    x_97 = 'b000000110;
    x_98 = 'b000000011;
    x_99 = 'b111111111;
    x_100 = 'b000001100;
    x_101 = 'b111011111;
    x_102 = 'b000100001;
    x_103 = 'b000010010;
    x_104 = 'b000100111;
    x_105 = 'b000000110;
    x_106 = 'b000101110;
    x_107 = 'b000001100;
    x_108 = 'b000110110;
    x_109 = 'b000011010;
    x_110 = 'b000110100;
    x_111 = 'b000101011;
    x_112 = 'b000100010;
    x_113 = 'b000011111;
    x_114 = 'b000011111;
    x_115 = 'b000101001;
    x_116 = 'b000100111;
    x_117 = 'b000100101;
    x_118 = 'b000100101;
    x_119 = 'b000100111;
    x_120 = 'b000100101;
    x_121 = 'b000100101;
    x_122 = 'b000110100;
    x_123 = 'b000101100;
    x_124 = 'b000011011;
    x_125 = 'b000110011;
    x_126 = 'b000110010;
    x_127 = 'b000101010;
    x_128 = 'b000100110;
    x_129 = 'b000100001;
    x_130 = 'b000001011;
    x_131 = 'b000010001;
    x_132 = 'b000001101;
    x_133 = 'b000001110;
    x_134 = 'b000010100;
    x_135 = 'b000110110;
    x_136 = 'b000011101;
    x_137 = 'b000010110;
    x_138 = 'b000010101;
    x_139 = 'b000010011;
    x_140 = 'b000011001;
    x_141 = 'b000011100;
    x_142 = 'b000110001;
    x_143 = 'b000100100;
    x_144 = 'b000011100;
    x_145 = 'b000011101;
    x_146 = 'b000011011;
    x_147 = 'b000100010;
    x_148 = 'b000101001;
    x_149 = 'b000001110;
    x_150 = 'b000010101;
    x_151 = 'b000010111;
    x_152 = 'b000010111;
    x_153 = 'b000010111;
    x_154 = 'b000000011;
    x_155 = 'b000001010;
    x_156 = 'b000011110;
    x_157 = 'b000011010;
    x_158 = 'b000100111;
    x_159 = 'b000001100;
    x_160 = 'b000001001;
    x_161 = 'b000000110;
    x_162 = 'b000000011;
    x_163 = 'b111111111;
    x_164 = 'b000001100;
    x_165 = 'b111011111;
    x_166 = 'b000100001;
    x_167 = 'b000010010;
    x_168 = 'b000100111;
    x_169 = 'b000000110;
    x_170 = 'b000101110;
    x_171 = 'b000001100;
    x_172 = 'b000110110;
    x_173 = 'b000011010;
    x_174 = 'b000110100;
    x_175 = 'b000101011;
    x_176 = 'b000100010;
    x_177 = 'b000011111;
    x_178 = 'b000011111;
    x_179 = 'b000101001;
    x_180 = 'b000100111;
    x_181 = 'b000100101;
    x_182 = 'b000100101;
    x_183 = 'b000100111;
    x_184 = 'b000100101;
    x_185 = 'b000100101;
    x_186 = 'b000110100;
    x_187 = 'b000101100;
    x_188 = 'b000011011;
    x_189 = 'b000110011;
    x_190 = 'b000110010;
    x_191 = 'b000101010;
    x_192 = 'b000100110;
    x_193 = 'b000100001;
    x_194 = 'b000001011;
    x_195 = 'b000010001;
    x_196 = 'b000001101;
    x_197 = 'b000001110;
    x_198 = 'b000010100;
    x_199 = 'b000110110;
    x_200 = 'b000011101;
    x_201 = 'b000010110;
    x_202 = 'b000010101;
    x_203 = 'b000010011;
    x_204 = 'b000011001;
    x_205 = 'b000011100;
    x_206 = 'b000110001;
    x_207 = 'b000100100;
    x_208 = 'b000011100;
    x_209 = 'b000011101;
    x_210 = 'b000011011;
    x_211 = 'b000100010;
    x_212 = 'b000101001;
    x_213 = 'b000001110;
    x_214 = 'b000010101;
    x_215 = 'b000010111;
    x_216 = 'b000010111;
    x_217 = 'b000010111;
    x_218 = 'b000000011;
    x_219 = 'b000001010;
    x_220 = 'b000011110;
    x_221 = 'b000011010;
    x_222 = 'b000100111;
    x_223 = 'b000001100;
    x_224 = 'b000001001;
    x_225 = 'b000000110;
    x_226 = 'b000000011;
    x_227 = 'b111111111;
    x_228 = 'b000001100;
    x_229 = 'b111011111;
    x_230 = 'b000100001;
    x_231 = 'b000010010;
    x_232 = 'b000100111;
    x_233 = 'b000000110;
    x_234 = 'b000101110;
    x_235 = 'b000001100;
    x_236 = 'b000110110;
    x_237 = 'b000011010;
    x_238 = 'b000110100;
    x_239 = 'b000101011;
    x_240 = 'b000100010;
    x_241 = 'b000011111;
    x_242 = 'b000011111;
    x_243 = 'b000101001;
    x_244 = 'b000100111;
    x_245 = 'b000100101;
    x_246 = 'b000100101;
    x_247 = 'b000100111;
    x_248 = 'b000100101;
    x_249 = 'b000100101;
    x_250 = 'b000110100;
    x_251 = 'b000101100;
    x_252 = 'b000011011;
    x_253 = 'b000110011;
    x_254 = 'b000110010;
    x_255 = 'b000101010;

    h_0 = 'b000100110;
    h_1 = 'b000100001;
    h_2 = 'b000001011;
    h_3 = 'b000010001;
    h_4 = 'b000001101;
    h_5 = 'b000001110;
    h_6 = 'b000010100;
    h_7 = 'b000110110;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000001001;
    x_1 = 'b000001110;
    x_2 = 'b111111111;
    x_3 = 'b000000111;
    x_4 = 'b111111111;
    x_5 = 'b111111100;
    x_6 = 'b000000011;
    x_7 = 'b000011010;
    x_8 = 'b000001011;
    x_9 = 'b000001100;
    x_10 = 'b000001100;
    x_11 = 'b000000001;
    x_12 = 'b000001000;
    x_13 = 'b000000011;
    x_14 = 'b000100100;
    x_15 = 'b000011000;
    x_16 = 'b000010010;
    x_17 = 'b000010101;
    x_18 = 'b000001111;
    x_19 = 'b000010101;
    x_20 = 'b000011000;
    x_21 = 'b111110101;
    x_22 = 'b111111110;
    x_23 = 'b000000101;
    x_24 = 'b111111010;
    x_25 = 'b111111010;
    x_26 = 'b111101111;
    x_27 = 'b111110101;
    x_28 = 'b000001010;
    x_29 = 'b111111000;
    x_30 = 'b000001101;
    x_31 = 'b111111100;
    x_32 = 'b111111010;
    x_33 = 'b111110110;
    x_34 = 'b111110010;
    x_35 = 'b111101011;
    x_36 = 'b111110100;
    x_37 = 'b111010101;
    x_38 = 'b111111111;
    x_39 = 'b111111011;
    x_40 = 'b000101010;
    x_41 = 'b111011101;
    x_42 = 'b000101001;
    x_43 = 'b000010001;
    x_44 = 'b000110110;
    x_45 = 'b000100100;
    x_46 = 'b000110001;
    x_47 = 'b000100111;
    x_48 = 'b000100001;
    x_49 = 'b000011110;
    x_50 = 'b000011100;
    x_51 = 'b000101000;
    x_52 = 'b000100111;
    x_53 = 'b000100110;
    x_54 = 'b000101101;
    x_55 = 'b000011111;
    x_56 = 'b000100001;
    x_57 = 'b000100011;
    x_58 = 'b000110110;
    x_59 = 'b000110011;
    x_60 = 'b000011011;
    x_61 = 'b000110011;
    x_62 = 'b000110000;
    x_63 = 'b000101001;
    x_64 = 'b000001001;
    x_65 = 'b000001110;
    x_66 = 'b111111111;
    x_67 = 'b000000111;
    x_68 = 'b111111111;
    x_69 = 'b111111100;
    x_70 = 'b000000011;
    x_71 = 'b000011010;
    x_72 = 'b000001011;
    x_73 = 'b000001100;
    x_74 = 'b000001100;
    x_75 = 'b000000001;
    x_76 = 'b000001000;
    x_77 = 'b000000011;
    x_78 = 'b000100100;
    x_79 = 'b000011000;
    x_80 = 'b000010010;
    x_81 = 'b000010101;
    x_82 = 'b000001111;
    x_83 = 'b000010101;
    x_84 = 'b000011000;
    x_85 = 'b111110101;
    x_86 = 'b111111110;
    x_87 = 'b000000101;
    x_88 = 'b111111010;
    x_89 = 'b111111010;
    x_90 = 'b111101111;
    x_91 = 'b111110101;
    x_92 = 'b000001010;
    x_93 = 'b111111000;
    x_94 = 'b000001101;
    x_95 = 'b111111100;
    x_96 = 'b111111010;
    x_97 = 'b111110110;
    x_98 = 'b111110010;
    x_99 = 'b111101011;
    x_100 = 'b111110100;
    x_101 = 'b111010101;
    x_102 = 'b111111111;
    x_103 = 'b111111011;
    x_104 = 'b000101010;
    x_105 = 'b111011101;
    x_106 = 'b000101001;
    x_107 = 'b000010001;
    x_108 = 'b000110110;
    x_109 = 'b000100100;
    x_110 = 'b000110001;
    x_111 = 'b000100111;
    x_112 = 'b000100001;
    x_113 = 'b000011110;
    x_114 = 'b000011100;
    x_115 = 'b000101000;
    x_116 = 'b000100111;
    x_117 = 'b000100110;
    x_118 = 'b000101101;
    x_119 = 'b000011111;
    x_120 = 'b000100001;
    x_121 = 'b000100011;
    x_122 = 'b000110110;
    x_123 = 'b000110011;
    x_124 = 'b000011011;
    x_125 = 'b000110011;
    x_126 = 'b000110000;
    x_127 = 'b000101001;
    x_128 = 'b000001001;
    x_129 = 'b000001110;
    x_130 = 'b111111111;
    x_131 = 'b000000111;
    x_132 = 'b111111111;
    x_133 = 'b111111100;
    x_134 = 'b000000011;
    x_135 = 'b000011010;
    x_136 = 'b000001011;
    x_137 = 'b000001100;
    x_138 = 'b000001100;
    x_139 = 'b000000001;
    x_140 = 'b000001000;
    x_141 = 'b000000011;
    x_142 = 'b000100100;
    x_143 = 'b000011000;
    x_144 = 'b000010010;
    x_145 = 'b000010101;
    x_146 = 'b000001111;
    x_147 = 'b000010101;
    x_148 = 'b000011000;
    x_149 = 'b111110101;
    x_150 = 'b111111110;
    x_151 = 'b000000101;
    x_152 = 'b111111010;
    x_153 = 'b111111010;
    x_154 = 'b111101111;
    x_155 = 'b111110101;
    x_156 = 'b000001010;
    x_157 = 'b111111000;
    x_158 = 'b000001101;
    x_159 = 'b111111100;
    x_160 = 'b111111010;
    x_161 = 'b111110110;
    x_162 = 'b111110010;
    x_163 = 'b111101011;
    x_164 = 'b111110100;
    x_165 = 'b111010101;
    x_166 = 'b111111111;
    x_167 = 'b111111011;
    x_168 = 'b000101010;
    x_169 = 'b111011101;
    x_170 = 'b000101001;
    x_171 = 'b000010001;
    x_172 = 'b000110110;
    x_173 = 'b000100100;
    x_174 = 'b000110001;
    x_175 = 'b000100111;
    x_176 = 'b000100001;
    x_177 = 'b000011110;
    x_178 = 'b000011100;
    x_179 = 'b000101000;
    x_180 = 'b000100111;
    x_181 = 'b000100110;
    x_182 = 'b000101101;
    x_183 = 'b000011111;
    x_184 = 'b000100001;
    x_185 = 'b000100011;
    x_186 = 'b000110110;
    x_187 = 'b000110011;
    x_188 = 'b000011011;
    x_189 = 'b000110011;
    x_190 = 'b000110000;
    x_191 = 'b000101001;
    x_192 = 'b000001001;
    x_193 = 'b000001110;
    x_194 = 'b111111111;
    x_195 = 'b000000111;
    x_196 = 'b111111111;
    x_197 = 'b111111100;
    x_198 = 'b000000011;
    x_199 = 'b000011010;
    x_200 = 'b000001011;
    x_201 = 'b000001100;
    x_202 = 'b000001100;
    x_203 = 'b000000001;
    x_204 = 'b000001000;
    x_205 = 'b000000011;
    x_206 = 'b000100100;
    x_207 = 'b000011000;
    x_208 = 'b000010010;
    x_209 = 'b000010101;
    x_210 = 'b000001111;
    x_211 = 'b000010101;
    x_212 = 'b000011000;
    x_213 = 'b111110101;
    x_214 = 'b111111110;
    x_215 = 'b000000101;
    x_216 = 'b111111010;
    x_217 = 'b111111010;
    x_218 = 'b111101111;
    x_219 = 'b111110101;
    x_220 = 'b000001010;
    x_221 = 'b111111000;
    x_222 = 'b000001101;
    x_223 = 'b111111100;
    x_224 = 'b111111010;
    x_225 = 'b111110110;
    x_226 = 'b111110010;
    x_227 = 'b111101011;
    x_228 = 'b111110100;
    x_229 = 'b111010101;
    x_230 = 'b111111111;
    x_231 = 'b111111011;
    x_232 = 'b000101010;
    x_233 = 'b111011101;
    x_234 = 'b000101001;
    x_235 = 'b000010001;
    x_236 = 'b000110110;
    x_237 = 'b000100100;
    x_238 = 'b000110001;
    x_239 = 'b000100111;
    x_240 = 'b000100001;
    x_241 = 'b000011110;
    x_242 = 'b000011100;
    x_243 = 'b000101000;
    x_244 = 'b000100111;
    x_245 = 'b000100110;
    x_246 = 'b000101101;
    x_247 = 'b000011111;
    x_248 = 'b000100001;
    x_249 = 'b000100011;
    x_250 = 'b000110110;
    x_251 = 'b000110011;
    x_252 = 'b000011011;
    x_253 = 'b000110011;
    x_254 = 'b000110000;
    x_255 = 'b000101001;

    h_0 = 'b000001001;
    h_1 = 'b000001110;
    h_2 = 'b111111111;
    h_3 = 'b000000111;
    h_4 = 'b111111111;
    h_5 = 'b111111100;
    h_6 = 'b000000011;
    h_7 = 'b000011010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000001001;
    x_1 = 'b000010010;
    x_2 = 'b000000100;
    x_3 = 'b000001010;
    x_4 = 'b000000000;
    x_5 = 'b111111001;
    x_6 = 'b111110101;
    x_7 = 'b000101010;
    x_8 = 'b000010110;
    x_9 = 'b000010110;
    x_10 = 'b000010100;
    x_11 = 'b000001010;
    x_12 = 'b000001011;
    x_13 = 'b111111111;
    x_14 = 'b000110001;
    x_15 = 'b000100111;
    x_16 = 'b000011100;
    x_17 = 'b000011111;
    x_18 = 'b000010110;
    x_19 = 'b000011001;
    x_20 = 'b000011101;
    x_21 = 'b111111110;
    x_22 = 'b000000001;
    x_23 = 'b000000101;
    x_24 = 'b000000111;
    x_25 = 'b000000101;
    x_26 = 'b111110111;
    x_27 = 'b111110110;
    x_28 = 'b000000100;
    x_29 = 'b000000000;
    x_30 = 'b000011000;
    x_31 = 'b000000100;
    x_32 = 'b000001000;
    x_33 = 'b000000100;
    x_34 = 'b111111011;
    x_35 = 'b111110111;
    x_36 = 'b111110111;
    x_37 = 'b111010100;
    x_38 = 'b000001011;
    x_39 = 'b111110111;
    x_40 = 'b000010011;
    x_41 = 'b111100100;
    x_42 = 'b000011110;
    x_43 = 'b000010100;
    x_44 = 'b000100011;
    x_45 = 'b000101001;
    x_46 = 'b000101011;
    x_47 = 'b000101011;
    x_48 = 'b000100111;
    x_49 = 'b000100101;
    x_50 = 'b000100100;
    x_51 = 'b000101010;
    x_52 = 'b000101001;
    x_53 = 'b000100111;
    x_54 = 'b000101010;
    x_55 = 'b000100011;
    x_56 = 'b000100011;
    x_57 = 'b000100011;
    x_58 = 'b000110100;
    x_59 = 'b000101110;
    x_60 = 'b000011001;
    x_61 = 'b000110000;
    x_62 = 'b000101100;
    x_63 = 'b000100011;
    x_64 = 'b000001001;
    x_65 = 'b000010010;
    x_66 = 'b000000100;
    x_67 = 'b000001010;
    x_68 = 'b000000000;
    x_69 = 'b111111001;
    x_70 = 'b111110101;
    x_71 = 'b000101010;
    x_72 = 'b000010110;
    x_73 = 'b000010110;
    x_74 = 'b000010100;
    x_75 = 'b000001010;
    x_76 = 'b000001011;
    x_77 = 'b111111111;
    x_78 = 'b000110001;
    x_79 = 'b000100111;
    x_80 = 'b000011100;
    x_81 = 'b000011111;
    x_82 = 'b000010110;
    x_83 = 'b000011001;
    x_84 = 'b000011101;
    x_85 = 'b111111110;
    x_86 = 'b000000001;
    x_87 = 'b000000101;
    x_88 = 'b000000111;
    x_89 = 'b000000101;
    x_90 = 'b111110111;
    x_91 = 'b111110110;
    x_92 = 'b000000100;
    x_93 = 'b000000000;
    x_94 = 'b000011000;
    x_95 = 'b000000100;
    x_96 = 'b000001000;
    x_97 = 'b000000100;
    x_98 = 'b111111011;
    x_99 = 'b111110111;
    x_100 = 'b111110111;
    x_101 = 'b111010100;
    x_102 = 'b000001011;
    x_103 = 'b111110111;
    x_104 = 'b000010011;
    x_105 = 'b111100100;
    x_106 = 'b000011110;
    x_107 = 'b000010100;
    x_108 = 'b000100011;
    x_109 = 'b000101001;
    x_110 = 'b000101011;
    x_111 = 'b000101011;
    x_112 = 'b000100111;
    x_113 = 'b000100101;
    x_114 = 'b000100100;
    x_115 = 'b000101010;
    x_116 = 'b000101001;
    x_117 = 'b000100111;
    x_118 = 'b000101010;
    x_119 = 'b000100011;
    x_120 = 'b000100011;
    x_121 = 'b000100011;
    x_122 = 'b000110100;
    x_123 = 'b000101110;
    x_124 = 'b000011001;
    x_125 = 'b000110000;
    x_126 = 'b000101100;
    x_127 = 'b000100011;
    x_128 = 'b000001001;
    x_129 = 'b000010010;
    x_130 = 'b000000100;
    x_131 = 'b000001010;
    x_132 = 'b000000000;
    x_133 = 'b111111001;
    x_134 = 'b111110101;
    x_135 = 'b000101010;
    x_136 = 'b000010110;
    x_137 = 'b000010110;
    x_138 = 'b000010100;
    x_139 = 'b000001010;
    x_140 = 'b000001011;
    x_141 = 'b111111111;
    x_142 = 'b000110001;
    x_143 = 'b000100111;
    x_144 = 'b000011100;
    x_145 = 'b000011111;
    x_146 = 'b000010110;
    x_147 = 'b000011001;
    x_148 = 'b000011101;
    x_149 = 'b111111110;
    x_150 = 'b000000001;
    x_151 = 'b000000101;
    x_152 = 'b000000111;
    x_153 = 'b000000101;
    x_154 = 'b111110111;
    x_155 = 'b111110110;
    x_156 = 'b000000100;
    x_157 = 'b000000000;
    x_158 = 'b000011000;
    x_159 = 'b000000100;
    x_160 = 'b000001000;
    x_161 = 'b000000100;
    x_162 = 'b111111011;
    x_163 = 'b111110111;
    x_164 = 'b111110111;
    x_165 = 'b111010100;
    x_166 = 'b000001011;
    x_167 = 'b111110111;
    x_168 = 'b000010011;
    x_169 = 'b111100100;
    x_170 = 'b000011110;
    x_171 = 'b000010100;
    x_172 = 'b000100011;
    x_173 = 'b000101001;
    x_174 = 'b000101011;
    x_175 = 'b000101011;
    x_176 = 'b000100111;
    x_177 = 'b000100101;
    x_178 = 'b000100100;
    x_179 = 'b000101010;
    x_180 = 'b000101001;
    x_181 = 'b000100111;
    x_182 = 'b000101010;
    x_183 = 'b000100011;
    x_184 = 'b000100011;
    x_185 = 'b000100011;
    x_186 = 'b000110100;
    x_187 = 'b000101110;
    x_188 = 'b000011001;
    x_189 = 'b000110000;
    x_190 = 'b000101100;
    x_191 = 'b000100011;
    x_192 = 'b000001001;
    x_193 = 'b000010010;
    x_194 = 'b000000100;
    x_195 = 'b000001010;
    x_196 = 'b000000000;
    x_197 = 'b111111001;
    x_198 = 'b111110101;
    x_199 = 'b000101010;
    x_200 = 'b000010110;
    x_201 = 'b000010110;
    x_202 = 'b000010100;
    x_203 = 'b000001010;
    x_204 = 'b000001011;
    x_205 = 'b111111111;
    x_206 = 'b000110001;
    x_207 = 'b000100111;
    x_208 = 'b000011100;
    x_209 = 'b000011111;
    x_210 = 'b000010110;
    x_211 = 'b000011001;
    x_212 = 'b000011101;
    x_213 = 'b111111110;
    x_214 = 'b000000001;
    x_215 = 'b000000101;
    x_216 = 'b000000111;
    x_217 = 'b000000101;
    x_218 = 'b111110111;
    x_219 = 'b111110110;
    x_220 = 'b000000100;
    x_221 = 'b000000000;
    x_222 = 'b000011000;
    x_223 = 'b000000100;
    x_224 = 'b000001000;
    x_225 = 'b000000100;
    x_226 = 'b111111011;
    x_227 = 'b111110111;
    x_228 = 'b111110111;
    x_229 = 'b111010100;
    x_230 = 'b000001011;
    x_231 = 'b111110111;
    x_232 = 'b000010011;
    x_233 = 'b111100100;
    x_234 = 'b000011110;
    x_235 = 'b000010100;
    x_236 = 'b000100011;
    x_237 = 'b000101001;
    x_238 = 'b000101011;
    x_239 = 'b000101011;
    x_240 = 'b000100111;
    x_241 = 'b000100101;
    x_242 = 'b000100100;
    x_243 = 'b000101010;
    x_244 = 'b000101001;
    x_245 = 'b000100111;
    x_246 = 'b000101010;
    x_247 = 'b000100011;
    x_248 = 'b000100011;
    x_249 = 'b000100011;
    x_250 = 'b000110100;
    x_251 = 'b000101110;
    x_252 = 'b000011001;
    x_253 = 'b000110000;
    x_254 = 'b000101100;
    x_255 = 'b000100011;

    h_0 = 'b000001001;
    h_1 = 'b000010010;
    h_2 = 'b000000100;
    h_3 = 'b000001010;
    h_4 = 'b000000000;
    h_5 = 'b111111001;
    h_6 = 'b111110101;
    h_7 = 'b000101010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000001010;
    x_1 = 'b000011001;
    x_2 = 'b000001110;
    x_3 = 'b000010110;
    x_4 = 'b000001010;
    x_5 = 'b000000110;
    x_6 = 'b000000011;
    x_7 = 'b000100001;
    x_8 = 'b000010111;
    x_9 = 'b000010111;
    x_10 = 'b000010101;
    x_11 = 'b000001111;
    x_12 = 'b000010001;
    x_13 = 'b000000110;
    x_14 = 'b000100000;
    x_15 = 'b000011011;
    x_16 = 'b000010110;
    x_17 = 'b000011100;
    x_18 = 'b000010100;
    x_19 = 'b000010110;
    x_20 = 'b000011010;
    x_21 = 'b111111000;
    x_22 = 'b111111111;
    x_23 = 'b000000100;
    x_24 = 'b111111100;
    x_25 = 'b111111101;
    x_26 = 'b111111100;
    x_27 = 'b111111010;
    x_28 = 'b000000110;
    x_29 = 'b111101011;
    x_30 = 'b000001100;
    x_31 = 'b000000011;
    x_32 = 'b000000110;
    x_33 = 'b000000100;
    x_34 = 'b111111101;
    x_35 = 'b111110101;
    x_36 = 'b111111011;
    x_37 = 'b111010111;
    x_38 = 'b111110101;
    x_39 = 'b000000001;
    x_40 = 'b000000001;
    x_41 = 'b111110110;
    x_42 = 'b000001100;
    x_43 = 'b111101111;
    x_44 = 'b000010010;
    x_45 = 'b000010101;
    x_46 = 'b000010010;
    x_47 = 'b000010010;
    x_48 = 'b000010101;
    x_49 = 'b000010001;
    x_50 = 'b000010101;
    x_51 = 'b000011010;
    x_52 = 'b000011001;
    x_53 = 'b000010111;
    x_54 = 'b000011001;
    x_55 = 'b000010000;
    x_56 = 'b000010010;
    x_57 = 'b000010010;
    x_58 = 'b000100100;
    x_59 = 'b000011111;
    x_60 = 'b000001111;
    x_61 = 'b000100011;
    x_62 = 'b000011101;
    x_63 = 'b000010000;
    x_64 = 'b000001010;
    x_65 = 'b000011001;
    x_66 = 'b000001110;
    x_67 = 'b000010110;
    x_68 = 'b000001010;
    x_69 = 'b000000110;
    x_70 = 'b000000011;
    x_71 = 'b000100001;
    x_72 = 'b000010111;
    x_73 = 'b000010111;
    x_74 = 'b000010101;
    x_75 = 'b000001111;
    x_76 = 'b000010001;
    x_77 = 'b000000110;
    x_78 = 'b000100000;
    x_79 = 'b000011011;
    x_80 = 'b000010110;
    x_81 = 'b000011100;
    x_82 = 'b000010100;
    x_83 = 'b000010110;
    x_84 = 'b000011010;
    x_85 = 'b111111000;
    x_86 = 'b111111111;
    x_87 = 'b000000100;
    x_88 = 'b111111100;
    x_89 = 'b111111101;
    x_90 = 'b111111100;
    x_91 = 'b111111010;
    x_92 = 'b000000110;
    x_93 = 'b111101011;
    x_94 = 'b000001100;
    x_95 = 'b000000011;
    x_96 = 'b000000110;
    x_97 = 'b000000100;
    x_98 = 'b111111101;
    x_99 = 'b111110101;
    x_100 = 'b111111011;
    x_101 = 'b111010111;
    x_102 = 'b111110101;
    x_103 = 'b000000001;
    x_104 = 'b000000001;
    x_105 = 'b111110110;
    x_106 = 'b000001100;
    x_107 = 'b111101111;
    x_108 = 'b000010010;
    x_109 = 'b000010101;
    x_110 = 'b000010010;
    x_111 = 'b000010010;
    x_112 = 'b000010101;
    x_113 = 'b000010001;
    x_114 = 'b000010101;
    x_115 = 'b000011010;
    x_116 = 'b000011001;
    x_117 = 'b000010111;
    x_118 = 'b000011001;
    x_119 = 'b000010000;
    x_120 = 'b000010010;
    x_121 = 'b000010010;
    x_122 = 'b000100100;
    x_123 = 'b000011111;
    x_124 = 'b000001111;
    x_125 = 'b000100011;
    x_126 = 'b000011101;
    x_127 = 'b000010000;
    x_128 = 'b000001010;
    x_129 = 'b000011001;
    x_130 = 'b000001110;
    x_131 = 'b000010110;
    x_132 = 'b000001010;
    x_133 = 'b000000110;
    x_134 = 'b000000011;
    x_135 = 'b000100001;
    x_136 = 'b000010111;
    x_137 = 'b000010111;
    x_138 = 'b000010101;
    x_139 = 'b000001111;
    x_140 = 'b000010001;
    x_141 = 'b000000110;
    x_142 = 'b000100000;
    x_143 = 'b000011011;
    x_144 = 'b000010110;
    x_145 = 'b000011100;
    x_146 = 'b000010100;
    x_147 = 'b000010110;
    x_148 = 'b000011010;
    x_149 = 'b111111000;
    x_150 = 'b111111111;
    x_151 = 'b000000100;
    x_152 = 'b111111100;
    x_153 = 'b111111101;
    x_154 = 'b111111100;
    x_155 = 'b111111010;
    x_156 = 'b000000110;
    x_157 = 'b111101011;
    x_158 = 'b000001100;
    x_159 = 'b000000011;
    x_160 = 'b000000110;
    x_161 = 'b000000100;
    x_162 = 'b111111101;
    x_163 = 'b111110101;
    x_164 = 'b111111011;
    x_165 = 'b111010111;
    x_166 = 'b111110101;
    x_167 = 'b000000001;
    x_168 = 'b000000001;
    x_169 = 'b111110110;
    x_170 = 'b000001100;
    x_171 = 'b111101111;
    x_172 = 'b000010010;
    x_173 = 'b000010101;
    x_174 = 'b000010010;
    x_175 = 'b000010010;
    x_176 = 'b000010101;
    x_177 = 'b000010001;
    x_178 = 'b000010101;
    x_179 = 'b000011010;
    x_180 = 'b000011001;
    x_181 = 'b000010111;
    x_182 = 'b000011001;
    x_183 = 'b000010000;
    x_184 = 'b000010010;
    x_185 = 'b000010010;
    x_186 = 'b000100100;
    x_187 = 'b000011111;
    x_188 = 'b000001111;
    x_189 = 'b000100011;
    x_190 = 'b000011101;
    x_191 = 'b000010000;
    x_192 = 'b000001010;
    x_193 = 'b000011001;
    x_194 = 'b000001110;
    x_195 = 'b000010110;
    x_196 = 'b000001010;
    x_197 = 'b000000110;
    x_198 = 'b000000011;
    x_199 = 'b000100001;
    x_200 = 'b000010111;
    x_201 = 'b000010111;
    x_202 = 'b000010101;
    x_203 = 'b000001111;
    x_204 = 'b000010001;
    x_205 = 'b000000110;
    x_206 = 'b000100000;
    x_207 = 'b000011011;
    x_208 = 'b000010110;
    x_209 = 'b000011100;
    x_210 = 'b000010100;
    x_211 = 'b000010110;
    x_212 = 'b000011010;
    x_213 = 'b111111000;
    x_214 = 'b111111111;
    x_215 = 'b000000100;
    x_216 = 'b111111100;
    x_217 = 'b111111101;
    x_218 = 'b111111100;
    x_219 = 'b111111010;
    x_220 = 'b000000110;
    x_221 = 'b111101011;
    x_222 = 'b000001100;
    x_223 = 'b000000011;
    x_224 = 'b000000110;
    x_225 = 'b000000100;
    x_226 = 'b111111101;
    x_227 = 'b111110101;
    x_228 = 'b111111011;
    x_229 = 'b111010111;
    x_230 = 'b111110101;
    x_231 = 'b000000001;
    x_232 = 'b000000001;
    x_233 = 'b111110110;
    x_234 = 'b000001100;
    x_235 = 'b111101111;
    x_236 = 'b000010010;
    x_237 = 'b000010101;
    x_238 = 'b000010010;
    x_239 = 'b000010010;
    x_240 = 'b000010101;
    x_241 = 'b000010001;
    x_242 = 'b000010101;
    x_243 = 'b000011010;
    x_244 = 'b000011001;
    x_245 = 'b000010111;
    x_246 = 'b000011001;
    x_247 = 'b000010000;
    x_248 = 'b000010010;
    x_249 = 'b000010010;
    x_250 = 'b000100100;
    x_251 = 'b000011111;
    x_252 = 'b000001111;
    x_253 = 'b000100011;
    x_254 = 'b000011101;
    x_255 = 'b000010000;

    h_0 = 'b000001010;
    h_1 = 'b000011001;
    h_2 = 'b000001110;
    h_3 = 'b000010110;
    h_4 = 'b000001010;
    h_5 = 'b000000110;
    h_6 = 'b000000011;
    h_7 = 'b000100001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111111010;
    x_1 = 'b000000110;
    x_2 = 'b000000001;
    x_3 = 'b000001001;
    x_4 = 'b000000000;
    x_5 = 'b111111110;
    x_6 = 'b000000001;
    x_7 = 'b000000101;
    x_8 = 'b111111111;
    x_9 = 'b000001000;
    x_10 = 'b000001001;
    x_11 = 'b000000001;
    x_12 = 'b000000110;
    x_13 = 'b000000011;
    x_14 = 'b000000101;
    x_15 = 'b000001001;
    x_16 = 'b000001000;
    x_17 = 'b000001111;
    x_18 = 'b000000110;
    x_19 = 'b000001001;
    x_20 = 'b000010011;
    x_21 = 'b111111110;
    x_22 = 'b000000100;
    x_23 = 'b000001010;
    x_24 = 'b000000001;
    x_25 = 'b000000001;
    x_26 = 'b111111011;
    x_27 = 'b111111101;
    x_28 = 'b000001100;
    x_29 = 'b111111011;
    x_30 = 'b000001100;
    x_31 = 'b000000010;
    x_32 = 'b000000000;
    x_33 = 'b000000000;
    x_34 = 'b111111001;
    x_35 = 'b111110010;
    x_36 = 'b111111111;
    x_37 = 'b111011111;
    x_38 = 'b000000100;
    x_39 = 'b000000111;
    x_40 = 'b000010101;
    x_41 = 'b111101111;
    x_42 = 'b000010010;
    x_43 = 'b111110101;
    x_44 = 'b000010001;
    x_45 = 'b000100100;
    x_46 = 'b000010000;
    x_47 = 'b000010000;
    x_48 = 'b000010101;
    x_49 = 'b000010000;
    x_50 = 'b000001111;
    x_51 = 'b000010011;
    x_52 = 'b000010010;
    x_53 = 'b000010010;
    x_54 = 'b000011110;
    x_55 = 'b000010001;
    x_56 = 'b000010111;
    x_57 = 'b000010001;
    x_58 = 'b000011101;
    x_59 = 'b000011100;
    x_60 = 'b000001001;
    x_61 = 'b000011010;
    x_62 = 'b000010001;
    x_63 = 'b000001000;
    x_64 = 'b111111010;
    x_65 = 'b000000110;
    x_66 = 'b000000001;
    x_67 = 'b000001001;
    x_68 = 'b000000000;
    x_69 = 'b111111110;
    x_70 = 'b000000001;
    x_71 = 'b000000101;
    x_72 = 'b111111111;
    x_73 = 'b000001000;
    x_74 = 'b000001001;
    x_75 = 'b000000001;
    x_76 = 'b000000110;
    x_77 = 'b000000011;
    x_78 = 'b000000101;
    x_79 = 'b000001001;
    x_80 = 'b000001000;
    x_81 = 'b000001111;
    x_82 = 'b000000110;
    x_83 = 'b000001001;
    x_84 = 'b000010011;
    x_85 = 'b111111110;
    x_86 = 'b000000100;
    x_87 = 'b000001010;
    x_88 = 'b000000001;
    x_89 = 'b000000001;
    x_90 = 'b111111011;
    x_91 = 'b111111101;
    x_92 = 'b000001100;
    x_93 = 'b111111011;
    x_94 = 'b000001100;
    x_95 = 'b000000010;
    x_96 = 'b000000000;
    x_97 = 'b000000000;
    x_98 = 'b111111001;
    x_99 = 'b111110010;
    x_100 = 'b111111111;
    x_101 = 'b111011111;
    x_102 = 'b000000100;
    x_103 = 'b000000111;
    x_104 = 'b000010101;
    x_105 = 'b111101111;
    x_106 = 'b000010010;
    x_107 = 'b111110101;
    x_108 = 'b000010001;
    x_109 = 'b000100100;
    x_110 = 'b000010000;
    x_111 = 'b000010000;
    x_112 = 'b000010101;
    x_113 = 'b000010000;
    x_114 = 'b000001111;
    x_115 = 'b000010011;
    x_116 = 'b000010010;
    x_117 = 'b000010010;
    x_118 = 'b000011110;
    x_119 = 'b000010001;
    x_120 = 'b000010111;
    x_121 = 'b000010001;
    x_122 = 'b000011101;
    x_123 = 'b000011100;
    x_124 = 'b000001001;
    x_125 = 'b000011010;
    x_126 = 'b000010001;
    x_127 = 'b000001000;
    x_128 = 'b111111010;
    x_129 = 'b000000110;
    x_130 = 'b000000001;
    x_131 = 'b000001001;
    x_132 = 'b000000000;
    x_133 = 'b111111110;
    x_134 = 'b000000001;
    x_135 = 'b000000101;
    x_136 = 'b111111111;
    x_137 = 'b000001000;
    x_138 = 'b000001001;
    x_139 = 'b000000001;
    x_140 = 'b000000110;
    x_141 = 'b000000011;
    x_142 = 'b000000101;
    x_143 = 'b000001001;
    x_144 = 'b000001000;
    x_145 = 'b000001111;
    x_146 = 'b000000110;
    x_147 = 'b000001001;
    x_148 = 'b000010011;
    x_149 = 'b111111110;
    x_150 = 'b000000100;
    x_151 = 'b000001010;
    x_152 = 'b000000001;
    x_153 = 'b000000001;
    x_154 = 'b111111011;
    x_155 = 'b111111101;
    x_156 = 'b000001100;
    x_157 = 'b111111011;
    x_158 = 'b000001100;
    x_159 = 'b000000010;
    x_160 = 'b000000000;
    x_161 = 'b000000000;
    x_162 = 'b111111001;
    x_163 = 'b111110010;
    x_164 = 'b111111111;
    x_165 = 'b111011111;
    x_166 = 'b000000100;
    x_167 = 'b000000111;
    x_168 = 'b000010101;
    x_169 = 'b111101111;
    x_170 = 'b000010010;
    x_171 = 'b111110101;
    x_172 = 'b000010001;
    x_173 = 'b000100100;
    x_174 = 'b000010000;
    x_175 = 'b000010000;
    x_176 = 'b000010101;
    x_177 = 'b000010000;
    x_178 = 'b000001111;
    x_179 = 'b000010011;
    x_180 = 'b000010010;
    x_181 = 'b000010010;
    x_182 = 'b000011110;
    x_183 = 'b000010001;
    x_184 = 'b000010111;
    x_185 = 'b000010001;
    x_186 = 'b000011101;
    x_187 = 'b000011100;
    x_188 = 'b000001001;
    x_189 = 'b000011010;
    x_190 = 'b000010001;
    x_191 = 'b000001000;
    x_192 = 'b111111010;
    x_193 = 'b000000110;
    x_194 = 'b000000001;
    x_195 = 'b000001001;
    x_196 = 'b000000000;
    x_197 = 'b111111110;
    x_198 = 'b000000001;
    x_199 = 'b000000101;
    x_200 = 'b111111111;
    x_201 = 'b000001000;
    x_202 = 'b000001001;
    x_203 = 'b000000001;
    x_204 = 'b000000110;
    x_205 = 'b000000011;
    x_206 = 'b000000101;
    x_207 = 'b000001001;
    x_208 = 'b000001000;
    x_209 = 'b000001111;
    x_210 = 'b000000110;
    x_211 = 'b000001001;
    x_212 = 'b000010011;
    x_213 = 'b111111110;
    x_214 = 'b000000100;
    x_215 = 'b000001010;
    x_216 = 'b000000001;
    x_217 = 'b000000001;
    x_218 = 'b111111011;
    x_219 = 'b111111101;
    x_220 = 'b000001100;
    x_221 = 'b111111011;
    x_222 = 'b000001100;
    x_223 = 'b000000010;
    x_224 = 'b000000000;
    x_225 = 'b000000000;
    x_226 = 'b111111001;
    x_227 = 'b111110010;
    x_228 = 'b111111111;
    x_229 = 'b111011111;
    x_230 = 'b000000100;
    x_231 = 'b000000111;
    x_232 = 'b000010101;
    x_233 = 'b111101111;
    x_234 = 'b000010010;
    x_235 = 'b111110101;
    x_236 = 'b000010001;
    x_237 = 'b000100100;
    x_238 = 'b000010000;
    x_239 = 'b000010000;
    x_240 = 'b000010101;
    x_241 = 'b000010000;
    x_242 = 'b000001111;
    x_243 = 'b000010011;
    x_244 = 'b000010010;
    x_245 = 'b000010010;
    x_246 = 'b000011110;
    x_247 = 'b000010001;
    x_248 = 'b000010111;
    x_249 = 'b000010001;
    x_250 = 'b000011101;
    x_251 = 'b000011100;
    x_252 = 'b000001001;
    x_253 = 'b000011010;
    x_254 = 'b000010001;
    x_255 = 'b000001000;

    h_0 = 'b111111010;
    h_1 = 'b000000110;
    h_2 = 'b000000001;
    h_3 = 'b000001001;
    h_4 = 'b000000000;
    h_5 = 'b111111110;
    h_6 = 'b000000001;
    h_7 = 'b000000101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000001001;
    x_1 = 'b000001001;
    x_2 = 'b111111110;
    x_3 = 'b000000001;
    x_4 = 'b111111000;
    x_5 = 'b111110111;
    x_6 = 'b111111100;
    x_7 = 'b000011000;
    x_8 = 'b000000110;
    x_9 = 'b000001001;
    x_10 = 'b000001001;
    x_11 = 'b111111011;
    x_12 = 'b111111101;
    x_13 = 'b111111001;
    x_14 = 'b000010011;
    x_15 = 'b000010001;
    x_16 = 'b000001100;
    x_17 = 'b000001111;
    x_18 = 'b000000000;
    x_19 = 'b111111111;
    x_20 = 'b000001010;
    x_21 = 'b000000101;
    x_22 = 'b000001010;
    x_23 = 'b000001110;
    x_24 = 'b000001011;
    x_25 = 'b000001011;
    x_26 = 'b111110111;
    x_27 = 'b111111010;
    x_28 = 'b000001000;
    x_29 = 'b000000010;
    x_30 = 'b000010101;
    x_31 = 'b111111010;
    x_32 = 'b111111010;
    x_33 = 'b111111001;
    x_34 = 'b111110010;
    x_35 = 'b111101100;
    x_36 = 'b111110110;
    x_37 = 'b111011100;
    x_38 = 'b000010000;
    x_39 = 'b111110110;
    x_40 = 'b000011010;
    x_41 = 'b111100100;
    x_42 = 'b000001111;
    x_43 = 'b000011000;
    x_44 = 'b000010110;
    x_45 = 'b000010000;
    x_46 = 'b000010110;
    x_47 = 'b000010100;
    x_48 = 'b000010101;
    x_49 = 'b000001111;
    x_50 = 'b000000101;
    x_51 = 'b000000011;
    x_52 = 'b111111110;
    x_53 = 'b111111101;
    x_54 = 'b000001010;
    x_55 = 'b000010110;
    x_56 = 'b000011001;
    x_57 = 'b000001001;
    x_58 = 'b000001001;
    x_59 = 'b000001000;
    x_60 = 'b000001010;
    x_61 = 'b000010110;
    x_62 = 'b000001010;
    x_63 = 'b000001001;
    x_64 = 'b000001001;
    x_65 = 'b000001001;
    x_66 = 'b111111110;
    x_67 = 'b000000001;
    x_68 = 'b111111000;
    x_69 = 'b111110111;
    x_70 = 'b111111100;
    x_71 = 'b000011000;
    x_72 = 'b000000110;
    x_73 = 'b000001001;
    x_74 = 'b000001001;
    x_75 = 'b111111011;
    x_76 = 'b111111101;
    x_77 = 'b111111001;
    x_78 = 'b000010011;
    x_79 = 'b000010001;
    x_80 = 'b000001100;
    x_81 = 'b000001111;
    x_82 = 'b000000000;
    x_83 = 'b111111111;
    x_84 = 'b000001010;
    x_85 = 'b000000101;
    x_86 = 'b000001010;
    x_87 = 'b000001110;
    x_88 = 'b000001011;
    x_89 = 'b000001011;
    x_90 = 'b111110111;
    x_91 = 'b111111010;
    x_92 = 'b000001000;
    x_93 = 'b000000010;
    x_94 = 'b000010101;
    x_95 = 'b111111010;
    x_96 = 'b111111010;
    x_97 = 'b111111001;
    x_98 = 'b111110010;
    x_99 = 'b111101100;
    x_100 = 'b111110110;
    x_101 = 'b111011100;
    x_102 = 'b000010000;
    x_103 = 'b111110110;
    x_104 = 'b000011010;
    x_105 = 'b111100100;
    x_106 = 'b000001111;
    x_107 = 'b000011000;
    x_108 = 'b000010110;
    x_109 = 'b000010000;
    x_110 = 'b000010110;
    x_111 = 'b000010100;
    x_112 = 'b000010101;
    x_113 = 'b000001111;
    x_114 = 'b000000101;
    x_115 = 'b000000011;
    x_116 = 'b111111110;
    x_117 = 'b111111101;
    x_118 = 'b000001010;
    x_119 = 'b000010110;
    x_120 = 'b000011001;
    x_121 = 'b000001001;
    x_122 = 'b000001001;
    x_123 = 'b000001000;
    x_124 = 'b000001010;
    x_125 = 'b000010110;
    x_126 = 'b000001010;
    x_127 = 'b000001001;
    x_128 = 'b000001001;
    x_129 = 'b000001001;
    x_130 = 'b111111110;
    x_131 = 'b000000001;
    x_132 = 'b111111000;
    x_133 = 'b111110111;
    x_134 = 'b111111100;
    x_135 = 'b000011000;
    x_136 = 'b000000110;
    x_137 = 'b000001001;
    x_138 = 'b000001001;
    x_139 = 'b111111011;
    x_140 = 'b111111101;
    x_141 = 'b111111001;
    x_142 = 'b000010011;
    x_143 = 'b000010001;
    x_144 = 'b000001100;
    x_145 = 'b000001111;
    x_146 = 'b000000000;
    x_147 = 'b111111111;
    x_148 = 'b000001010;
    x_149 = 'b000000101;
    x_150 = 'b000001010;
    x_151 = 'b000001110;
    x_152 = 'b000001011;
    x_153 = 'b000001011;
    x_154 = 'b111110111;
    x_155 = 'b111111010;
    x_156 = 'b000001000;
    x_157 = 'b000000010;
    x_158 = 'b000010101;
    x_159 = 'b111111010;
    x_160 = 'b111111010;
    x_161 = 'b111111001;
    x_162 = 'b111110010;
    x_163 = 'b111101100;
    x_164 = 'b111110110;
    x_165 = 'b111011100;
    x_166 = 'b000010000;
    x_167 = 'b111110110;
    x_168 = 'b000011010;
    x_169 = 'b111100100;
    x_170 = 'b000001111;
    x_171 = 'b000011000;
    x_172 = 'b000010110;
    x_173 = 'b000010000;
    x_174 = 'b000010110;
    x_175 = 'b000010100;
    x_176 = 'b000010101;
    x_177 = 'b000001111;
    x_178 = 'b000000101;
    x_179 = 'b000000011;
    x_180 = 'b111111110;
    x_181 = 'b111111101;
    x_182 = 'b000001010;
    x_183 = 'b000010110;
    x_184 = 'b000011001;
    x_185 = 'b000001001;
    x_186 = 'b000001001;
    x_187 = 'b000001000;
    x_188 = 'b000001010;
    x_189 = 'b000010110;
    x_190 = 'b000001010;
    x_191 = 'b000001001;
    x_192 = 'b000001001;
    x_193 = 'b000001001;
    x_194 = 'b111111110;
    x_195 = 'b000000001;
    x_196 = 'b111111000;
    x_197 = 'b111110111;
    x_198 = 'b111111100;
    x_199 = 'b000011000;
    x_200 = 'b000000110;
    x_201 = 'b000001001;
    x_202 = 'b000001001;
    x_203 = 'b111111011;
    x_204 = 'b111111101;
    x_205 = 'b111111001;
    x_206 = 'b000010011;
    x_207 = 'b000010001;
    x_208 = 'b000001100;
    x_209 = 'b000001111;
    x_210 = 'b000000000;
    x_211 = 'b111111111;
    x_212 = 'b000001010;
    x_213 = 'b000000101;
    x_214 = 'b000001010;
    x_215 = 'b000001110;
    x_216 = 'b000001011;
    x_217 = 'b000001011;
    x_218 = 'b111110111;
    x_219 = 'b111111010;
    x_220 = 'b000001000;
    x_221 = 'b000000010;
    x_222 = 'b000010101;
    x_223 = 'b111111010;
    x_224 = 'b111111010;
    x_225 = 'b111111001;
    x_226 = 'b111110010;
    x_227 = 'b111101100;
    x_228 = 'b111110110;
    x_229 = 'b111011100;
    x_230 = 'b000010000;
    x_231 = 'b111110110;
    x_232 = 'b000011010;
    x_233 = 'b111100100;
    x_234 = 'b000001111;
    x_235 = 'b000011000;
    x_236 = 'b000010110;
    x_237 = 'b000010000;
    x_238 = 'b000010110;
    x_239 = 'b000010100;
    x_240 = 'b000010101;
    x_241 = 'b000001111;
    x_242 = 'b000000101;
    x_243 = 'b000000011;
    x_244 = 'b111111110;
    x_245 = 'b111111101;
    x_246 = 'b000001010;
    x_247 = 'b000010110;
    x_248 = 'b000011001;
    x_249 = 'b000001001;
    x_250 = 'b000001001;
    x_251 = 'b000001000;
    x_252 = 'b000001010;
    x_253 = 'b000010110;
    x_254 = 'b000001010;
    x_255 = 'b000001001;

    h_0 = 'b000001001;
    h_1 = 'b000001001;
    h_2 = 'b111111110;
    h_3 = 'b000000001;
    h_4 = 'b111111000;
    h_5 = 'b111110111;
    h_6 = 'b111111100;
    h_7 = 'b000011000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000001010;
    x_1 = 'b000001010;
    x_2 = 'b111111011;
    x_3 = 'b111111101;
    x_4 = 'b111110000;
    x_5 = 'b111101001;
    x_6 = 'b111110000;
    x_7 = 'b000011011;
    x_8 = 'b000001101;
    x_9 = 'b000001000;
    x_10 = 'b000000011;
    x_11 = 'b111111010;
    x_12 = 'b111110000;
    x_13 = 'b111101010;
    x_14 = 'b000010110;
    x_15 = 'b000010000;
    x_16 = 'b000001011;
    x_17 = 'b000001010;
    x_18 = 'b111110111;
    x_19 = 'b111110010;
    x_20 = 'b111111001;
    x_21 = 'b000000001;
    x_22 = 'b000000111;
    x_23 = 'b000001001;
    x_24 = 'b000001001;
    x_25 = 'b000001001;
    x_26 = 'b111111010;
    x_27 = 'b111111000;
    x_28 = 'b000000011;
    x_29 = 'b000000111;
    x_30 = 'b000010011;
    x_31 = 'b111111111;
    x_32 = 'b111111111;
    x_33 = 'b000000000;
    x_34 = 'b111110111;
    x_35 = 'b111101111;
    x_36 = 'b111111000;
    x_37 = 'b111011100;
    x_38 = 'b000010011;
    x_39 = 'b111110111;
    x_40 = 'b000011101;
    x_41 = 'b000000101;
    x_42 = 'b000101100;
    x_43 = 'b111111010;
    x_44 = 'b000100101;
    x_45 = 'b000000100;
    x_46 = 'b000100010;
    x_47 = 'b000011011;
    x_48 = 'b000011010;
    x_49 = 'b000010011;
    x_50 = 'b000001010;
    x_51 = 'b000000000;
    x_52 = 'b111111100;
    x_53 = 'b111110111;
    x_54 = 'b000000001;
    x_55 = 'b000100001;
    x_56 = 'b000100001;
    x_57 = 'b000001010;
    x_58 = 'b111111110;
    x_59 = 'b000000000;
    x_60 = 'b000010010;
    x_61 = 'b000010110;
    x_62 = 'b000000001;
    x_63 = 'b000001100;
    x_64 = 'b000001010;
    x_65 = 'b000001010;
    x_66 = 'b111111011;
    x_67 = 'b111111101;
    x_68 = 'b111110000;
    x_69 = 'b111101001;
    x_70 = 'b111110000;
    x_71 = 'b000011011;
    x_72 = 'b000001101;
    x_73 = 'b000001000;
    x_74 = 'b000000011;
    x_75 = 'b111111010;
    x_76 = 'b111110000;
    x_77 = 'b111101010;
    x_78 = 'b000010110;
    x_79 = 'b000010000;
    x_80 = 'b000001011;
    x_81 = 'b000001010;
    x_82 = 'b111110111;
    x_83 = 'b111110010;
    x_84 = 'b111111001;
    x_85 = 'b000000001;
    x_86 = 'b000000111;
    x_87 = 'b000001001;
    x_88 = 'b000001001;
    x_89 = 'b000001001;
    x_90 = 'b111111010;
    x_91 = 'b111111000;
    x_92 = 'b000000011;
    x_93 = 'b000000111;
    x_94 = 'b000010011;
    x_95 = 'b111111111;
    x_96 = 'b111111111;
    x_97 = 'b000000000;
    x_98 = 'b111110111;
    x_99 = 'b111101111;
    x_100 = 'b111111000;
    x_101 = 'b111011100;
    x_102 = 'b000010011;
    x_103 = 'b111110111;
    x_104 = 'b000011101;
    x_105 = 'b000000101;
    x_106 = 'b000101100;
    x_107 = 'b111111010;
    x_108 = 'b000100101;
    x_109 = 'b000000100;
    x_110 = 'b000100010;
    x_111 = 'b000011011;
    x_112 = 'b000011010;
    x_113 = 'b000010011;
    x_114 = 'b000001010;
    x_115 = 'b000000000;
    x_116 = 'b111111100;
    x_117 = 'b111110111;
    x_118 = 'b000000001;
    x_119 = 'b000100001;
    x_120 = 'b000100001;
    x_121 = 'b000001010;
    x_122 = 'b111111110;
    x_123 = 'b000000000;
    x_124 = 'b000010010;
    x_125 = 'b000010110;
    x_126 = 'b000000001;
    x_127 = 'b000001100;
    x_128 = 'b000001010;
    x_129 = 'b000001010;
    x_130 = 'b111111011;
    x_131 = 'b111111101;
    x_132 = 'b111110000;
    x_133 = 'b111101001;
    x_134 = 'b111110000;
    x_135 = 'b000011011;
    x_136 = 'b000001101;
    x_137 = 'b000001000;
    x_138 = 'b000000011;
    x_139 = 'b111111010;
    x_140 = 'b111110000;
    x_141 = 'b111101010;
    x_142 = 'b000010110;
    x_143 = 'b000010000;
    x_144 = 'b000001011;
    x_145 = 'b000001010;
    x_146 = 'b111110111;
    x_147 = 'b111110010;
    x_148 = 'b111111001;
    x_149 = 'b000000001;
    x_150 = 'b000000111;
    x_151 = 'b000001001;
    x_152 = 'b000001001;
    x_153 = 'b000001001;
    x_154 = 'b111111010;
    x_155 = 'b111111000;
    x_156 = 'b000000011;
    x_157 = 'b000000111;
    x_158 = 'b000010011;
    x_159 = 'b111111111;
    x_160 = 'b111111111;
    x_161 = 'b000000000;
    x_162 = 'b111110111;
    x_163 = 'b111101111;
    x_164 = 'b111111000;
    x_165 = 'b111011100;
    x_166 = 'b000010011;
    x_167 = 'b111110111;
    x_168 = 'b000011101;
    x_169 = 'b000000101;
    x_170 = 'b000101100;
    x_171 = 'b111111010;
    x_172 = 'b000100101;
    x_173 = 'b000000100;
    x_174 = 'b000100010;
    x_175 = 'b000011011;
    x_176 = 'b000011010;
    x_177 = 'b000010011;
    x_178 = 'b000001010;
    x_179 = 'b000000000;
    x_180 = 'b111111100;
    x_181 = 'b111110111;
    x_182 = 'b000000001;
    x_183 = 'b000100001;
    x_184 = 'b000100001;
    x_185 = 'b000001010;
    x_186 = 'b111111110;
    x_187 = 'b000000000;
    x_188 = 'b000010010;
    x_189 = 'b000010110;
    x_190 = 'b000000001;
    x_191 = 'b000001100;
    x_192 = 'b000001010;
    x_193 = 'b000001010;
    x_194 = 'b111111011;
    x_195 = 'b111111101;
    x_196 = 'b111110000;
    x_197 = 'b111101001;
    x_198 = 'b111110000;
    x_199 = 'b000011011;
    x_200 = 'b000001101;
    x_201 = 'b000001000;
    x_202 = 'b000000011;
    x_203 = 'b111111010;
    x_204 = 'b111110000;
    x_205 = 'b111101010;
    x_206 = 'b000010110;
    x_207 = 'b000010000;
    x_208 = 'b000001011;
    x_209 = 'b000001010;
    x_210 = 'b111110111;
    x_211 = 'b111110010;
    x_212 = 'b111111001;
    x_213 = 'b000000001;
    x_214 = 'b000000111;
    x_215 = 'b000001001;
    x_216 = 'b000001001;
    x_217 = 'b000001001;
    x_218 = 'b111111010;
    x_219 = 'b111111000;
    x_220 = 'b000000011;
    x_221 = 'b000000111;
    x_222 = 'b000010011;
    x_223 = 'b111111111;
    x_224 = 'b111111111;
    x_225 = 'b000000000;
    x_226 = 'b111110111;
    x_227 = 'b111101111;
    x_228 = 'b111111000;
    x_229 = 'b111011100;
    x_230 = 'b000010011;
    x_231 = 'b111110111;
    x_232 = 'b000011101;
    x_233 = 'b000000101;
    x_234 = 'b000101100;
    x_235 = 'b111111010;
    x_236 = 'b000100101;
    x_237 = 'b000000100;
    x_238 = 'b000100010;
    x_239 = 'b000011011;
    x_240 = 'b000011010;
    x_241 = 'b000010011;
    x_242 = 'b000001010;
    x_243 = 'b000000000;
    x_244 = 'b111111100;
    x_245 = 'b111110111;
    x_246 = 'b000000001;
    x_247 = 'b000100001;
    x_248 = 'b000100001;
    x_249 = 'b000001010;
    x_250 = 'b111111110;
    x_251 = 'b000000000;
    x_252 = 'b000010010;
    x_253 = 'b000010110;
    x_254 = 'b000000001;
    x_255 = 'b000001100;

    h_0 = 'b000001010;
    h_1 = 'b000001010;
    h_2 = 'b111111011;
    h_3 = 'b111111101;
    h_4 = 'b111110000;
    h_5 = 'b111101001;
    h_6 = 'b111110000;
    h_7 = 'b000011011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000011000;
    x_1 = 'b000011100;
    x_2 = 'b000001101;
    x_3 = 'b000001111;
    x_4 = 'b000000111;
    x_5 = 'b111111101;
    x_6 = 'b000000110;
    x_7 = 'b000101101;
    x_8 = 'b000011101;
    x_9 = 'b000011001;
    x_10 = 'b000010101;
    x_11 = 'b000001001;
    x_12 = 'b000000000;
    x_13 = 'b000000111;
    x_14 = 'b000100001;
    x_15 = 'b000011100;
    x_16 = 'b000010110;
    x_17 = 'b000010111;
    x_18 = 'b000000100;
    x_19 = 'b111111010;
    x_20 = 'b000000010;
    x_21 = 'b000010011;
    x_22 = 'b000011001;
    x_23 = 'b000011000;
    x_24 = 'b000011100;
    x_25 = 'b000011100;
    x_26 = 'b000001110;
    x_27 = 'b000001011;
    x_28 = 'b000010100;
    x_29 = 'b000011110;
    x_30 = 'b000100011;
    x_31 = 'b000010001;
    x_32 = 'b000010010;
    x_33 = 'b000010100;
    x_34 = 'b000001100;
    x_35 = 'b000000011;
    x_36 = 'b000001010;
    x_37 = 'b111101011;
    x_38 = 'b000100100;
    x_39 = 'b000010001;
    x_40 = 'b000100101;
    x_41 = 'b000010001;
    x_42 = 'b000111101;
    x_43 = 'b111110101;
    x_44 = 'b000101111;
    x_45 = 'b111111011;
    x_46 = 'b000101100;
    x_47 = 'b000011111;
    x_48 = 'b000011011;
    x_49 = 'b000010010;
    x_50 = 'b000000100;
    x_51 = 'b111101110;
    x_52 = 'b111101010;
    x_53 = 'b111100001;
    x_54 = 'b111101100;
    x_55 = 'b000100100;
    x_56 = 'b000100000;
    x_57 = 'b111111011;
    x_58 = 'b111011011;
    x_59 = 'b111100110;
    x_60 = 'b000011000;
    x_61 = 'b000010010;
    x_62 = 'b111110000;
    x_63 = 'b000001101;
    x_64 = 'b000011000;
    x_65 = 'b000011100;
    x_66 = 'b000001101;
    x_67 = 'b000001111;
    x_68 = 'b000000111;
    x_69 = 'b111111101;
    x_70 = 'b000000110;
    x_71 = 'b000101101;
    x_72 = 'b000011101;
    x_73 = 'b000011001;
    x_74 = 'b000010101;
    x_75 = 'b000001001;
    x_76 = 'b000000000;
    x_77 = 'b000000111;
    x_78 = 'b000100001;
    x_79 = 'b000011100;
    x_80 = 'b000010110;
    x_81 = 'b000010111;
    x_82 = 'b000000100;
    x_83 = 'b111111010;
    x_84 = 'b000000010;
    x_85 = 'b000010011;
    x_86 = 'b000011001;
    x_87 = 'b000011000;
    x_88 = 'b000011100;
    x_89 = 'b000011100;
    x_90 = 'b000001110;
    x_91 = 'b000001011;
    x_92 = 'b000010100;
    x_93 = 'b000011110;
    x_94 = 'b000100011;
    x_95 = 'b000010001;
    x_96 = 'b000010010;
    x_97 = 'b000010100;
    x_98 = 'b000001100;
    x_99 = 'b000000011;
    x_100 = 'b000001010;
    x_101 = 'b111101011;
    x_102 = 'b000100100;
    x_103 = 'b000010001;
    x_104 = 'b000100101;
    x_105 = 'b000010001;
    x_106 = 'b000111101;
    x_107 = 'b111110101;
    x_108 = 'b000101111;
    x_109 = 'b111111011;
    x_110 = 'b000101100;
    x_111 = 'b000011111;
    x_112 = 'b000011011;
    x_113 = 'b000010010;
    x_114 = 'b000000100;
    x_115 = 'b111101110;
    x_116 = 'b111101010;
    x_117 = 'b111100001;
    x_118 = 'b111101100;
    x_119 = 'b000100100;
    x_120 = 'b000100000;
    x_121 = 'b111111011;
    x_122 = 'b111011011;
    x_123 = 'b111100110;
    x_124 = 'b000011000;
    x_125 = 'b000010010;
    x_126 = 'b111110000;
    x_127 = 'b000001101;
    x_128 = 'b000011000;
    x_129 = 'b000011100;
    x_130 = 'b000001101;
    x_131 = 'b000001111;
    x_132 = 'b000000111;
    x_133 = 'b111111101;
    x_134 = 'b000000110;
    x_135 = 'b000101101;
    x_136 = 'b000011101;
    x_137 = 'b000011001;
    x_138 = 'b000010101;
    x_139 = 'b000001001;
    x_140 = 'b000000000;
    x_141 = 'b000000111;
    x_142 = 'b000100001;
    x_143 = 'b000011100;
    x_144 = 'b000010110;
    x_145 = 'b000010111;
    x_146 = 'b000000100;
    x_147 = 'b111111010;
    x_148 = 'b000000010;
    x_149 = 'b000010011;
    x_150 = 'b000011001;
    x_151 = 'b000011000;
    x_152 = 'b000011100;
    x_153 = 'b000011100;
    x_154 = 'b000001110;
    x_155 = 'b000001011;
    x_156 = 'b000010100;
    x_157 = 'b000011110;
    x_158 = 'b000100011;
    x_159 = 'b000010001;
    x_160 = 'b000010010;
    x_161 = 'b000010100;
    x_162 = 'b000001100;
    x_163 = 'b000000011;
    x_164 = 'b000001010;
    x_165 = 'b111101011;
    x_166 = 'b000100100;
    x_167 = 'b000010001;
    x_168 = 'b000100101;
    x_169 = 'b000010001;
    x_170 = 'b000111101;
    x_171 = 'b111110101;
    x_172 = 'b000101111;
    x_173 = 'b111111011;
    x_174 = 'b000101100;
    x_175 = 'b000011111;
    x_176 = 'b000011011;
    x_177 = 'b000010010;
    x_178 = 'b000000100;
    x_179 = 'b111101110;
    x_180 = 'b111101010;
    x_181 = 'b111100001;
    x_182 = 'b111101100;
    x_183 = 'b000100100;
    x_184 = 'b000100000;
    x_185 = 'b111111011;
    x_186 = 'b111011011;
    x_187 = 'b111100110;
    x_188 = 'b000011000;
    x_189 = 'b000010010;
    x_190 = 'b111110000;
    x_191 = 'b000001101;
    x_192 = 'b000011000;
    x_193 = 'b000011100;
    x_194 = 'b000001101;
    x_195 = 'b000001111;
    x_196 = 'b000000111;
    x_197 = 'b111111101;
    x_198 = 'b000000110;
    x_199 = 'b000101101;
    x_200 = 'b000011101;
    x_201 = 'b000011001;
    x_202 = 'b000010101;
    x_203 = 'b000001001;
    x_204 = 'b000000000;
    x_205 = 'b000000111;
    x_206 = 'b000100001;
    x_207 = 'b000011100;
    x_208 = 'b000010110;
    x_209 = 'b000010111;
    x_210 = 'b000000100;
    x_211 = 'b111111010;
    x_212 = 'b000000010;
    x_213 = 'b000010011;
    x_214 = 'b000011001;
    x_215 = 'b000011000;
    x_216 = 'b000011100;
    x_217 = 'b000011100;
    x_218 = 'b000001110;
    x_219 = 'b000001011;
    x_220 = 'b000010100;
    x_221 = 'b000011110;
    x_222 = 'b000100011;
    x_223 = 'b000010001;
    x_224 = 'b000010010;
    x_225 = 'b000010100;
    x_226 = 'b000001100;
    x_227 = 'b000000011;
    x_228 = 'b000001010;
    x_229 = 'b111101011;
    x_230 = 'b000100100;
    x_231 = 'b000010001;
    x_232 = 'b000100101;
    x_233 = 'b000010001;
    x_234 = 'b000111101;
    x_235 = 'b111110101;
    x_236 = 'b000101111;
    x_237 = 'b111111011;
    x_238 = 'b000101100;
    x_239 = 'b000011111;
    x_240 = 'b000011011;
    x_241 = 'b000010010;
    x_242 = 'b000000100;
    x_243 = 'b111101110;
    x_244 = 'b111101010;
    x_245 = 'b111100001;
    x_246 = 'b111101100;
    x_247 = 'b000100100;
    x_248 = 'b000100000;
    x_249 = 'b111111011;
    x_250 = 'b111011011;
    x_251 = 'b111100110;
    x_252 = 'b000011000;
    x_253 = 'b000010010;
    x_254 = 'b111110000;
    x_255 = 'b000001101;

    h_0 = 'b000011000;
    h_1 = 'b000011100;
    h_2 = 'b000001101;
    h_3 = 'b000001111;
    h_4 = 'b000000111;
    h_5 = 'b111111101;
    h_6 = 'b000000110;
    h_7 = 'b000101101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000011111;
    x_1 = 'b000100000;
    x_2 = 'b000001110;
    x_3 = 'b000010111;
    x_4 = 'b000001011;
    x_5 = 'b000000000;
    x_6 = 'b000000000;
    x_7 = 'b000101001;
    x_8 = 'b000011001;
    x_9 = 'b000010110;
    x_10 = 'b000010010;
    x_11 = 'b111111111;
    x_12 = 'b111110111;
    x_13 = 'b111110010;
    x_14 = 'b000011110;
    x_15 = 'b000010011;
    x_16 = 'b000001100;
    x_17 = 'b000001001;
    x_18 = 'b111110101;
    x_19 = 'b111101000;
    x_20 = 'b111101001;
    x_21 = 'b000010100;
    x_22 = 'b000011010;
    x_23 = 'b000011011;
    x_24 = 'b000010111;
    x_25 = 'b000011000;
    x_26 = 'b000001100;
    x_27 = 'b000001010;
    x_28 = 'b000010011;
    x_29 = 'b000010111;
    x_30 = 'b000011001;
    x_31 = 'b000001010;
    x_32 = 'b000001101;
    x_33 = 'b000001110;
    x_34 = 'b000001000;
    x_35 = 'b111111110;
    x_36 = 'b000000100;
    x_37 = 'b111100010;
    x_38 = 'b000010100;
    x_39 = 'b111111111;
    x_40 = 'b000100010;
    x_41 = 'b111011000;
    x_42 = 'b000101001;
    x_43 = 'b000010100;
    x_44 = 'b000101010;
    x_45 = 'b111101011;
    x_46 = 'b000101000;
    x_47 = 'b000010010;
    x_48 = 'b000001000;
    x_49 = 'b000000001;
    x_50 = 'b111101111;
    x_51 = 'b111010101;
    x_52 = 'b111010000;
    x_53 = 'b111001100;
    x_54 = 'b111011111;
    x_55 = 'b000011011;
    x_56 = 'b000010101;
    x_57 = 'b111101010;
    x_58 = 'b111000011;
    x_59 = 'b111011000;
    x_60 = 'b000010101;
    x_61 = 'b000000101;
    x_62 = 'b111011010;
    x_63 = 'b000001101;
    x_64 = 'b000011111;
    x_65 = 'b000100000;
    x_66 = 'b000001110;
    x_67 = 'b000010111;
    x_68 = 'b000001011;
    x_69 = 'b000000000;
    x_70 = 'b000000000;
    x_71 = 'b000101001;
    x_72 = 'b000011001;
    x_73 = 'b000010110;
    x_74 = 'b000010010;
    x_75 = 'b111111111;
    x_76 = 'b111110111;
    x_77 = 'b111110010;
    x_78 = 'b000011110;
    x_79 = 'b000010011;
    x_80 = 'b000001100;
    x_81 = 'b000001001;
    x_82 = 'b111110101;
    x_83 = 'b111101000;
    x_84 = 'b111101001;
    x_85 = 'b000010100;
    x_86 = 'b000011010;
    x_87 = 'b000011011;
    x_88 = 'b000010111;
    x_89 = 'b000011000;
    x_90 = 'b000001100;
    x_91 = 'b000001010;
    x_92 = 'b000010011;
    x_93 = 'b000010111;
    x_94 = 'b000011001;
    x_95 = 'b000001010;
    x_96 = 'b000001101;
    x_97 = 'b000001110;
    x_98 = 'b000001000;
    x_99 = 'b111111110;
    x_100 = 'b000000100;
    x_101 = 'b111100010;
    x_102 = 'b000010100;
    x_103 = 'b111111111;
    x_104 = 'b000100010;
    x_105 = 'b111011000;
    x_106 = 'b000101001;
    x_107 = 'b000010100;
    x_108 = 'b000101010;
    x_109 = 'b111101011;
    x_110 = 'b000101000;
    x_111 = 'b000010010;
    x_112 = 'b000001000;
    x_113 = 'b000000001;
    x_114 = 'b111101111;
    x_115 = 'b111010101;
    x_116 = 'b111010000;
    x_117 = 'b111001100;
    x_118 = 'b111011111;
    x_119 = 'b000011011;
    x_120 = 'b000010101;
    x_121 = 'b111101010;
    x_122 = 'b111000011;
    x_123 = 'b111011000;
    x_124 = 'b000010101;
    x_125 = 'b000000101;
    x_126 = 'b111011010;
    x_127 = 'b000001101;
    x_128 = 'b000011111;
    x_129 = 'b000100000;
    x_130 = 'b000001110;
    x_131 = 'b000010111;
    x_132 = 'b000001011;
    x_133 = 'b000000000;
    x_134 = 'b000000000;
    x_135 = 'b000101001;
    x_136 = 'b000011001;
    x_137 = 'b000010110;
    x_138 = 'b000010010;
    x_139 = 'b111111111;
    x_140 = 'b111110111;
    x_141 = 'b111110010;
    x_142 = 'b000011110;
    x_143 = 'b000010011;
    x_144 = 'b000001100;
    x_145 = 'b000001001;
    x_146 = 'b111110101;
    x_147 = 'b111101000;
    x_148 = 'b111101001;
    x_149 = 'b000010100;
    x_150 = 'b000011010;
    x_151 = 'b000011011;
    x_152 = 'b000010111;
    x_153 = 'b000011000;
    x_154 = 'b000001100;
    x_155 = 'b000001010;
    x_156 = 'b000010011;
    x_157 = 'b000010111;
    x_158 = 'b000011001;
    x_159 = 'b000001010;
    x_160 = 'b000001101;
    x_161 = 'b000001110;
    x_162 = 'b000001000;
    x_163 = 'b111111110;
    x_164 = 'b000000100;
    x_165 = 'b111100010;
    x_166 = 'b000010100;
    x_167 = 'b111111111;
    x_168 = 'b000100010;
    x_169 = 'b111011000;
    x_170 = 'b000101001;
    x_171 = 'b000010100;
    x_172 = 'b000101010;
    x_173 = 'b111101011;
    x_174 = 'b000101000;
    x_175 = 'b000010010;
    x_176 = 'b000001000;
    x_177 = 'b000000001;
    x_178 = 'b111101111;
    x_179 = 'b111010101;
    x_180 = 'b111010000;
    x_181 = 'b111001100;
    x_182 = 'b111011111;
    x_183 = 'b000011011;
    x_184 = 'b000010101;
    x_185 = 'b111101010;
    x_186 = 'b111000011;
    x_187 = 'b111011000;
    x_188 = 'b000010101;
    x_189 = 'b000000101;
    x_190 = 'b111011010;
    x_191 = 'b000001101;
    x_192 = 'b000011111;
    x_193 = 'b000100000;
    x_194 = 'b000001110;
    x_195 = 'b000010111;
    x_196 = 'b000001011;
    x_197 = 'b000000000;
    x_198 = 'b000000000;
    x_199 = 'b000101001;
    x_200 = 'b000011001;
    x_201 = 'b000010110;
    x_202 = 'b000010010;
    x_203 = 'b111111111;
    x_204 = 'b111110111;
    x_205 = 'b111110010;
    x_206 = 'b000011110;
    x_207 = 'b000010011;
    x_208 = 'b000001100;
    x_209 = 'b000001001;
    x_210 = 'b111110101;
    x_211 = 'b111101000;
    x_212 = 'b111101001;
    x_213 = 'b000010100;
    x_214 = 'b000011010;
    x_215 = 'b000011011;
    x_216 = 'b000010111;
    x_217 = 'b000011000;
    x_218 = 'b000001100;
    x_219 = 'b000001010;
    x_220 = 'b000010011;
    x_221 = 'b000010111;
    x_222 = 'b000011001;
    x_223 = 'b000001010;
    x_224 = 'b000001101;
    x_225 = 'b000001110;
    x_226 = 'b000001000;
    x_227 = 'b111111110;
    x_228 = 'b000000100;
    x_229 = 'b111100010;
    x_230 = 'b000010100;
    x_231 = 'b111111111;
    x_232 = 'b000100010;
    x_233 = 'b111011000;
    x_234 = 'b000101001;
    x_235 = 'b000010100;
    x_236 = 'b000101010;
    x_237 = 'b111101011;
    x_238 = 'b000101000;
    x_239 = 'b000010010;
    x_240 = 'b000001000;
    x_241 = 'b000000001;
    x_242 = 'b111101111;
    x_243 = 'b111010101;
    x_244 = 'b111010000;
    x_245 = 'b111001100;
    x_246 = 'b111011111;
    x_247 = 'b000011011;
    x_248 = 'b000010101;
    x_249 = 'b111101010;
    x_250 = 'b111000011;
    x_251 = 'b111011000;
    x_252 = 'b000010101;
    x_253 = 'b000000101;
    x_254 = 'b111011010;
    x_255 = 'b000001101;

    h_0 = 'b000011111;
    h_1 = 'b000100000;
    h_2 = 'b000001110;
    h_3 = 'b000010111;
    h_4 = 'b000001011;
    h_5 = 'b000000000;
    h_6 = 'b000000000;
    h_7 = 'b000101001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000001100;
    x_1 = 'b000010101;
    x_2 = 'b111111110;
    x_3 = 'b000010010;
    x_4 = 'b000000110;
    x_5 = 'b111111000;
    x_6 = 'b111111011;
    x_7 = 'b000011101;
    x_8 = 'b000001110;
    x_9 = 'b000001101;
    x_10 = 'b000001001;
    x_11 = 'b111111011;
    x_12 = 'b111111000;
    x_13 = 'b111101101;
    x_14 = 'b000010110;
    x_15 = 'b000001011;
    x_16 = 'b000000010;
    x_17 = 'b111111111;
    x_18 = 'b111110001;
    x_19 = 'b111101100;
    x_20 = 'b111101111;
    x_21 = 'b000001000;
    x_22 = 'b000010000;
    x_23 = 'b000010011;
    x_24 = 'b000001110;
    x_25 = 'b000001110;
    x_26 = 'b000000101;
    x_27 = 'b000000010;
    x_28 = 'b000001101;
    x_29 = 'b000000101;
    x_30 = 'b000001111;
    x_31 = 'b000001000;
    x_32 = 'b000001010;
    x_33 = 'b000001110;
    x_34 = 'b000000101;
    x_35 = 'b111111000;
    x_36 = 'b000000011;
    x_37 = 'b111011100;
    x_38 = 'b111111111;
    x_39 = 'b000000110;
    x_40 = 'b000010011;
    x_41 = 'b111101100;
    x_42 = 'b000011010;
    x_43 = 'b111110000;
    x_44 = 'b000011000;
    x_45 = 'b111111101;
    x_46 = 'b000011000;
    x_47 = 'b000001101;
    x_48 = 'b000001000;
    x_49 = 'b111111010;
    x_50 = 'b111101110;
    x_51 = 'b111011011;
    x_52 = 'b111011001;
    x_53 = 'b111010101;
    x_54 = 'b111100011;
    x_55 = 'b000010110;
    x_56 = 'b000001111;
    x_57 = 'b111100101;
    x_58 = 'b111001001;
    x_59 = 'b111011001;
    x_60 = 'b000001111;
    x_61 = 'b111111000;
    x_62 = 'b111001110;
    x_63 = 'b000001011;
    x_64 = 'b000001100;
    x_65 = 'b000010101;
    x_66 = 'b111111110;
    x_67 = 'b000010010;
    x_68 = 'b000000110;
    x_69 = 'b111111000;
    x_70 = 'b111111011;
    x_71 = 'b000011101;
    x_72 = 'b000001110;
    x_73 = 'b000001101;
    x_74 = 'b000001001;
    x_75 = 'b111111011;
    x_76 = 'b111111000;
    x_77 = 'b111101101;
    x_78 = 'b000010110;
    x_79 = 'b000001011;
    x_80 = 'b000000010;
    x_81 = 'b111111111;
    x_82 = 'b111110001;
    x_83 = 'b111101100;
    x_84 = 'b111101111;
    x_85 = 'b000001000;
    x_86 = 'b000010000;
    x_87 = 'b000010011;
    x_88 = 'b000001110;
    x_89 = 'b000001110;
    x_90 = 'b000000101;
    x_91 = 'b000000010;
    x_92 = 'b000001101;
    x_93 = 'b000000101;
    x_94 = 'b000001111;
    x_95 = 'b000001000;
    x_96 = 'b000001010;
    x_97 = 'b000001110;
    x_98 = 'b000000101;
    x_99 = 'b111111000;
    x_100 = 'b000000011;
    x_101 = 'b111011100;
    x_102 = 'b111111111;
    x_103 = 'b000000110;
    x_104 = 'b000010011;
    x_105 = 'b111101100;
    x_106 = 'b000011010;
    x_107 = 'b111110000;
    x_108 = 'b000011000;
    x_109 = 'b111111101;
    x_110 = 'b000011000;
    x_111 = 'b000001101;
    x_112 = 'b000001000;
    x_113 = 'b111111010;
    x_114 = 'b111101110;
    x_115 = 'b111011011;
    x_116 = 'b111011001;
    x_117 = 'b111010101;
    x_118 = 'b111100011;
    x_119 = 'b000010110;
    x_120 = 'b000001111;
    x_121 = 'b111100101;
    x_122 = 'b111001001;
    x_123 = 'b111011001;
    x_124 = 'b000001111;
    x_125 = 'b111111000;
    x_126 = 'b111001110;
    x_127 = 'b000001011;
    x_128 = 'b000001100;
    x_129 = 'b000010101;
    x_130 = 'b111111110;
    x_131 = 'b000010010;
    x_132 = 'b000000110;
    x_133 = 'b111111000;
    x_134 = 'b111111011;
    x_135 = 'b000011101;
    x_136 = 'b000001110;
    x_137 = 'b000001101;
    x_138 = 'b000001001;
    x_139 = 'b111111011;
    x_140 = 'b111111000;
    x_141 = 'b111101101;
    x_142 = 'b000010110;
    x_143 = 'b000001011;
    x_144 = 'b000000010;
    x_145 = 'b111111111;
    x_146 = 'b111110001;
    x_147 = 'b111101100;
    x_148 = 'b111101111;
    x_149 = 'b000001000;
    x_150 = 'b000010000;
    x_151 = 'b000010011;
    x_152 = 'b000001110;
    x_153 = 'b000001110;
    x_154 = 'b000000101;
    x_155 = 'b000000010;
    x_156 = 'b000001101;
    x_157 = 'b000000101;
    x_158 = 'b000001111;
    x_159 = 'b000001000;
    x_160 = 'b000001010;
    x_161 = 'b000001110;
    x_162 = 'b000000101;
    x_163 = 'b111111000;
    x_164 = 'b000000011;
    x_165 = 'b111011100;
    x_166 = 'b111111111;
    x_167 = 'b000000110;
    x_168 = 'b000010011;
    x_169 = 'b111101100;
    x_170 = 'b000011010;
    x_171 = 'b111110000;
    x_172 = 'b000011000;
    x_173 = 'b111111101;
    x_174 = 'b000011000;
    x_175 = 'b000001101;
    x_176 = 'b000001000;
    x_177 = 'b111111010;
    x_178 = 'b111101110;
    x_179 = 'b111011011;
    x_180 = 'b111011001;
    x_181 = 'b111010101;
    x_182 = 'b111100011;
    x_183 = 'b000010110;
    x_184 = 'b000001111;
    x_185 = 'b111100101;
    x_186 = 'b111001001;
    x_187 = 'b111011001;
    x_188 = 'b000001111;
    x_189 = 'b111111000;
    x_190 = 'b111001110;
    x_191 = 'b000001011;
    x_192 = 'b000001100;
    x_193 = 'b000010101;
    x_194 = 'b111111110;
    x_195 = 'b000010010;
    x_196 = 'b000000110;
    x_197 = 'b111111000;
    x_198 = 'b111111011;
    x_199 = 'b000011101;
    x_200 = 'b000001110;
    x_201 = 'b000001101;
    x_202 = 'b000001001;
    x_203 = 'b111111011;
    x_204 = 'b111111000;
    x_205 = 'b111101101;
    x_206 = 'b000010110;
    x_207 = 'b000001011;
    x_208 = 'b000000010;
    x_209 = 'b111111111;
    x_210 = 'b111110001;
    x_211 = 'b111101100;
    x_212 = 'b111101111;
    x_213 = 'b000001000;
    x_214 = 'b000010000;
    x_215 = 'b000010011;
    x_216 = 'b000001110;
    x_217 = 'b000001110;
    x_218 = 'b000000101;
    x_219 = 'b000000010;
    x_220 = 'b000001101;
    x_221 = 'b000000101;
    x_222 = 'b000001111;
    x_223 = 'b000001000;
    x_224 = 'b000001010;
    x_225 = 'b000001110;
    x_226 = 'b000000101;
    x_227 = 'b111111000;
    x_228 = 'b000000011;
    x_229 = 'b111011100;
    x_230 = 'b111111111;
    x_231 = 'b000000110;
    x_232 = 'b000010011;
    x_233 = 'b111101100;
    x_234 = 'b000011010;
    x_235 = 'b111110000;
    x_236 = 'b000011000;
    x_237 = 'b111111101;
    x_238 = 'b000011000;
    x_239 = 'b000001101;
    x_240 = 'b000001000;
    x_241 = 'b111111010;
    x_242 = 'b111101110;
    x_243 = 'b111011011;
    x_244 = 'b111011001;
    x_245 = 'b111010101;
    x_246 = 'b111100011;
    x_247 = 'b000010110;
    x_248 = 'b000001111;
    x_249 = 'b111100101;
    x_250 = 'b111001001;
    x_251 = 'b111011001;
    x_252 = 'b000001111;
    x_253 = 'b111111000;
    x_254 = 'b111001110;
    x_255 = 'b000001011;

    h_0 = 'b000001100;
    h_1 = 'b000010101;
    h_2 = 'b111111110;
    h_3 = 'b000010010;
    h_4 = 'b000000110;
    h_5 = 'b111111000;
    h_6 = 'b111111011;
    h_7 = 'b000011101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111110101;
    x_1 = 'b111110101;
    x_2 = 'b111110000;
    x_3 = 'b111110001;
    x_4 = 'b111101100;
    x_5 = 'b111011100;
    x_6 = 'b111011000;
    x_7 = 'b111111101;
    x_8 = 'b111110001;
    x_9 = 'b111101101;
    x_10 = 'b111101100;
    x_11 = 'b111100101;
    x_12 = 'b111011101;
    x_13 = 'b111001000;
    x_14 = 'b111111101;
    x_15 = 'b111110011;
    x_16 = 'b111101110;
    x_17 = 'b111101001;
    x_18 = 'b111101001;
    x_19 = 'b111100101;
    x_20 = 'b111100001;
    x_21 = 'b111110110;
    x_22 = 'b111101010;
    x_23 = 'b111110001;
    x_24 = 'b111110101;
    x_25 = 'b111110110;
    x_26 = 'b111100110;
    x_27 = 'b111101010;
    x_28 = 'b111101010;
    x_29 = 'b111110111;
    x_30 = 'b111101001;
    x_31 = 'b111110110;
    x_32 = 'b111110001;
    x_33 = 'b111101001;
    x_34 = 'b111100011;
    x_35 = 'b111011110;
    x_36 = 'b111011100;
    x_37 = 'b111000011;
    x_38 = 'b111110001;
    x_39 = 'b111000111;
    x_40 = 'b111110000;
    x_41 = 'b111010101;
    x_42 = 'b111111100;
    x_43 = 'b111110110;
    x_44 = 'b111011100;
    x_45 = 'b111011000;
    x_46 = 'b111111110;
    x_47 = 'b111111000;
    x_48 = 'b111110011;
    x_49 = 'b111111010;
    x_50 = 'b111110001;
    x_51 = 'b111110010;
    x_52 = 'b111110010;
    x_53 = 'b111101000;
    x_54 = 'b111100100;
    x_55 = 'b111111000;
    x_56 = 'b111111110;
    x_57 = 'b111111110;
    x_58 = 'b000000010;
    x_59 = 'b000000001;
    x_60 = 'b111110110;
    x_61 = 'b111101110;
    x_62 = 'b111110100;
    x_63 = 'b111100001;
    x_64 = 'b111110101;
    x_65 = 'b111110101;
    x_66 = 'b111110000;
    x_67 = 'b111110001;
    x_68 = 'b111101100;
    x_69 = 'b111011100;
    x_70 = 'b111011000;
    x_71 = 'b111111101;
    x_72 = 'b111110001;
    x_73 = 'b111101101;
    x_74 = 'b111101100;
    x_75 = 'b111100101;
    x_76 = 'b111011101;
    x_77 = 'b111001000;
    x_78 = 'b111111101;
    x_79 = 'b111110011;
    x_80 = 'b111101110;
    x_81 = 'b111101001;
    x_82 = 'b111101001;
    x_83 = 'b111100101;
    x_84 = 'b111100001;
    x_85 = 'b111110110;
    x_86 = 'b111101010;
    x_87 = 'b111110001;
    x_88 = 'b111110101;
    x_89 = 'b111110110;
    x_90 = 'b111100110;
    x_91 = 'b111101010;
    x_92 = 'b111101010;
    x_93 = 'b111110111;
    x_94 = 'b111101001;
    x_95 = 'b111110110;
    x_96 = 'b111110001;
    x_97 = 'b111101001;
    x_98 = 'b111100011;
    x_99 = 'b111011110;
    x_100 = 'b111011100;
    x_101 = 'b111000011;
    x_102 = 'b111110001;
    x_103 = 'b111000111;
    x_104 = 'b111110000;
    x_105 = 'b111010101;
    x_106 = 'b111111100;
    x_107 = 'b111110110;
    x_108 = 'b111011100;
    x_109 = 'b111011000;
    x_110 = 'b111111110;
    x_111 = 'b111111000;
    x_112 = 'b111110011;
    x_113 = 'b111111010;
    x_114 = 'b111110001;
    x_115 = 'b111110010;
    x_116 = 'b111110010;
    x_117 = 'b111101000;
    x_118 = 'b111100100;
    x_119 = 'b111111000;
    x_120 = 'b111111110;
    x_121 = 'b111111110;
    x_122 = 'b000000010;
    x_123 = 'b000000001;
    x_124 = 'b111110110;
    x_125 = 'b111101110;
    x_126 = 'b111110100;
    x_127 = 'b111100001;
    x_128 = 'b111110101;
    x_129 = 'b111110101;
    x_130 = 'b111110000;
    x_131 = 'b111110001;
    x_132 = 'b111101100;
    x_133 = 'b111011100;
    x_134 = 'b111011000;
    x_135 = 'b111111101;
    x_136 = 'b111110001;
    x_137 = 'b111101101;
    x_138 = 'b111101100;
    x_139 = 'b111100101;
    x_140 = 'b111011101;
    x_141 = 'b111001000;
    x_142 = 'b111111101;
    x_143 = 'b111110011;
    x_144 = 'b111101110;
    x_145 = 'b111101001;
    x_146 = 'b111101001;
    x_147 = 'b111100101;
    x_148 = 'b111100001;
    x_149 = 'b111110110;
    x_150 = 'b111101010;
    x_151 = 'b111110001;
    x_152 = 'b111110101;
    x_153 = 'b111110110;
    x_154 = 'b111100110;
    x_155 = 'b111101010;
    x_156 = 'b111101010;
    x_157 = 'b111110111;
    x_158 = 'b111101001;
    x_159 = 'b111110110;
    x_160 = 'b111110001;
    x_161 = 'b111101001;
    x_162 = 'b111100011;
    x_163 = 'b111011110;
    x_164 = 'b111011100;
    x_165 = 'b111000011;
    x_166 = 'b111110001;
    x_167 = 'b111000111;
    x_168 = 'b111110000;
    x_169 = 'b111010101;
    x_170 = 'b111111100;
    x_171 = 'b111110110;
    x_172 = 'b111011100;
    x_173 = 'b111011000;
    x_174 = 'b111111110;
    x_175 = 'b111111000;
    x_176 = 'b111110011;
    x_177 = 'b111111010;
    x_178 = 'b111110001;
    x_179 = 'b111110010;
    x_180 = 'b111110010;
    x_181 = 'b111101000;
    x_182 = 'b111100100;
    x_183 = 'b111111000;
    x_184 = 'b111111110;
    x_185 = 'b111111110;
    x_186 = 'b000000010;
    x_187 = 'b000000001;
    x_188 = 'b111110110;
    x_189 = 'b111101110;
    x_190 = 'b111110100;
    x_191 = 'b111100001;
    x_192 = 'b111110101;
    x_193 = 'b111110101;
    x_194 = 'b111110000;
    x_195 = 'b111110001;
    x_196 = 'b111101100;
    x_197 = 'b111011100;
    x_198 = 'b111011000;
    x_199 = 'b111111101;
    x_200 = 'b111110001;
    x_201 = 'b111101101;
    x_202 = 'b111101100;
    x_203 = 'b111100101;
    x_204 = 'b111011101;
    x_205 = 'b111001000;
    x_206 = 'b111111101;
    x_207 = 'b111110011;
    x_208 = 'b111101110;
    x_209 = 'b111101001;
    x_210 = 'b111101001;
    x_211 = 'b111100101;
    x_212 = 'b111100001;
    x_213 = 'b111110110;
    x_214 = 'b111101010;
    x_215 = 'b111110001;
    x_216 = 'b111110101;
    x_217 = 'b111110110;
    x_218 = 'b111100110;
    x_219 = 'b111101010;
    x_220 = 'b111101010;
    x_221 = 'b111110111;
    x_222 = 'b111101001;
    x_223 = 'b111110110;
    x_224 = 'b111110001;
    x_225 = 'b111101001;
    x_226 = 'b111100011;
    x_227 = 'b111011110;
    x_228 = 'b111011100;
    x_229 = 'b111000011;
    x_230 = 'b111110001;
    x_231 = 'b111000111;
    x_232 = 'b111110000;
    x_233 = 'b111010101;
    x_234 = 'b111111100;
    x_235 = 'b111110110;
    x_236 = 'b111011100;
    x_237 = 'b111011000;
    x_238 = 'b111111110;
    x_239 = 'b111111000;
    x_240 = 'b111110011;
    x_241 = 'b111111010;
    x_242 = 'b111110001;
    x_243 = 'b111110010;
    x_244 = 'b111110010;
    x_245 = 'b111101000;
    x_246 = 'b111100100;
    x_247 = 'b111111000;
    x_248 = 'b111111110;
    x_249 = 'b111111110;
    x_250 = 'b000000010;
    x_251 = 'b000000001;
    x_252 = 'b111110110;
    x_253 = 'b111101110;
    x_254 = 'b111110100;
    x_255 = 'b111100001;

    h_0 = 'b111110101;
    h_1 = 'b111110101;
    h_2 = 'b111110000;
    h_3 = 'b111110001;
    h_4 = 'b111101100;
    h_5 = 'b111011100;
    h_6 = 'b111011000;
    h_7 = 'b111111101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111100100;
    x_1 = 'b111100100;
    x_2 = 'b111011111;
    x_3 = 'b111011101;
    x_4 = 'b111011011;
    x_5 = 'b111001111;
    x_6 = 'b111001111;
    x_7 = 'b111110101;
    x_8 = 'b111101000;
    x_9 = 'b111100010;
    x_10 = 'b111100010;
    x_11 = 'b111100000;
    x_12 = 'b111011110;
    x_13 = 'b111010001;
    x_14 = 'b111110110;
    x_15 = 'b111101110;
    x_16 = 'b111101001;
    x_17 = 'b111100101;
    x_18 = 'b111101010;
    x_19 = 'b111101101;
    x_20 = 'b111101010;
    x_21 = 'b111101010;
    x_22 = 'b111011111;
    x_23 = 'b111100110;
    x_24 = 'b111101011;
    x_25 = 'b111101011;
    x_26 = 'b111010110;
    x_27 = 'b111011011;
    x_28 = 'b111011110;
    x_29 = 'b111101000;
    x_30 = 'b111011010;
    x_31 = 'b111101000;
    x_32 = 'b111100000;
    x_33 = 'b111011000;
    x_34 = 'b111010011;
    x_35 = 'b111001101;
    x_36 = 'b111001111;
    x_37 = 'b111000100;
    x_38 = 'b111100011;
    x_39 = 'b111001100;
    x_40 = 'b111100100;
    x_41 = 'b111100110;
    x_42 = 'b111100001;
    x_43 = 'b111001010;
    x_44 = 'b111001111;
    x_45 = 'b111101001;
    x_46 = 'b111110010;
    x_47 = 'b111111000;
    x_48 = 'b111111001;
    x_49 = 'b000000100;
    x_50 = 'b111111001;
    x_51 = 'b111111111;
    x_52 = 'b000000000;
    x_53 = 'b111110111;
    x_54 = 'b111110101;
    x_55 = 'b111111110;
    x_56 = 'b000000110;
    x_57 = 'b000001011;
    x_58 = 'b000001111;
    x_59 = 'b000010000;
    x_60 = 'b111111010;
    x_61 = 'b111110111;
    x_62 = 'b000000001;
    x_63 = 'b111101101;
    x_64 = 'b111100100;
    x_65 = 'b111100100;
    x_66 = 'b111011111;
    x_67 = 'b111011101;
    x_68 = 'b111011011;
    x_69 = 'b111001111;
    x_70 = 'b111001111;
    x_71 = 'b111110101;
    x_72 = 'b111101000;
    x_73 = 'b111100010;
    x_74 = 'b111100010;
    x_75 = 'b111100000;
    x_76 = 'b111011110;
    x_77 = 'b111010001;
    x_78 = 'b111110110;
    x_79 = 'b111101110;
    x_80 = 'b111101001;
    x_81 = 'b111100101;
    x_82 = 'b111101010;
    x_83 = 'b111101101;
    x_84 = 'b111101010;
    x_85 = 'b111101010;
    x_86 = 'b111011111;
    x_87 = 'b111100110;
    x_88 = 'b111101011;
    x_89 = 'b111101011;
    x_90 = 'b111010110;
    x_91 = 'b111011011;
    x_92 = 'b111011110;
    x_93 = 'b111101000;
    x_94 = 'b111011010;
    x_95 = 'b111101000;
    x_96 = 'b111100000;
    x_97 = 'b111011000;
    x_98 = 'b111010011;
    x_99 = 'b111001101;
    x_100 = 'b111001111;
    x_101 = 'b111000100;
    x_102 = 'b111100011;
    x_103 = 'b111001100;
    x_104 = 'b111100100;
    x_105 = 'b111100110;
    x_106 = 'b111100001;
    x_107 = 'b111001010;
    x_108 = 'b111001111;
    x_109 = 'b111101001;
    x_110 = 'b111110010;
    x_111 = 'b111111000;
    x_112 = 'b111111001;
    x_113 = 'b000000100;
    x_114 = 'b111111001;
    x_115 = 'b111111111;
    x_116 = 'b000000000;
    x_117 = 'b111110111;
    x_118 = 'b111110101;
    x_119 = 'b111111110;
    x_120 = 'b000000110;
    x_121 = 'b000001011;
    x_122 = 'b000001111;
    x_123 = 'b000010000;
    x_124 = 'b111111010;
    x_125 = 'b111110111;
    x_126 = 'b000000001;
    x_127 = 'b111101101;
    x_128 = 'b111100100;
    x_129 = 'b111100100;
    x_130 = 'b111011111;
    x_131 = 'b111011101;
    x_132 = 'b111011011;
    x_133 = 'b111001111;
    x_134 = 'b111001111;
    x_135 = 'b111110101;
    x_136 = 'b111101000;
    x_137 = 'b111100010;
    x_138 = 'b111100010;
    x_139 = 'b111100000;
    x_140 = 'b111011110;
    x_141 = 'b111010001;
    x_142 = 'b111110110;
    x_143 = 'b111101110;
    x_144 = 'b111101001;
    x_145 = 'b111100101;
    x_146 = 'b111101010;
    x_147 = 'b111101101;
    x_148 = 'b111101010;
    x_149 = 'b111101010;
    x_150 = 'b111011111;
    x_151 = 'b111100110;
    x_152 = 'b111101011;
    x_153 = 'b111101011;
    x_154 = 'b111010110;
    x_155 = 'b111011011;
    x_156 = 'b111011110;
    x_157 = 'b111101000;
    x_158 = 'b111011010;
    x_159 = 'b111101000;
    x_160 = 'b111100000;
    x_161 = 'b111011000;
    x_162 = 'b111010011;
    x_163 = 'b111001101;
    x_164 = 'b111001111;
    x_165 = 'b111000100;
    x_166 = 'b111100011;
    x_167 = 'b111001100;
    x_168 = 'b111100100;
    x_169 = 'b111100110;
    x_170 = 'b111100001;
    x_171 = 'b111001010;
    x_172 = 'b111001111;
    x_173 = 'b111101001;
    x_174 = 'b111110010;
    x_175 = 'b111111000;
    x_176 = 'b111111001;
    x_177 = 'b000000100;
    x_178 = 'b111111001;
    x_179 = 'b111111111;
    x_180 = 'b000000000;
    x_181 = 'b111110111;
    x_182 = 'b111110101;
    x_183 = 'b111111110;
    x_184 = 'b000000110;
    x_185 = 'b000001011;
    x_186 = 'b000001111;
    x_187 = 'b000010000;
    x_188 = 'b111111010;
    x_189 = 'b111110111;
    x_190 = 'b000000001;
    x_191 = 'b111101101;
    x_192 = 'b111100100;
    x_193 = 'b111100100;
    x_194 = 'b111011111;
    x_195 = 'b111011101;
    x_196 = 'b111011011;
    x_197 = 'b111001111;
    x_198 = 'b111001111;
    x_199 = 'b111110101;
    x_200 = 'b111101000;
    x_201 = 'b111100010;
    x_202 = 'b111100010;
    x_203 = 'b111100000;
    x_204 = 'b111011110;
    x_205 = 'b111010001;
    x_206 = 'b111110110;
    x_207 = 'b111101110;
    x_208 = 'b111101001;
    x_209 = 'b111100101;
    x_210 = 'b111101010;
    x_211 = 'b111101101;
    x_212 = 'b111101010;
    x_213 = 'b111101010;
    x_214 = 'b111011111;
    x_215 = 'b111100110;
    x_216 = 'b111101011;
    x_217 = 'b111101011;
    x_218 = 'b111010110;
    x_219 = 'b111011011;
    x_220 = 'b111011110;
    x_221 = 'b111101000;
    x_222 = 'b111011010;
    x_223 = 'b111101000;
    x_224 = 'b111100000;
    x_225 = 'b111011000;
    x_226 = 'b111010011;
    x_227 = 'b111001101;
    x_228 = 'b111001111;
    x_229 = 'b111000100;
    x_230 = 'b111100011;
    x_231 = 'b111001100;
    x_232 = 'b111100100;
    x_233 = 'b111100110;
    x_234 = 'b111100001;
    x_235 = 'b111001010;
    x_236 = 'b111001111;
    x_237 = 'b111101001;
    x_238 = 'b111110010;
    x_239 = 'b111111000;
    x_240 = 'b111111001;
    x_241 = 'b000000100;
    x_242 = 'b111111001;
    x_243 = 'b111111111;
    x_244 = 'b000000000;
    x_245 = 'b111110111;
    x_246 = 'b111110101;
    x_247 = 'b111111110;
    x_248 = 'b000000110;
    x_249 = 'b000001011;
    x_250 = 'b000001111;
    x_251 = 'b000010000;
    x_252 = 'b111111010;
    x_253 = 'b111110111;
    x_254 = 'b000000001;
    x_255 = 'b111101101;

    h_0 = 'b111100100;
    h_1 = 'b111100100;
    h_2 = 'b111011111;
    h_3 = 'b111011101;
    h_4 = 'b111011011;
    h_5 = 'b111001111;
    h_6 = 'b111001111;
    h_7 = 'b111110101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111100010;
    x_1 = 'b111100001;
    x_2 = 'b111011011;
    x_3 = 'b111011101;
    x_4 = 'b111011011;
    x_5 = 'b111010011;
    x_6 = 'b111001110;
    x_7 = 'b111110001;
    x_8 = 'b111101000;
    x_9 = 'b111100111;
    x_10 = 'b111101101;
    x_11 = 'b111101111;
    x_12 = 'b111101010;
    x_13 = 'b111100010;
    x_14 = 'b111101110;
    x_15 = 'b111110001;
    x_16 = 'b111110001;
    x_17 = 'b111101111;
    x_18 = 'b111110101;
    x_19 = 'b111111010;
    x_20 = 'b111111000;
    x_21 = 'b111100111;
    x_22 = 'b111011011;
    x_23 = 'b111100011;
    x_24 = 'b111101000;
    x_25 = 'b111101001;
    x_26 = 'b111011000;
    x_27 = 'b111011011;
    x_28 = 'b111011001;
    x_29 = 'b111100111;
    x_30 = 'b111011010;
    x_31 = 'b111101111;
    x_32 = 'b111101000;
    x_33 = 'b111100010;
    x_34 = 'b111011100;
    x_35 = 'b111010110;
    x_36 = 'b111011000;
    x_37 = 'b111000110;
    x_38 = 'b111101010;
    x_39 = 'b111011011;
    x_40 = 'b111110011;
    x_41 = 'b111111110;
    x_42 = 'b111110101;
    x_43 = 'b110111011;
    x_44 = 'b111011011;
    x_45 = 'b111110001;
    x_46 = 'b000000000;
    x_47 = 'b000000101;
    x_48 = 'b000000111;
    x_49 = 'b000010101;
    x_50 = 'b000001001;
    x_51 = 'b000001011;
    x_52 = 'b000001010;
    x_53 = 'b000000011;
    x_54 = 'b000000100;
    x_55 = 'b000001111;
    x_56 = 'b000011000;
    x_57 = 'b000011011;
    x_58 = 'b000010111;
    x_59 = 'b000011100;
    x_60 = 'b000001010;
    x_61 = 'b000001000;
    x_62 = 'b000010001;
    x_63 = 'b000000011;
    x_64 = 'b111100010;
    x_65 = 'b111100001;
    x_66 = 'b111011011;
    x_67 = 'b111011101;
    x_68 = 'b111011011;
    x_69 = 'b111010011;
    x_70 = 'b111001110;
    x_71 = 'b111110001;
    x_72 = 'b111101000;
    x_73 = 'b111100111;
    x_74 = 'b111101101;
    x_75 = 'b111101111;
    x_76 = 'b111101010;
    x_77 = 'b111100010;
    x_78 = 'b111101110;
    x_79 = 'b111110001;
    x_80 = 'b111110001;
    x_81 = 'b111101111;
    x_82 = 'b111110101;
    x_83 = 'b111111010;
    x_84 = 'b111111000;
    x_85 = 'b111100111;
    x_86 = 'b111011011;
    x_87 = 'b111100011;
    x_88 = 'b111101000;
    x_89 = 'b111101001;
    x_90 = 'b111011000;
    x_91 = 'b111011011;
    x_92 = 'b111011001;
    x_93 = 'b111100111;
    x_94 = 'b111011010;
    x_95 = 'b111101111;
    x_96 = 'b111101000;
    x_97 = 'b111100010;
    x_98 = 'b111011100;
    x_99 = 'b111010110;
    x_100 = 'b111011000;
    x_101 = 'b111000110;
    x_102 = 'b111101010;
    x_103 = 'b111011011;
    x_104 = 'b111110011;
    x_105 = 'b111111110;
    x_106 = 'b111110101;
    x_107 = 'b110111011;
    x_108 = 'b111011011;
    x_109 = 'b111110001;
    x_110 = 'b000000000;
    x_111 = 'b000000101;
    x_112 = 'b000000111;
    x_113 = 'b000010101;
    x_114 = 'b000001001;
    x_115 = 'b000001011;
    x_116 = 'b000001010;
    x_117 = 'b000000011;
    x_118 = 'b000000100;
    x_119 = 'b000001111;
    x_120 = 'b000011000;
    x_121 = 'b000011011;
    x_122 = 'b000010111;
    x_123 = 'b000011100;
    x_124 = 'b000001010;
    x_125 = 'b000001000;
    x_126 = 'b000010001;
    x_127 = 'b000000011;
    x_128 = 'b111100010;
    x_129 = 'b111100001;
    x_130 = 'b111011011;
    x_131 = 'b111011101;
    x_132 = 'b111011011;
    x_133 = 'b111010011;
    x_134 = 'b111001110;
    x_135 = 'b111110001;
    x_136 = 'b111101000;
    x_137 = 'b111100111;
    x_138 = 'b111101101;
    x_139 = 'b111101111;
    x_140 = 'b111101010;
    x_141 = 'b111100010;
    x_142 = 'b111101110;
    x_143 = 'b111110001;
    x_144 = 'b111110001;
    x_145 = 'b111101111;
    x_146 = 'b111110101;
    x_147 = 'b111111010;
    x_148 = 'b111111000;
    x_149 = 'b111100111;
    x_150 = 'b111011011;
    x_151 = 'b111100011;
    x_152 = 'b111101000;
    x_153 = 'b111101001;
    x_154 = 'b111011000;
    x_155 = 'b111011011;
    x_156 = 'b111011001;
    x_157 = 'b111100111;
    x_158 = 'b111011010;
    x_159 = 'b111101111;
    x_160 = 'b111101000;
    x_161 = 'b111100010;
    x_162 = 'b111011100;
    x_163 = 'b111010110;
    x_164 = 'b111011000;
    x_165 = 'b111000110;
    x_166 = 'b111101010;
    x_167 = 'b111011011;
    x_168 = 'b111110011;
    x_169 = 'b111111110;
    x_170 = 'b111110101;
    x_171 = 'b110111011;
    x_172 = 'b111011011;
    x_173 = 'b111110001;
    x_174 = 'b000000000;
    x_175 = 'b000000101;
    x_176 = 'b000000111;
    x_177 = 'b000010101;
    x_178 = 'b000001001;
    x_179 = 'b000001011;
    x_180 = 'b000001010;
    x_181 = 'b000000011;
    x_182 = 'b000000100;
    x_183 = 'b000001111;
    x_184 = 'b000011000;
    x_185 = 'b000011011;
    x_186 = 'b000010111;
    x_187 = 'b000011100;
    x_188 = 'b000001010;
    x_189 = 'b000001000;
    x_190 = 'b000010001;
    x_191 = 'b000000011;
    x_192 = 'b111100010;
    x_193 = 'b111100001;
    x_194 = 'b111011011;
    x_195 = 'b111011101;
    x_196 = 'b111011011;
    x_197 = 'b111010011;
    x_198 = 'b111001110;
    x_199 = 'b111110001;
    x_200 = 'b111101000;
    x_201 = 'b111100111;
    x_202 = 'b111101101;
    x_203 = 'b111101111;
    x_204 = 'b111101010;
    x_205 = 'b111100010;
    x_206 = 'b111101110;
    x_207 = 'b111110001;
    x_208 = 'b111110001;
    x_209 = 'b111101111;
    x_210 = 'b111110101;
    x_211 = 'b111111010;
    x_212 = 'b111111000;
    x_213 = 'b111100111;
    x_214 = 'b111011011;
    x_215 = 'b111100011;
    x_216 = 'b111101000;
    x_217 = 'b111101001;
    x_218 = 'b111011000;
    x_219 = 'b111011011;
    x_220 = 'b111011001;
    x_221 = 'b111100111;
    x_222 = 'b111011010;
    x_223 = 'b111101111;
    x_224 = 'b111101000;
    x_225 = 'b111100010;
    x_226 = 'b111011100;
    x_227 = 'b111010110;
    x_228 = 'b111011000;
    x_229 = 'b111000110;
    x_230 = 'b111101010;
    x_231 = 'b111011011;
    x_232 = 'b111110011;
    x_233 = 'b111111110;
    x_234 = 'b111110101;
    x_235 = 'b110111011;
    x_236 = 'b111011011;
    x_237 = 'b111110001;
    x_238 = 'b000000000;
    x_239 = 'b000000101;
    x_240 = 'b000000111;
    x_241 = 'b000010101;
    x_242 = 'b000001001;
    x_243 = 'b000001011;
    x_244 = 'b000001010;
    x_245 = 'b000000011;
    x_246 = 'b000000100;
    x_247 = 'b000001111;
    x_248 = 'b000011000;
    x_249 = 'b000011011;
    x_250 = 'b000010111;
    x_251 = 'b000011100;
    x_252 = 'b000001010;
    x_253 = 'b000001000;
    x_254 = 'b000010001;
    x_255 = 'b000000011;

    h_0 = 'b111100010;
    h_1 = 'b111100001;
    h_2 = 'b111011011;
    h_3 = 'b111011101;
    h_4 = 'b111011011;
    h_5 = 'b111010011;
    h_6 = 'b111001110;
    h_7 = 'b111110001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111101101;
    x_1 = 'b111110101;
    x_2 = 'b111110011;
    x_3 = 'b111110100;
    x_4 = 'b111110011;
    x_5 = 'b111101100;
    x_6 = 'b111100111;
    x_7 = 'b000000101;
    x_8 = 'b111111110;
    x_9 = 'b111111110;
    x_10 = 'b000000100;
    x_11 = 'b000000110;
    x_12 = 'b111111111;
    x_13 = 'b111110011;
    x_14 = 'b000001000;
    x_15 = 'b000001000;
    x_16 = 'b000001000;
    x_17 = 'b000000101;
    x_18 = 'b000001010;
    x_19 = 'b000001100;
    x_20 = 'b000001001;
    x_21 = 'b111110011;
    x_22 = 'b111100111;
    x_23 = 'b111101100;
    x_24 = 'b111110011;
    x_25 = 'b111110100;
    x_26 = 'b111101100;
    x_27 = 'b111101101;
    x_28 = 'b111100110;
    x_29 = 'b111110010;
    x_30 = 'b111101000;
    x_31 = 'b000000010;
    x_32 = 'b111111111;
    x_33 = 'b111111000;
    x_34 = 'b111110000;
    x_35 = 'b111101110;
    x_36 = 'b111101111;
    x_37 = 'b111010011;
    x_38 = 'b111111111;
    x_39 = 'b111101000;
    x_40 = 'b000000110;
    x_41 = 'b111111100;
    x_42 = 'b000001010;
    x_43 = 'b111110110;
    x_44 = 'b111110010;
    x_45 = 'b111111101;
    x_46 = 'b000011000;
    x_47 = 'b000011101;
    x_48 = 'b000011100;
    x_49 = 'b000101001;
    x_50 = 'b000011111;
    x_51 = 'b000011011;
    x_52 = 'b000010111;
    x_53 = 'b000001110;
    x_54 = 'b000010011;
    x_55 = 'b000100100;
    x_56 = 'b000101100;
    x_57 = 'b000101111;
    x_58 = 'b000100010;
    x_59 = 'b000100011;
    x_60 = 'b000100011;
    x_61 = 'b000100001;
    x_62 = 'b000100001;
    x_63 = 'b000011110;
    x_64 = 'b111101101;
    x_65 = 'b111110101;
    x_66 = 'b111110011;
    x_67 = 'b111110100;
    x_68 = 'b111110011;
    x_69 = 'b111101100;
    x_70 = 'b111100111;
    x_71 = 'b000000101;
    x_72 = 'b111111110;
    x_73 = 'b111111110;
    x_74 = 'b000000100;
    x_75 = 'b000000110;
    x_76 = 'b111111111;
    x_77 = 'b111110011;
    x_78 = 'b000001000;
    x_79 = 'b000001000;
    x_80 = 'b000001000;
    x_81 = 'b000000101;
    x_82 = 'b000001010;
    x_83 = 'b000001100;
    x_84 = 'b000001001;
    x_85 = 'b111110011;
    x_86 = 'b111100111;
    x_87 = 'b111101100;
    x_88 = 'b111110011;
    x_89 = 'b111110100;
    x_90 = 'b111101100;
    x_91 = 'b111101101;
    x_92 = 'b111100110;
    x_93 = 'b111110010;
    x_94 = 'b111101000;
    x_95 = 'b000000010;
    x_96 = 'b111111111;
    x_97 = 'b111111000;
    x_98 = 'b111110000;
    x_99 = 'b111101110;
    x_100 = 'b111101111;
    x_101 = 'b111010011;
    x_102 = 'b111111111;
    x_103 = 'b111101000;
    x_104 = 'b000000110;
    x_105 = 'b111111100;
    x_106 = 'b000001010;
    x_107 = 'b111110110;
    x_108 = 'b111110010;
    x_109 = 'b111111101;
    x_110 = 'b000011000;
    x_111 = 'b000011101;
    x_112 = 'b000011100;
    x_113 = 'b000101001;
    x_114 = 'b000011111;
    x_115 = 'b000011011;
    x_116 = 'b000010111;
    x_117 = 'b000001110;
    x_118 = 'b000010011;
    x_119 = 'b000100100;
    x_120 = 'b000101100;
    x_121 = 'b000101111;
    x_122 = 'b000100010;
    x_123 = 'b000100011;
    x_124 = 'b000100011;
    x_125 = 'b000100001;
    x_126 = 'b000100001;
    x_127 = 'b000011110;
    x_128 = 'b111101101;
    x_129 = 'b111110101;
    x_130 = 'b111110011;
    x_131 = 'b111110100;
    x_132 = 'b111110011;
    x_133 = 'b111101100;
    x_134 = 'b111100111;
    x_135 = 'b000000101;
    x_136 = 'b111111110;
    x_137 = 'b111111110;
    x_138 = 'b000000100;
    x_139 = 'b000000110;
    x_140 = 'b111111111;
    x_141 = 'b111110011;
    x_142 = 'b000001000;
    x_143 = 'b000001000;
    x_144 = 'b000001000;
    x_145 = 'b000000101;
    x_146 = 'b000001010;
    x_147 = 'b000001100;
    x_148 = 'b000001001;
    x_149 = 'b111110011;
    x_150 = 'b111100111;
    x_151 = 'b111101100;
    x_152 = 'b111110011;
    x_153 = 'b111110100;
    x_154 = 'b111101100;
    x_155 = 'b111101101;
    x_156 = 'b111100110;
    x_157 = 'b111110010;
    x_158 = 'b111101000;
    x_159 = 'b000000010;
    x_160 = 'b111111111;
    x_161 = 'b111111000;
    x_162 = 'b111110000;
    x_163 = 'b111101110;
    x_164 = 'b111101111;
    x_165 = 'b111010011;
    x_166 = 'b111111111;
    x_167 = 'b111101000;
    x_168 = 'b000000110;
    x_169 = 'b111111100;
    x_170 = 'b000001010;
    x_171 = 'b111110110;
    x_172 = 'b111110010;
    x_173 = 'b111111101;
    x_174 = 'b000011000;
    x_175 = 'b000011101;
    x_176 = 'b000011100;
    x_177 = 'b000101001;
    x_178 = 'b000011111;
    x_179 = 'b000011011;
    x_180 = 'b000010111;
    x_181 = 'b000001110;
    x_182 = 'b000010011;
    x_183 = 'b000100100;
    x_184 = 'b000101100;
    x_185 = 'b000101111;
    x_186 = 'b000100010;
    x_187 = 'b000100011;
    x_188 = 'b000100011;
    x_189 = 'b000100001;
    x_190 = 'b000100001;
    x_191 = 'b000011110;
    x_192 = 'b111101101;
    x_193 = 'b111110101;
    x_194 = 'b111110011;
    x_195 = 'b111110100;
    x_196 = 'b111110011;
    x_197 = 'b111101100;
    x_198 = 'b111100111;
    x_199 = 'b000000101;
    x_200 = 'b111111110;
    x_201 = 'b111111110;
    x_202 = 'b000000100;
    x_203 = 'b000000110;
    x_204 = 'b111111111;
    x_205 = 'b111110011;
    x_206 = 'b000001000;
    x_207 = 'b000001000;
    x_208 = 'b000001000;
    x_209 = 'b000000101;
    x_210 = 'b000001010;
    x_211 = 'b000001100;
    x_212 = 'b000001001;
    x_213 = 'b111110011;
    x_214 = 'b111100111;
    x_215 = 'b111101100;
    x_216 = 'b111110011;
    x_217 = 'b111110100;
    x_218 = 'b111101100;
    x_219 = 'b111101101;
    x_220 = 'b111100110;
    x_221 = 'b111110010;
    x_222 = 'b111101000;
    x_223 = 'b000000010;
    x_224 = 'b111111111;
    x_225 = 'b111111000;
    x_226 = 'b111110000;
    x_227 = 'b111101110;
    x_228 = 'b111101111;
    x_229 = 'b111010011;
    x_230 = 'b111111111;
    x_231 = 'b111101000;
    x_232 = 'b000000110;
    x_233 = 'b111111100;
    x_234 = 'b000001010;
    x_235 = 'b111110110;
    x_236 = 'b111110010;
    x_237 = 'b111111101;
    x_238 = 'b000011000;
    x_239 = 'b000011101;
    x_240 = 'b000011100;
    x_241 = 'b000101001;
    x_242 = 'b000011111;
    x_243 = 'b000011011;
    x_244 = 'b000010111;
    x_245 = 'b000001110;
    x_246 = 'b000010011;
    x_247 = 'b000100100;
    x_248 = 'b000101100;
    x_249 = 'b000101111;
    x_250 = 'b000100010;
    x_251 = 'b000100011;
    x_252 = 'b000100011;
    x_253 = 'b000100001;
    x_254 = 'b000100001;
    x_255 = 'b000011110;

    h_0 = 'b111101101;
    h_1 = 'b111110101;
    h_2 = 'b111110011;
    h_3 = 'b111110100;
    h_4 = 'b111110011;
    h_5 = 'b111101100;
    h_6 = 'b111100111;
    h_7 = 'b000000101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111111100;
    x_1 = 'b000000110;
    x_2 = 'b111111111;
    x_3 = 'b111111100;
    x_4 = 'b111111000;
    x_5 = 'b111110001;
    x_6 = 'b111101111;
    x_7 = 'b000011000;
    x_8 = 'b000001011;
    x_9 = 'b000001000;
    x_10 = 'b000001010;
    x_11 = 'b000000010;
    x_12 = 'b111111101;
    x_13 = 'b111100111;
    x_14 = 'b000010111;
    x_15 = 'b000010011;
    x_16 = 'b000010000;
    x_17 = 'b000001011;
    x_18 = 'b000001101;
    x_19 = 'b000001010;
    x_20 = 'b000000001;
    x_21 = 'b111110011;
    x_22 = 'b111101011;
    x_23 = 'b111101110;
    x_24 = 'b111110100;
    x_25 = 'b111110110;
    x_26 = 'b111101101;
    x_27 = 'b111110000;
    x_28 = 'b111101010;
    x_29 = 'b111111111;
    x_30 = 'b111100001;
    x_31 = 'b000000100;
    x_32 = 'b111111110;
    x_33 = 'b111110100;
    x_34 = 'b111101101;
    x_35 = 'b111101011;
    x_36 = 'b111110000;
    x_37 = 'b111010100;
    x_38 = 'b000000100;
    x_39 = 'b111100011;
    x_40 = 'b000001110;
    x_41 = 'b111101010;
    x_42 = 'b000000111;
    x_43 = 'b111100011;
    x_44 = 'b111110111;
    x_45 = 'b111110101;
    x_46 = 'b000011111;
    x_47 = 'b000100010;
    x_48 = 'b000100010;
    x_49 = 'b000101010;
    x_50 = 'b000100000;
    x_51 = 'b000011010;
    x_52 = 'b000010100;
    x_53 = 'b000000111;
    x_54 = 'b000000100;
    x_55 = 'b000101100;
    x_56 = 'b000110010;
    x_57 = 'b000110110;
    x_58 = 'b000100000;
    x_59 = 'b000011011;
    x_60 = 'b000110111;
    x_61 = 'b000110001;
    x_62 = 'b000100111;
    x_63 = 'b000101100;
    x_64 = 'b111111100;
    x_65 = 'b000000110;
    x_66 = 'b111111111;
    x_67 = 'b111111100;
    x_68 = 'b111111000;
    x_69 = 'b111110001;
    x_70 = 'b111101111;
    x_71 = 'b000011000;
    x_72 = 'b000001011;
    x_73 = 'b000001000;
    x_74 = 'b000001010;
    x_75 = 'b000000010;
    x_76 = 'b111111101;
    x_77 = 'b111100111;
    x_78 = 'b000010111;
    x_79 = 'b000010011;
    x_80 = 'b000010000;
    x_81 = 'b000001011;
    x_82 = 'b000001101;
    x_83 = 'b000001010;
    x_84 = 'b000000001;
    x_85 = 'b111110011;
    x_86 = 'b111101011;
    x_87 = 'b111101110;
    x_88 = 'b111110100;
    x_89 = 'b111110110;
    x_90 = 'b111101101;
    x_91 = 'b111110000;
    x_92 = 'b111101010;
    x_93 = 'b111111111;
    x_94 = 'b111100001;
    x_95 = 'b000000100;
    x_96 = 'b111111110;
    x_97 = 'b111110100;
    x_98 = 'b111101101;
    x_99 = 'b111101011;
    x_100 = 'b111110000;
    x_101 = 'b111010100;
    x_102 = 'b000000100;
    x_103 = 'b111100011;
    x_104 = 'b000001110;
    x_105 = 'b111101010;
    x_106 = 'b000000111;
    x_107 = 'b111100011;
    x_108 = 'b111110111;
    x_109 = 'b111110101;
    x_110 = 'b000011111;
    x_111 = 'b000100010;
    x_112 = 'b000100010;
    x_113 = 'b000101010;
    x_114 = 'b000100000;
    x_115 = 'b000011010;
    x_116 = 'b000010100;
    x_117 = 'b000000111;
    x_118 = 'b000000100;
    x_119 = 'b000101100;
    x_120 = 'b000110010;
    x_121 = 'b000110110;
    x_122 = 'b000100000;
    x_123 = 'b000011011;
    x_124 = 'b000110111;
    x_125 = 'b000110001;
    x_126 = 'b000100111;
    x_127 = 'b000101100;
    x_128 = 'b111111100;
    x_129 = 'b000000110;
    x_130 = 'b111111111;
    x_131 = 'b111111100;
    x_132 = 'b111111000;
    x_133 = 'b111110001;
    x_134 = 'b111101111;
    x_135 = 'b000011000;
    x_136 = 'b000001011;
    x_137 = 'b000001000;
    x_138 = 'b000001010;
    x_139 = 'b000000010;
    x_140 = 'b111111101;
    x_141 = 'b111100111;
    x_142 = 'b000010111;
    x_143 = 'b000010011;
    x_144 = 'b000010000;
    x_145 = 'b000001011;
    x_146 = 'b000001101;
    x_147 = 'b000001010;
    x_148 = 'b000000001;
    x_149 = 'b111110011;
    x_150 = 'b111101011;
    x_151 = 'b111101110;
    x_152 = 'b111110100;
    x_153 = 'b111110110;
    x_154 = 'b111101101;
    x_155 = 'b111110000;
    x_156 = 'b111101010;
    x_157 = 'b111111111;
    x_158 = 'b111100001;
    x_159 = 'b000000100;
    x_160 = 'b111111110;
    x_161 = 'b111110100;
    x_162 = 'b111101101;
    x_163 = 'b111101011;
    x_164 = 'b111110000;
    x_165 = 'b111010100;
    x_166 = 'b000000100;
    x_167 = 'b111100011;
    x_168 = 'b000001110;
    x_169 = 'b111101010;
    x_170 = 'b000000111;
    x_171 = 'b111100011;
    x_172 = 'b111110111;
    x_173 = 'b111110101;
    x_174 = 'b000011111;
    x_175 = 'b000100010;
    x_176 = 'b000100010;
    x_177 = 'b000101010;
    x_178 = 'b000100000;
    x_179 = 'b000011010;
    x_180 = 'b000010100;
    x_181 = 'b000000111;
    x_182 = 'b000000100;
    x_183 = 'b000101100;
    x_184 = 'b000110010;
    x_185 = 'b000110110;
    x_186 = 'b000100000;
    x_187 = 'b000011011;
    x_188 = 'b000110111;
    x_189 = 'b000110001;
    x_190 = 'b000100111;
    x_191 = 'b000101100;
    x_192 = 'b111111100;
    x_193 = 'b000000110;
    x_194 = 'b111111111;
    x_195 = 'b111111100;
    x_196 = 'b111111000;
    x_197 = 'b111110001;
    x_198 = 'b111101111;
    x_199 = 'b000011000;
    x_200 = 'b000001011;
    x_201 = 'b000001000;
    x_202 = 'b000001010;
    x_203 = 'b000000010;
    x_204 = 'b111111101;
    x_205 = 'b111100111;
    x_206 = 'b000010111;
    x_207 = 'b000010011;
    x_208 = 'b000010000;
    x_209 = 'b000001011;
    x_210 = 'b000001101;
    x_211 = 'b000001010;
    x_212 = 'b000000001;
    x_213 = 'b111110011;
    x_214 = 'b111101011;
    x_215 = 'b111101110;
    x_216 = 'b111110100;
    x_217 = 'b111110110;
    x_218 = 'b111101101;
    x_219 = 'b111110000;
    x_220 = 'b111101010;
    x_221 = 'b111111111;
    x_222 = 'b111100001;
    x_223 = 'b000000100;
    x_224 = 'b111111110;
    x_225 = 'b111110100;
    x_226 = 'b111101101;
    x_227 = 'b111101011;
    x_228 = 'b111110000;
    x_229 = 'b111010100;
    x_230 = 'b000000100;
    x_231 = 'b111100011;
    x_232 = 'b000001110;
    x_233 = 'b111101010;
    x_234 = 'b000000111;
    x_235 = 'b111100011;
    x_236 = 'b111110111;
    x_237 = 'b111110101;
    x_238 = 'b000011111;
    x_239 = 'b000100010;
    x_240 = 'b000100010;
    x_241 = 'b000101010;
    x_242 = 'b000100000;
    x_243 = 'b000011010;
    x_244 = 'b000010100;
    x_245 = 'b000000111;
    x_246 = 'b000000100;
    x_247 = 'b000101100;
    x_248 = 'b000110010;
    x_249 = 'b000110110;
    x_250 = 'b000100000;
    x_251 = 'b000011011;
    x_252 = 'b000110111;
    x_253 = 'b000110001;
    x_254 = 'b000100111;
    x_255 = 'b000101100;

    h_0 = 'b111111100;
    h_1 = 'b000000110;
    h_2 = 'b111111111;
    h_3 = 'b111111100;
    h_4 = 'b111111000;
    h_5 = 'b111110001;
    h_6 = 'b111101111;
    h_7 = 'b000011000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000000010;
    x_1 = 'b000000010;
    x_2 = 'b111111001;
    x_3 = 'b111110010;
    x_4 = 'b111101110;
    x_5 = 'b111101000;
    x_6 = 'b111101001;
    x_7 = 'b000011001;
    x_8 = 'b000001010;
    x_9 = 'b000000011;
    x_10 = 'b111111111;
    x_11 = 'b111110011;
    x_12 = 'b111110011;
    x_13 = 'b111100011;
    x_14 = 'b000011100;
    x_15 = 'b000010101;
    x_16 = 'b000001110;
    x_17 = 'b000001000;
    x_18 = 'b000001000;
    x_19 = 'b000000100;
    x_20 = 'b111111111;
    x_21 = 'b111110101;
    x_22 = 'b111101101;
    x_23 = 'b111110001;
    x_24 = 'b111111000;
    x_25 = 'b111111010;
    x_26 = 'b111101101;
    x_27 = 'b111110010;
    x_28 = 'b111101110;
    x_29 = 'b000000111;
    x_30 = 'b111101101;
    x_31 = 'b000000100;
    x_32 = 'b000000000;
    x_33 = 'b111110111;
    x_34 = 'b111101111;
    x_35 = 'b111101110;
    x_36 = 'b111110001;
    x_37 = 'b111010110;
    x_38 = 'b000011000;
    x_39 = 'b111101100;
    x_40 = 'b000011101;
    x_41 = 'b000000110;
    x_42 = 'b000011000;
    x_43 = 'b111010100;
    x_44 = 'b000000001;
    x_45 = 'b111110100;
    x_46 = 'b000101110;
    x_47 = 'b000101110;
    x_48 = 'b000101100;
    x_49 = 'b000110011;
    x_50 = 'b000100101;
    x_51 = 'b000011110;
    x_52 = 'b000011001;
    x_53 = 'b000001011;
    x_54 = 'b000000100;
    x_55 = 'b000111001;
    x_56 = 'b000111100;
    x_57 = 'b000111110;
    x_58 = 'b000100011;
    x_59 = 'b000011110;
    x_60 = 'b001000011;
    x_61 = 'b000111001;
    x_62 = 'b000100110;
    x_63 = 'b000101110;
    x_64 = 'b000000010;
    x_65 = 'b000000010;
    x_66 = 'b111111001;
    x_67 = 'b111110010;
    x_68 = 'b111101110;
    x_69 = 'b111101000;
    x_70 = 'b111101001;
    x_71 = 'b000011001;
    x_72 = 'b000001010;
    x_73 = 'b000000011;
    x_74 = 'b111111111;
    x_75 = 'b111110011;
    x_76 = 'b111110011;
    x_77 = 'b111100011;
    x_78 = 'b000011100;
    x_79 = 'b000010101;
    x_80 = 'b000001110;
    x_81 = 'b000001000;
    x_82 = 'b000001000;
    x_83 = 'b000000100;
    x_84 = 'b111111111;
    x_85 = 'b111110101;
    x_86 = 'b111101101;
    x_87 = 'b111110001;
    x_88 = 'b111111000;
    x_89 = 'b111111010;
    x_90 = 'b111101101;
    x_91 = 'b111110010;
    x_92 = 'b111101110;
    x_93 = 'b000000111;
    x_94 = 'b111101101;
    x_95 = 'b000000100;
    x_96 = 'b000000000;
    x_97 = 'b111110111;
    x_98 = 'b111101111;
    x_99 = 'b111101110;
    x_100 = 'b111110001;
    x_101 = 'b111010110;
    x_102 = 'b000011000;
    x_103 = 'b111101100;
    x_104 = 'b000011101;
    x_105 = 'b000000110;
    x_106 = 'b000011000;
    x_107 = 'b111010100;
    x_108 = 'b000000001;
    x_109 = 'b111110100;
    x_110 = 'b000101110;
    x_111 = 'b000101110;
    x_112 = 'b000101100;
    x_113 = 'b000110011;
    x_114 = 'b000100101;
    x_115 = 'b000011110;
    x_116 = 'b000011001;
    x_117 = 'b000001011;
    x_118 = 'b000000100;
    x_119 = 'b000111001;
    x_120 = 'b000111100;
    x_121 = 'b000111110;
    x_122 = 'b000100011;
    x_123 = 'b000011110;
    x_124 = 'b001000011;
    x_125 = 'b000111001;
    x_126 = 'b000100110;
    x_127 = 'b000101110;
    x_128 = 'b000000010;
    x_129 = 'b000000010;
    x_130 = 'b111111001;
    x_131 = 'b111110010;
    x_132 = 'b111101110;
    x_133 = 'b111101000;
    x_134 = 'b111101001;
    x_135 = 'b000011001;
    x_136 = 'b000001010;
    x_137 = 'b000000011;
    x_138 = 'b111111111;
    x_139 = 'b111110011;
    x_140 = 'b111110011;
    x_141 = 'b111100011;
    x_142 = 'b000011100;
    x_143 = 'b000010101;
    x_144 = 'b000001110;
    x_145 = 'b000001000;
    x_146 = 'b000001000;
    x_147 = 'b000000100;
    x_148 = 'b111111111;
    x_149 = 'b111110101;
    x_150 = 'b111101101;
    x_151 = 'b111110001;
    x_152 = 'b111111000;
    x_153 = 'b111111010;
    x_154 = 'b111101101;
    x_155 = 'b111110010;
    x_156 = 'b111101110;
    x_157 = 'b000000111;
    x_158 = 'b111101101;
    x_159 = 'b000000100;
    x_160 = 'b000000000;
    x_161 = 'b111110111;
    x_162 = 'b111101111;
    x_163 = 'b111101110;
    x_164 = 'b111110001;
    x_165 = 'b111010110;
    x_166 = 'b000011000;
    x_167 = 'b111101100;
    x_168 = 'b000011101;
    x_169 = 'b000000110;
    x_170 = 'b000011000;
    x_171 = 'b111010100;
    x_172 = 'b000000001;
    x_173 = 'b111110100;
    x_174 = 'b000101110;
    x_175 = 'b000101110;
    x_176 = 'b000101100;
    x_177 = 'b000110011;
    x_178 = 'b000100101;
    x_179 = 'b000011110;
    x_180 = 'b000011001;
    x_181 = 'b000001011;
    x_182 = 'b000000100;
    x_183 = 'b000111001;
    x_184 = 'b000111100;
    x_185 = 'b000111110;
    x_186 = 'b000100011;
    x_187 = 'b000011110;
    x_188 = 'b001000011;
    x_189 = 'b000111001;
    x_190 = 'b000100110;
    x_191 = 'b000101110;
    x_192 = 'b000000010;
    x_193 = 'b000000010;
    x_194 = 'b111111001;
    x_195 = 'b111110010;
    x_196 = 'b111101110;
    x_197 = 'b111101000;
    x_198 = 'b111101001;
    x_199 = 'b000011001;
    x_200 = 'b000001010;
    x_201 = 'b000000011;
    x_202 = 'b111111111;
    x_203 = 'b111110011;
    x_204 = 'b111110011;
    x_205 = 'b111100011;
    x_206 = 'b000011100;
    x_207 = 'b000010101;
    x_208 = 'b000001110;
    x_209 = 'b000001000;
    x_210 = 'b000001000;
    x_211 = 'b000000100;
    x_212 = 'b111111111;
    x_213 = 'b111110101;
    x_214 = 'b111101101;
    x_215 = 'b111110001;
    x_216 = 'b111111000;
    x_217 = 'b111111010;
    x_218 = 'b111101101;
    x_219 = 'b111110010;
    x_220 = 'b111101110;
    x_221 = 'b000000111;
    x_222 = 'b111101101;
    x_223 = 'b000000100;
    x_224 = 'b000000000;
    x_225 = 'b111110111;
    x_226 = 'b111101111;
    x_227 = 'b111101110;
    x_228 = 'b111110001;
    x_229 = 'b111010110;
    x_230 = 'b000011000;
    x_231 = 'b111101100;
    x_232 = 'b000011101;
    x_233 = 'b000000110;
    x_234 = 'b000011000;
    x_235 = 'b111010100;
    x_236 = 'b000000001;
    x_237 = 'b111110100;
    x_238 = 'b000101110;
    x_239 = 'b000101110;
    x_240 = 'b000101100;
    x_241 = 'b000110011;
    x_242 = 'b000100101;
    x_243 = 'b000011110;
    x_244 = 'b000011001;
    x_245 = 'b000001011;
    x_246 = 'b000000100;
    x_247 = 'b000111001;
    x_248 = 'b000111100;
    x_249 = 'b000111110;
    x_250 = 'b000100011;
    x_251 = 'b000011110;
    x_252 = 'b001000011;
    x_253 = 'b000111001;
    x_254 = 'b000100110;
    x_255 = 'b000101110;

    h_0 = 'b000000010;
    h_1 = 'b000000010;
    h_2 = 'b111111001;
    h_3 = 'b111110010;
    h_4 = 'b111101110;
    h_5 = 'b111101000;
    h_6 = 'b111101001;
    h_7 = 'b000011001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000010011;
    x_1 = 'b000010010;
    x_2 = 'b000000110;
    x_3 = 'b111111101;
    x_4 = 'b111111000;
    x_5 = 'b111101111;
    x_6 = 'b111101110;
    x_7 = 'b000101101;
    x_8 = 'b000011101;
    x_9 = 'b000010011;
    x_10 = 'b000001011;
    x_11 = 'b111111101;
    x_12 = 'b111111011;
    x_13 = 'b111101110;
    x_14 = 'b000110000;
    x_15 = 'b000101000;
    x_16 = 'b000011101;
    x_17 = 'b000010100;
    x_18 = 'b000010010;
    x_19 = 'b000001110;
    x_20 = 'b000001001;
    x_21 = 'b111111100;
    x_22 = 'b111110001;
    x_23 = 'b111110100;
    x_24 = 'b111111110;
    x_25 = 'b111111111;
    x_26 = 'b111110011;
    x_27 = 'b111110101;
    x_28 = 'b111101101;
    x_29 = 'b000001101;
    x_30 = 'b111111001;
    x_31 = 'b000001001;
    x_32 = 'b000001000;
    x_33 = 'b111111110;
    x_34 = 'b111110110;
    x_35 = 'b111110011;
    x_36 = 'b111101101;
    x_37 = 'b111010001;
    x_38 = 'b000011100;
    x_39 = 'b111100101;
    x_40 = 'b000011100;
    x_41 = 'b111110011;
    x_42 = 'b000001110;
    x_43 = 'b111011011;
    x_44 = 'b000001111;
    x_45 = 'b111111000;
    x_46 = 'b000110110;
    x_47 = 'b000110111;
    x_48 = 'b000110101;
    x_49 = 'b000111100;
    x_50 = 'b000101101;
    x_51 = 'b000100101;
    x_52 = 'b000100000;
    x_53 = 'b000010011;
    x_54 = 'b000001101;
    x_55 = 'b000111101;
    x_56 = 'b001000000;
    x_57 = 'b001000001;
    x_58 = 'b000101000;
    x_59 = 'b000100101;
    x_60 = 'b001001000;
    x_61 = 'b000111110;
    x_62 = 'b000101001;
    x_63 = 'b000110011;
    x_64 = 'b000010011;
    x_65 = 'b000010010;
    x_66 = 'b000000110;
    x_67 = 'b111111101;
    x_68 = 'b111111000;
    x_69 = 'b111101111;
    x_70 = 'b111101110;
    x_71 = 'b000101101;
    x_72 = 'b000011101;
    x_73 = 'b000010011;
    x_74 = 'b000001011;
    x_75 = 'b111111101;
    x_76 = 'b111111011;
    x_77 = 'b111101110;
    x_78 = 'b000110000;
    x_79 = 'b000101000;
    x_80 = 'b000011101;
    x_81 = 'b000010100;
    x_82 = 'b000010010;
    x_83 = 'b000001110;
    x_84 = 'b000001001;
    x_85 = 'b111111100;
    x_86 = 'b111110001;
    x_87 = 'b111110100;
    x_88 = 'b111111110;
    x_89 = 'b111111111;
    x_90 = 'b111110011;
    x_91 = 'b111110101;
    x_92 = 'b111101101;
    x_93 = 'b000001101;
    x_94 = 'b111111001;
    x_95 = 'b000001001;
    x_96 = 'b000001000;
    x_97 = 'b111111110;
    x_98 = 'b111110110;
    x_99 = 'b111110011;
    x_100 = 'b111101101;
    x_101 = 'b111010001;
    x_102 = 'b000011100;
    x_103 = 'b111100101;
    x_104 = 'b000011100;
    x_105 = 'b111110011;
    x_106 = 'b000001110;
    x_107 = 'b111011011;
    x_108 = 'b000001111;
    x_109 = 'b111111000;
    x_110 = 'b000110110;
    x_111 = 'b000110111;
    x_112 = 'b000110101;
    x_113 = 'b000111100;
    x_114 = 'b000101101;
    x_115 = 'b000100101;
    x_116 = 'b000100000;
    x_117 = 'b000010011;
    x_118 = 'b000001101;
    x_119 = 'b000111101;
    x_120 = 'b001000000;
    x_121 = 'b001000001;
    x_122 = 'b000101000;
    x_123 = 'b000100101;
    x_124 = 'b001001000;
    x_125 = 'b000111110;
    x_126 = 'b000101001;
    x_127 = 'b000110011;
    x_128 = 'b000010011;
    x_129 = 'b000010010;
    x_130 = 'b000000110;
    x_131 = 'b111111101;
    x_132 = 'b111111000;
    x_133 = 'b111101111;
    x_134 = 'b111101110;
    x_135 = 'b000101101;
    x_136 = 'b000011101;
    x_137 = 'b000010011;
    x_138 = 'b000001011;
    x_139 = 'b111111101;
    x_140 = 'b111111011;
    x_141 = 'b111101110;
    x_142 = 'b000110000;
    x_143 = 'b000101000;
    x_144 = 'b000011101;
    x_145 = 'b000010100;
    x_146 = 'b000010010;
    x_147 = 'b000001110;
    x_148 = 'b000001001;
    x_149 = 'b111111100;
    x_150 = 'b111110001;
    x_151 = 'b111110100;
    x_152 = 'b111111110;
    x_153 = 'b111111111;
    x_154 = 'b111110011;
    x_155 = 'b111110101;
    x_156 = 'b111101101;
    x_157 = 'b000001101;
    x_158 = 'b111111001;
    x_159 = 'b000001001;
    x_160 = 'b000001000;
    x_161 = 'b111111110;
    x_162 = 'b111110110;
    x_163 = 'b111110011;
    x_164 = 'b111101101;
    x_165 = 'b111010001;
    x_166 = 'b000011100;
    x_167 = 'b111100101;
    x_168 = 'b000011100;
    x_169 = 'b111110011;
    x_170 = 'b000001110;
    x_171 = 'b111011011;
    x_172 = 'b000001111;
    x_173 = 'b111111000;
    x_174 = 'b000110110;
    x_175 = 'b000110111;
    x_176 = 'b000110101;
    x_177 = 'b000111100;
    x_178 = 'b000101101;
    x_179 = 'b000100101;
    x_180 = 'b000100000;
    x_181 = 'b000010011;
    x_182 = 'b000001101;
    x_183 = 'b000111101;
    x_184 = 'b001000000;
    x_185 = 'b001000001;
    x_186 = 'b000101000;
    x_187 = 'b000100101;
    x_188 = 'b001001000;
    x_189 = 'b000111110;
    x_190 = 'b000101001;
    x_191 = 'b000110011;
    x_192 = 'b000010011;
    x_193 = 'b000010010;
    x_194 = 'b000000110;
    x_195 = 'b111111101;
    x_196 = 'b111111000;
    x_197 = 'b111101111;
    x_198 = 'b111101110;
    x_199 = 'b000101101;
    x_200 = 'b000011101;
    x_201 = 'b000010011;
    x_202 = 'b000001011;
    x_203 = 'b111111101;
    x_204 = 'b111111011;
    x_205 = 'b111101110;
    x_206 = 'b000110000;
    x_207 = 'b000101000;
    x_208 = 'b000011101;
    x_209 = 'b000010100;
    x_210 = 'b000010010;
    x_211 = 'b000001110;
    x_212 = 'b000001001;
    x_213 = 'b111111100;
    x_214 = 'b111110001;
    x_215 = 'b111110100;
    x_216 = 'b111111110;
    x_217 = 'b111111111;
    x_218 = 'b111110011;
    x_219 = 'b111110101;
    x_220 = 'b111101101;
    x_221 = 'b000001101;
    x_222 = 'b111111001;
    x_223 = 'b000001001;
    x_224 = 'b000001000;
    x_225 = 'b111111110;
    x_226 = 'b111110110;
    x_227 = 'b111110011;
    x_228 = 'b111101101;
    x_229 = 'b111010001;
    x_230 = 'b000011100;
    x_231 = 'b111100101;
    x_232 = 'b000011100;
    x_233 = 'b111110011;
    x_234 = 'b000001110;
    x_235 = 'b111011011;
    x_236 = 'b000001111;
    x_237 = 'b111111000;
    x_238 = 'b000110110;
    x_239 = 'b000110111;
    x_240 = 'b000110101;
    x_241 = 'b000111100;
    x_242 = 'b000101101;
    x_243 = 'b000100101;
    x_244 = 'b000100000;
    x_245 = 'b000010011;
    x_246 = 'b000001101;
    x_247 = 'b000111101;
    x_248 = 'b001000000;
    x_249 = 'b001000001;
    x_250 = 'b000101000;
    x_251 = 'b000100101;
    x_252 = 'b001001000;
    x_253 = 'b000111110;
    x_254 = 'b000101001;
    x_255 = 'b000110011;

    h_0 = 'b000010011;
    h_1 = 'b000010010;
    h_2 = 'b000000110;
    h_3 = 'b111111101;
    h_4 = 'b111111000;
    h_5 = 'b111101111;
    h_6 = 'b111101110;
    h_7 = 'b000101101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000001111;
    x_1 = 'b000010011;
    x_2 = 'b000000110;
    x_3 = 'b000000001;
    x_4 = 'b111111011;
    x_5 = 'b111110000;
    x_6 = 'b111110000;
    x_7 = 'b000101001;
    x_8 = 'b000100000;
    x_9 = 'b000010110;
    x_10 = 'b000010100;
    x_11 = 'b000000110;
    x_12 = 'b000000011;
    x_13 = 'b111110011;
    x_14 = 'b000101011;
    x_15 = 'b000101010;
    x_16 = 'b000100011;
    x_17 = 'b000011001;
    x_18 = 'b000010111;
    x_19 = 'b000010010;
    x_20 = 'b000001100;
    x_21 = 'b111110111;
    x_22 = 'b111101011;
    x_23 = 'b111101110;
    x_24 = 'b111110111;
    x_25 = 'b111111001;
    x_26 = 'b111101010;
    x_27 = 'b111101101;
    x_28 = 'b111100110;
    x_29 = 'b000000011;
    x_30 = 'b111110011;
    x_31 = 'b000000010;
    x_32 = 'b111111101;
    x_33 = 'b111110011;
    x_34 = 'b111101101;
    x_35 = 'b111100111;
    x_36 = 'b111100110;
    x_37 = 'b111001110;
    x_38 = 'b000001111;
    x_39 = 'b111100000;
    x_40 = 'b000001100;
    x_41 = 'b111110101;
    x_42 = 'b000010100;
    x_43 = 'b111000110;
    x_44 = 'b000001110;
    x_45 = 'b111110001;
    x_46 = 'b000101000;
    x_47 = 'b000101110;
    x_48 = 'b000101111;
    x_49 = 'b000111000;
    x_50 = 'b000101001;
    x_51 = 'b000011111;
    x_52 = 'b000011010;
    x_53 = 'b000001100;
    x_54 = 'b000001100;
    x_55 = 'b000110111;
    x_56 = 'b000111011;
    x_57 = 'b000111011;
    x_58 = 'b000100010;
    x_59 = 'b000011111;
    x_60 = 'b001001000;
    x_61 = 'b000111111;
    x_62 = 'b000101111;
    x_63 = 'b000111010;
    x_64 = 'b000001111;
    x_65 = 'b000010011;
    x_66 = 'b000000110;
    x_67 = 'b000000001;
    x_68 = 'b111111011;
    x_69 = 'b111110000;
    x_70 = 'b111110000;
    x_71 = 'b000101001;
    x_72 = 'b000100000;
    x_73 = 'b000010110;
    x_74 = 'b000010100;
    x_75 = 'b000000110;
    x_76 = 'b000000011;
    x_77 = 'b111110011;
    x_78 = 'b000101011;
    x_79 = 'b000101010;
    x_80 = 'b000100011;
    x_81 = 'b000011001;
    x_82 = 'b000010111;
    x_83 = 'b000010010;
    x_84 = 'b000001100;
    x_85 = 'b111110111;
    x_86 = 'b111101011;
    x_87 = 'b111101110;
    x_88 = 'b111110111;
    x_89 = 'b111111001;
    x_90 = 'b111101010;
    x_91 = 'b111101101;
    x_92 = 'b111100110;
    x_93 = 'b000000011;
    x_94 = 'b111110011;
    x_95 = 'b000000010;
    x_96 = 'b111111101;
    x_97 = 'b111110011;
    x_98 = 'b111101101;
    x_99 = 'b111100111;
    x_100 = 'b111100110;
    x_101 = 'b111001110;
    x_102 = 'b000001111;
    x_103 = 'b111100000;
    x_104 = 'b000001100;
    x_105 = 'b111110101;
    x_106 = 'b000010100;
    x_107 = 'b111000110;
    x_108 = 'b000001110;
    x_109 = 'b111110001;
    x_110 = 'b000101000;
    x_111 = 'b000101110;
    x_112 = 'b000101111;
    x_113 = 'b000111000;
    x_114 = 'b000101001;
    x_115 = 'b000011111;
    x_116 = 'b000011010;
    x_117 = 'b000001100;
    x_118 = 'b000001100;
    x_119 = 'b000110111;
    x_120 = 'b000111011;
    x_121 = 'b000111011;
    x_122 = 'b000100010;
    x_123 = 'b000011111;
    x_124 = 'b001001000;
    x_125 = 'b000111111;
    x_126 = 'b000101111;
    x_127 = 'b000111010;
    x_128 = 'b000001111;
    x_129 = 'b000010011;
    x_130 = 'b000000110;
    x_131 = 'b000000001;
    x_132 = 'b111111011;
    x_133 = 'b111110000;
    x_134 = 'b111110000;
    x_135 = 'b000101001;
    x_136 = 'b000100000;
    x_137 = 'b000010110;
    x_138 = 'b000010100;
    x_139 = 'b000000110;
    x_140 = 'b000000011;
    x_141 = 'b111110011;
    x_142 = 'b000101011;
    x_143 = 'b000101010;
    x_144 = 'b000100011;
    x_145 = 'b000011001;
    x_146 = 'b000010111;
    x_147 = 'b000010010;
    x_148 = 'b000001100;
    x_149 = 'b111110111;
    x_150 = 'b111101011;
    x_151 = 'b111101110;
    x_152 = 'b111110111;
    x_153 = 'b111111001;
    x_154 = 'b111101010;
    x_155 = 'b111101101;
    x_156 = 'b111100110;
    x_157 = 'b000000011;
    x_158 = 'b111110011;
    x_159 = 'b000000010;
    x_160 = 'b111111101;
    x_161 = 'b111110011;
    x_162 = 'b111101101;
    x_163 = 'b111100111;
    x_164 = 'b111100110;
    x_165 = 'b111001110;
    x_166 = 'b000001111;
    x_167 = 'b111100000;
    x_168 = 'b000001100;
    x_169 = 'b111110101;
    x_170 = 'b000010100;
    x_171 = 'b111000110;
    x_172 = 'b000001110;
    x_173 = 'b111110001;
    x_174 = 'b000101000;
    x_175 = 'b000101110;
    x_176 = 'b000101111;
    x_177 = 'b000111000;
    x_178 = 'b000101001;
    x_179 = 'b000011111;
    x_180 = 'b000011010;
    x_181 = 'b000001100;
    x_182 = 'b000001100;
    x_183 = 'b000110111;
    x_184 = 'b000111011;
    x_185 = 'b000111011;
    x_186 = 'b000100010;
    x_187 = 'b000011111;
    x_188 = 'b001001000;
    x_189 = 'b000111111;
    x_190 = 'b000101111;
    x_191 = 'b000111010;
    x_192 = 'b000001111;
    x_193 = 'b000010011;
    x_194 = 'b000000110;
    x_195 = 'b000000001;
    x_196 = 'b111111011;
    x_197 = 'b111110000;
    x_198 = 'b111110000;
    x_199 = 'b000101001;
    x_200 = 'b000100000;
    x_201 = 'b000010110;
    x_202 = 'b000010100;
    x_203 = 'b000000110;
    x_204 = 'b000000011;
    x_205 = 'b111110011;
    x_206 = 'b000101011;
    x_207 = 'b000101010;
    x_208 = 'b000100011;
    x_209 = 'b000011001;
    x_210 = 'b000010111;
    x_211 = 'b000010010;
    x_212 = 'b000001100;
    x_213 = 'b111110111;
    x_214 = 'b111101011;
    x_215 = 'b111101110;
    x_216 = 'b111110111;
    x_217 = 'b111111001;
    x_218 = 'b111101010;
    x_219 = 'b111101101;
    x_220 = 'b111100110;
    x_221 = 'b000000011;
    x_222 = 'b111110011;
    x_223 = 'b000000010;
    x_224 = 'b111111101;
    x_225 = 'b111110011;
    x_226 = 'b111101101;
    x_227 = 'b111100111;
    x_228 = 'b111100110;
    x_229 = 'b111001110;
    x_230 = 'b000001111;
    x_231 = 'b111100000;
    x_232 = 'b000001100;
    x_233 = 'b111110101;
    x_234 = 'b000010100;
    x_235 = 'b111000110;
    x_236 = 'b000001110;
    x_237 = 'b111110001;
    x_238 = 'b000101000;
    x_239 = 'b000101110;
    x_240 = 'b000101111;
    x_241 = 'b000111000;
    x_242 = 'b000101001;
    x_243 = 'b000011111;
    x_244 = 'b000011010;
    x_245 = 'b000001100;
    x_246 = 'b000001100;
    x_247 = 'b000110111;
    x_248 = 'b000111011;
    x_249 = 'b000111011;
    x_250 = 'b000100010;
    x_251 = 'b000011111;
    x_252 = 'b001001000;
    x_253 = 'b000111111;
    x_254 = 'b000101111;
    x_255 = 'b000111010;

    h_0 = 'b000001111;
    h_1 = 'b000010011;
    h_2 = 'b000000110;
    h_3 = 'b000000001;
    h_4 = 'b111111011;
    h_5 = 'b111110000;
    h_6 = 'b111110000;
    h_7 = 'b000101001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000000011;
    x_1 = 'b000001001;
    x_2 = 'b000000010;
    x_3 = 'b111111101;
    x_4 = 'b111111001;
    x_5 = 'b111101101;
    x_6 = 'b111101011;
    x_7 = 'b000011011;
    x_8 = 'b000011001;
    x_9 = 'b000010100;
    x_10 = 'b000010101;
    x_11 = 'b000001001;
    x_12 = 'b111111110;
    x_13 = 'b111100100;
    x_14 = 'b000100101;
    x_15 = 'b000100110;
    x_16 = 'b000100000;
    x_17 = 'b000010101;
    x_18 = 'b000010011;
    x_19 = 'b000001010;
    x_20 = 'b111111100;
    x_21 = 'b111111000;
    x_22 = 'b111101101;
    x_23 = 'b111101111;
    x_24 = 'b111111001;
    x_25 = 'b111111011;
    x_26 = 'b111101101;
    x_27 = 'b111110000;
    x_28 = 'b111101011;
    x_29 = 'b000000110;
    x_30 = 'b111110111;
    x_31 = 'b000000111;
    x_32 = 'b000000101;
    x_33 = 'b111111100;
    x_34 = 'b111110100;
    x_35 = 'b111110001;
    x_36 = 'b111101101;
    x_37 = 'b111011011;
    x_38 = 'b000010000;
    x_39 = 'b111100111;
    x_40 = 'b000010100;
    x_41 = 'b111101001;
    x_42 = 'b000011011;
    x_43 = 'b111101000;
    x_44 = 'b000001101;
    x_45 = 'b111101110;
    x_46 = 'b000100110;
    x_47 = 'b000101101;
    x_48 = 'b000101110;
    x_49 = 'b000110100;
    x_50 = 'b000101000;
    x_51 = 'b000011010;
    x_52 = 'b000010011;
    x_53 = 'b000000011;
    x_54 = 'b000000100;
    x_55 = 'b000111001;
    x_56 = 'b000111100;
    x_57 = 'b000111000;
    x_58 = 'b000011011;
    x_59 = 'b000011001;
    x_60 = 'b001000011;
    x_61 = 'b000111001;
    x_62 = 'b000101110;
    x_63 = 'b000110011;
    x_64 = 'b000000011;
    x_65 = 'b000001001;
    x_66 = 'b000000010;
    x_67 = 'b111111101;
    x_68 = 'b111111001;
    x_69 = 'b111101101;
    x_70 = 'b111101011;
    x_71 = 'b000011011;
    x_72 = 'b000011001;
    x_73 = 'b000010100;
    x_74 = 'b000010101;
    x_75 = 'b000001001;
    x_76 = 'b111111110;
    x_77 = 'b111100100;
    x_78 = 'b000100101;
    x_79 = 'b000100110;
    x_80 = 'b000100000;
    x_81 = 'b000010101;
    x_82 = 'b000010011;
    x_83 = 'b000001010;
    x_84 = 'b111111100;
    x_85 = 'b111111000;
    x_86 = 'b111101101;
    x_87 = 'b111101111;
    x_88 = 'b111111001;
    x_89 = 'b111111011;
    x_90 = 'b111101101;
    x_91 = 'b111110000;
    x_92 = 'b111101011;
    x_93 = 'b000000110;
    x_94 = 'b111110111;
    x_95 = 'b000000111;
    x_96 = 'b000000101;
    x_97 = 'b111111100;
    x_98 = 'b111110100;
    x_99 = 'b111110001;
    x_100 = 'b111101101;
    x_101 = 'b111011011;
    x_102 = 'b000010000;
    x_103 = 'b111100111;
    x_104 = 'b000010100;
    x_105 = 'b111101001;
    x_106 = 'b000011011;
    x_107 = 'b111101000;
    x_108 = 'b000001101;
    x_109 = 'b111101110;
    x_110 = 'b000100110;
    x_111 = 'b000101101;
    x_112 = 'b000101110;
    x_113 = 'b000110100;
    x_114 = 'b000101000;
    x_115 = 'b000011010;
    x_116 = 'b000010011;
    x_117 = 'b000000011;
    x_118 = 'b000000100;
    x_119 = 'b000111001;
    x_120 = 'b000111100;
    x_121 = 'b000111000;
    x_122 = 'b000011011;
    x_123 = 'b000011001;
    x_124 = 'b001000011;
    x_125 = 'b000111001;
    x_126 = 'b000101110;
    x_127 = 'b000110011;
    x_128 = 'b000000011;
    x_129 = 'b000001001;
    x_130 = 'b000000010;
    x_131 = 'b111111101;
    x_132 = 'b111111001;
    x_133 = 'b111101101;
    x_134 = 'b111101011;
    x_135 = 'b000011011;
    x_136 = 'b000011001;
    x_137 = 'b000010100;
    x_138 = 'b000010101;
    x_139 = 'b000001001;
    x_140 = 'b111111110;
    x_141 = 'b111100100;
    x_142 = 'b000100101;
    x_143 = 'b000100110;
    x_144 = 'b000100000;
    x_145 = 'b000010101;
    x_146 = 'b000010011;
    x_147 = 'b000001010;
    x_148 = 'b111111100;
    x_149 = 'b111111000;
    x_150 = 'b111101101;
    x_151 = 'b111101111;
    x_152 = 'b111111001;
    x_153 = 'b111111011;
    x_154 = 'b111101101;
    x_155 = 'b111110000;
    x_156 = 'b111101011;
    x_157 = 'b000000110;
    x_158 = 'b111110111;
    x_159 = 'b000000111;
    x_160 = 'b000000101;
    x_161 = 'b111111100;
    x_162 = 'b111110100;
    x_163 = 'b111110001;
    x_164 = 'b111101101;
    x_165 = 'b111011011;
    x_166 = 'b000010000;
    x_167 = 'b111100111;
    x_168 = 'b000010100;
    x_169 = 'b111101001;
    x_170 = 'b000011011;
    x_171 = 'b111101000;
    x_172 = 'b000001101;
    x_173 = 'b111101110;
    x_174 = 'b000100110;
    x_175 = 'b000101101;
    x_176 = 'b000101110;
    x_177 = 'b000110100;
    x_178 = 'b000101000;
    x_179 = 'b000011010;
    x_180 = 'b000010011;
    x_181 = 'b000000011;
    x_182 = 'b000000100;
    x_183 = 'b000111001;
    x_184 = 'b000111100;
    x_185 = 'b000111000;
    x_186 = 'b000011011;
    x_187 = 'b000011001;
    x_188 = 'b001000011;
    x_189 = 'b000111001;
    x_190 = 'b000101110;
    x_191 = 'b000110011;
    x_192 = 'b000000011;
    x_193 = 'b000001001;
    x_194 = 'b000000010;
    x_195 = 'b111111101;
    x_196 = 'b111111001;
    x_197 = 'b111101101;
    x_198 = 'b111101011;
    x_199 = 'b000011011;
    x_200 = 'b000011001;
    x_201 = 'b000010100;
    x_202 = 'b000010101;
    x_203 = 'b000001001;
    x_204 = 'b111111110;
    x_205 = 'b111100100;
    x_206 = 'b000100101;
    x_207 = 'b000100110;
    x_208 = 'b000100000;
    x_209 = 'b000010101;
    x_210 = 'b000010011;
    x_211 = 'b000001010;
    x_212 = 'b111111100;
    x_213 = 'b111111000;
    x_214 = 'b111101101;
    x_215 = 'b111101111;
    x_216 = 'b111111001;
    x_217 = 'b111111011;
    x_218 = 'b111101101;
    x_219 = 'b111110000;
    x_220 = 'b111101011;
    x_221 = 'b000000110;
    x_222 = 'b111110111;
    x_223 = 'b000000111;
    x_224 = 'b000000101;
    x_225 = 'b111111100;
    x_226 = 'b111110100;
    x_227 = 'b111110001;
    x_228 = 'b111101101;
    x_229 = 'b111011011;
    x_230 = 'b000010000;
    x_231 = 'b111100111;
    x_232 = 'b000010100;
    x_233 = 'b111101001;
    x_234 = 'b000011011;
    x_235 = 'b111101000;
    x_236 = 'b000001101;
    x_237 = 'b111101110;
    x_238 = 'b000100110;
    x_239 = 'b000101101;
    x_240 = 'b000101110;
    x_241 = 'b000110100;
    x_242 = 'b000101000;
    x_243 = 'b000011010;
    x_244 = 'b000010011;
    x_245 = 'b000000011;
    x_246 = 'b000000100;
    x_247 = 'b000111001;
    x_248 = 'b000111100;
    x_249 = 'b000111000;
    x_250 = 'b000011011;
    x_251 = 'b000011001;
    x_252 = 'b001000011;
    x_253 = 'b000111001;
    x_254 = 'b000101110;
    x_255 = 'b000110011;

    h_0 = 'b000000011;
    h_1 = 'b000001001;
    h_2 = 'b000000010;
    h_3 = 'b111111101;
    h_4 = 'b111111001;
    h_5 = 'b111101101;
    h_6 = 'b111101011;
    h_7 = 'b000011011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000010001;
    x_1 = 'b000011101;
    x_2 = 'b000010111;
    x_3 = 'b000010011;
    x_4 = 'b000001011;
    x_5 = 'b111111011;
    x_6 = 'b111101111;
    x_7 = 'b000110010;
    x_8 = 'b000101100;
    x_9 = 'b000100111;
    x_10 = 'b000100010;
    x_11 = 'b000010111;
    x_12 = 'b000000110;
    x_13 = 'b111100011;
    x_14 = 'b000111100;
    x_15 = 'b000110100;
    x_16 = 'b000101101;
    x_17 = 'b000100001;
    x_18 = 'b000011101;
    x_19 = 'b000010010;
    x_20 = 'b000000001;
    x_21 = 'b111111001;
    x_22 = 'b111110000;
    x_23 = 'b111110100;
    x_24 = 'b111111110;
    x_25 = 'b000000000;
    x_26 = 'b111111010;
    x_27 = 'b111111010;
    x_28 = 'b111110010;
    x_29 = 'b000001110;
    x_30 = 'b000000000;
    x_31 = 'b000010110;
    x_32 = 'b000010011;
    x_33 = 'b000001011;
    x_34 = 'b000000011;
    x_35 = 'b111111101;
    x_36 = 'b111110110;
    x_37 = 'b111100000;
    x_38 = 'b000010101;
    x_39 = 'b111101011;
    x_40 = 'b000010011;
    x_41 = 'b111100111;
    x_42 = 'b000011111;
    x_43 = 'b111110010;
    x_44 = 'b000011100;
    x_45 = 'b000000001;
    x_46 = 'b000110111;
    x_47 = 'b000111100;
    x_48 = 'b000110111;
    x_49 = 'b001000000;
    x_50 = 'b000110011;
    x_51 = 'b000100111;
    x_52 = 'b000100010;
    x_53 = 'b000010001;
    x_54 = 'b000010001;
    x_55 = 'b001000011;
    x_56 = 'b001000110;
    x_57 = 'b001000001;
    x_58 = 'b000100011;
    x_59 = 'b000100000;
    x_60 = 'b001000011;
    x_61 = 'b000111000;
    x_62 = 'b000110000;
    x_63 = 'b000110100;
    x_64 = 'b000010001;
    x_65 = 'b000011101;
    x_66 = 'b000010111;
    x_67 = 'b000010011;
    x_68 = 'b000001011;
    x_69 = 'b111111011;
    x_70 = 'b111101111;
    x_71 = 'b000110010;
    x_72 = 'b000101100;
    x_73 = 'b000100111;
    x_74 = 'b000100010;
    x_75 = 'b000010111;
    x_76 = 'b000000110;
    x_77 = 'b111100011;
    x_78 = 'b000111100;
    x_79 = 'b000110100;
    x_80 = 'b000101101;
    x_81 = 'b000100001;
    x_82 = 'b000011101;
    x_83 = 'b000010010;
    x_84 = 'b000000001;
    x_85 = 'b111111001;
    x_86 = 'b111110000;
    x_87 = 'b111110100;
    x_88 = 'b111111110;
    x_89 = 'b000000000;
    x_90 = 'b111111010;
    x_91 = 'b111111010;
    x_92 = 'b111110010;
    x_93 = 'b000001110;
    x_94 = 'b000000000;
    x_95 = 'b000010110;
    x_96 = 'b000010011;
    x_97 = 'b000001011;
    x_98 = 'b000000011;
    x_99 = 'b111111101;
    x_100 = 'b111110110;
    x_101 = 'b111100000;
    x_102 = 'b000010101;
    x_103 = 'b111101011;
    x_104 = 'b000010011;
    x_105 = 'b111100111;
    x_106 = 'b000011111;
    x_107 = 'b111110010;
    x_108 = 'b000011100;
    x_109 = 'b000000001;
    x_110 = 'b000110111;
    x_111 = 'b000111100;
    x_112 = 'b000110111;
    x_113 = 'b001000000;
    x_114 = 'b000110011;
    x_115 = 'b000100111;
    x_116 = 'b000100010;
    x_117 = 'b000010001;
    x_118 = 'b000010001;
    x_119 = 'b001000011;
    x_120 = 'b001000110;
    x_121 = 'b001000001;
    x_122 = 'b000100011;
    x_123 = 'b000100000;
    x_124 = 'b001000011;
    x_125 = 'b000111000;
    x_126 = 'b000110000;
    x_127 = 'b000110100;
    x_128 = 'b000010001;
    x_129 = 'b000011101;
    x_130 = 'b000010111;
    x_131 = 'b000010011;
    x_132 = 'b000001011;
    x_133 = 'b111111011;
    x_134 = 'b111101111;
    x_135 = 'b000110010;
    x_136 = 'b000101100;
    x_137 = 'b000100111;
    x_138 = 'b000100010;
    x_139 = 'b000010111;
    x_140 = 'b000000110;
    x_141 = 'b111100011;
    x_142 = 'b000111100;
    x_143 = 'b000110100;
    x_144 = 'b000101101;
    x_145 = 'b000100001;
    x_146 = 'b000011101;
    x_147 = 'b000010010;
    x_148 = 'b000000001;
    x_149 = 'b111111001;
    x_150 = 'b111110000;
    x_151 = 'b111110100;
    x_152 = 'b111111110;
    x_153 = 'b000000000;
    x_154 = 'b111111010;
    x_155 = 'b111111010;
    x_156 = 'b111110010;
    x_157 = 'b000001110;
    x_158 = 'b000000000;
    x_159 = 'b000010110;
    x_160 = 'b000010011;
    x_161 = 'b000001011;
    x_162 = 'b000000011;
    x_163 = 'b111111101;
    x_164 = 'b111110110;
    x_165 = 'b111100000;
    x_166 = 'b000010101;
    x_167 = 'b111101011;
    x_168 = 'b000010011;
    x_169 = 'b111100111;
    x_170 = 'b000011111;
    x_171 = 'b111110010;
    x_172 = 'b000011100;
    x_173 = 'b000000001;
    x_174 = 'b000110111;
    x_175 = 'b000111100;
    x_176 = 'b000110111;
    x_177 = 'b001000000;
    x_178 = 'b000110011;
    x_179 = 'b000100111;
    x_180 = 'b000100010;
    x_181 = 'b000010001;
    x_182 = 'b000010001;
    x_183 = 'b001000011;
    x_184 = 'b001000110;
    x_185 = 'b001000001;
    x_186 = 'b000100011;
    x_187 = 'b000100000;
    x_188 = 'b001000011;
    x_189 = 'b000111000;
    x_190 = 'b000110000;
    x_191 = 'b000110100;
    x_192 = 'b000010001;
    x_193 = 'b000011101;
    x_194 = 'b000010111;
    x_195 = 'b000010011;
    x_196 = 'b000001011;
    x_197 = 'b111111011;
    x_198 = 'b111101111;
    x_199 = 'b000110010;
    x_200 = 'b000101100;
    x_201 = 'b000100111;
    x_202 = 'b000100010;
    x_203 = 'b000010111;
    x_204 = 'b000000110;
    x_205 = 'b111100011;
    x_206 = 'b000111100;
    x_207 = 'b000110100;
    x_208 = 'b000101101;
    x_209 = 'b000100001;
    x_210 = 'b000011101;
    x_211 = 'b000010010;
    x_212 = 'b000000001;
    x_213 = 'b111111001;
    x_214 = 'b111110000;
    x_215 = 'b111110100;
    x_216 = 'b111111110;
    x_217 = 'b000000000;
    x_218 = 'b111111010;
    x_219 = 'b111111010;
    x_220 = 'b111110010;
    x_221 = 'b000001110;
    x_222 = 'b000000000;
    x_223 = 'b000010110;
    x_224 = 'b000010011;
    x_225 = 'b000001011;
    x_226 = 'b000000011;
    x_227 = 'b111111101;
    x_228 = 'b111110110;
    x_229 = 'b111100000;
    x_230 = 'b000010101;
    x_231 = 'b111101011;
    x_232 = 'b000010011;
    x_233 = 'b111100111;
    x_234 = 'b000011111;
    x_235 = 'b111110010;
    x_236 = 'b000011100;
    x_237 = 'b000000001;
    x_238 = 'b000110111;
    x_239 = 'b000111100;
    x_240 = 'b000110111;
    x_241 = 'b001000000;
    x_242 = 'b000110011;
    x_243 = 'b000100111;
    x_244 = 'b000100010;
    x_245 = 'b000010001;
    x_246 = 'b000010001;
    x_247 = 'b001000011;
    x_248 = 'b001000110;
    x_249 = 'b001000001;
    x_250 = 'b000100011;
    x_251 = 'b000100000;
    x_252 = 'b001000011;
    x_253 = 'b000111000;
    x_254 = 'b000110000;
    x_255 = 'b000110100;

    h_0 = 'b000010001;
    h_1 = 'b000011101;
    h_2 = 'b000010111;
    h_3 = 'b000010011;
    h_4 = 'b000001011;
    h_5 = 'b111111011;
    h_6 = 'b111101111;
    h_7 = 'b000110010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000010110;
    x_1 = 'b000011011;
    x_2 = 'b000010101;
    x_3 = 'b000010101;
    x_4 = 'b000001110;
    x_5 = 'b000000001;
    x_6 = 'b111111100;
    x_7 = 'b000100111;
    x_8 = 'b000100011;
    x_9 = 'b000100000;
    x_10 = 'b000011111;
    x_11 = 'b000011001;
    x_12 = 'b000001101;
    x_13 = 'b111111000;
    x_14 = 'b000101100;
    x_15 = 'b000101001;
    x_16 = 'b000100111;
    x_17 = 'b000011101;
    x_18 = 'b000100001;
    x_19 = 'b000011100;
    x_20 = 'b000010010;
    x_21 = 'b111110110;
    x_22 = 'b111101100;
    x_23 = 'b111110010;
    x_24 = 'b111111001;
    x_25 = 'b111111011;
    x_26 = 'b111110011;
    x_27 = 'b111110111;
    x_28 = 'b111110001;
    x_29 = 'b000001110;
    x_30 = 'b111111101;
    x_31 = 'b000001111;
    x_32 = 'b000000111;
    x_33 = 'b000000010;
    x_34 = 'b111111100;
    x_35 = 'b111110110;
    x_36 = 'b111110011;
    x_37 = 'b111100001;
    x_38 = 'b000011100;
    x_39 = 'b111111000;
    x_40 = 'b000101001;
    x_41 = 'b000011011;
    x_42 = 'b000101101;
    x_43 = 'b111110101;
    x_44 = 'b000011110;
    x_45 = 'b000001101;
    x_46 = 'b000101100;
    x_47 = 'b000101101;
    x_48 = 'b000100110;
    x_49 = 'b000110101;
    x_50 = 'b000101000;
    x_51 = 'b000100010;
    x_52 = 'b000100001;
    x_53 = 'b000010101;
    x_54 = 'b000010110;
    x_55 = 'b000110100;
    x_56 = 'b000111001;
    x_57 = 'b000110111;
    x_58 = 'b000100001;
    x_59 = 'b000100000;
    x_60 = 'b001000010;
    x_61 = 'b000111001;
    x_62 = 'b000110001;
    x_63 = 'b000110101;
    x_64 = 'b000010110;
    x_65 = 'b000011011;
    x_66 = 'b000010101;
    x_67 = 'b000010101;
    x_68 = 'b000001110;
    x_69 = 'b000000001;
    x_70 = 'b111111100;
    x_71 = 'b000100111;
    x_72 = 'b000100011;
    x_73 = 'b000100000;
    x_74 = 'b000011111;
    x_75 = 'b000011001;
    x_76 = 'b000001101;
    x_77 = 'b111111000;
    x_78 = 'b000101100;
    x_79 = 'b000101001;
    x_80 = 'b000100111;
    x_81 = 'b000011101;
    x_82 = 'b000100001;
    x_83 = 'b000011100;
    x_84 = 'b000010010;
    x_85 = 'b111110110;
    x_86 = 'b111101100;
    x_87 = 'b111110010;
    x_88 = 'b111111001;
    x_89 = 'b111111011;
    x_90 = 'b111110011;
    x_91 = 'b111110111;
    x_92 = 'b111110001;
    x_93 = 'b000001110;
    x_94 = 'b111111101;
    x_95 = 'b000001111;
    x_96 = 'b000000111;
    x_97 = 'b000000010;
    x_98 = 'b111111100;
    x_99 = 'b111110110;
    x_100 = 'b111110011;
    x_101 = 'b111100001;
    x_102 = 'b000011100;
    x_103 = 'b111111000;
    x_104 = 'b000101001;
    x_105 = 'b000011011;
    x_106 = 'b000101101;
    x_107 = 'b111110101;
    x_108 = 'b000011110;
    x_109 = 'b000001101;
    x_110 = 'b000101100;
    x_111 = 'b000101101;
    x_112 = 'b000100110;
    x_113 = 'b000110101;
    x_114 = 'b000101000;
    x_115 = 'b000100010;
    x_116 = 'b000100001;
    x_117 = 'b000010101;
    x_118 = 'b000010110;
    x_119 = 'b000110100;
    x_120 = 'b000111001;
    x_121 = 'b000110111;
    x_122 = 'b000100001;
    x_123 = 'b000100000;
    x_124 = 'b001000010;
    x_125 = 'b000111001;
    x_126 = 'b000110001;
    x_127 = 'b000110101;
    x_128 = 'b000010110;
    x_129 = 'b000011011;
    x_130 = 'b000010101;
    x_131 = 'b000010101;
    x_132 = 'b000001110;
    x_133 = 'b000000001;
    x_134 = 'b111111100;
    x_135 = 'b000100111;
    x_136 = 'b000100011;
    x_137 = 'b000100000;
    x_138 = 'b000011111;
    x_139 = 'b000011001;
    x_140 = 'b000001101;
    x_141 = 'b111111000;
    x_142 = 'b000101100;
    x_143 = 'b000101001;
    x_144 = 'b000100111;
    x_145 = 'b000011101;
    x_146 = 'b000100001;
    x_147 = 'b000011100;
    x_148 = 'b000010010;
    x_149 = 'b111110110;
    x_150 = 'b111101100;
    x_151 = 'b111110010;
    x_152 = 'b111111001;
    x_153 = 'b111111011;
    x_154 = 'b111110011;
    x_155 = 'b111110111;
    x_156 = 'b111110001;
    x_157 = 'b000001110;
    x_158 = 'b111111101;
    x_159 = 'b000001111;
    x_160 = 'b000000111;
    x_161 = 'b000000010;
    x_162 = 'b111111100;
    x_163 = 'b111110110;
    x_164 = 'b111110011;
    x_165 = 'b111100001;
    x_166 = 'b000011100;
    x_167 = 'b111111000;
    x_168 = 'b000101001;
    x_169 = 'b000011011;
    x_170 = 'b000101101;
    x_171 = 'b111110101;
    x_172 = 'b000011110;
    x_173 = 'b000001101;
    x_174 = 'b000101100;
    x_175 = 'b000101101;
    x_176 = 'b000100110;
    x_177 = 'b000110101;
    x_178 = 'b000101000;
    x_179 = 'b000100010;
    x_180 = 'b000100001;
    x_181 = 'b000010101;
    x_182 = 'b000010110;
    x_183 = 'b000110100;
    x_184 = 'b000111001;
    x_185 = 'b000110111;
    x_186 = 'b000100001;
    x_187 = 'b000100000;
    x_188 = 'b001000010;
    x_189 = 'b000111001;
    x_190 = 'b000110001;
    x_191 = 'b000110101;
    x_192 = 'b000010110;
    x_193 = 'b000011011;
    x_194 = 'b000010101;
    x_195 = 'b000010101;
    x_196 = 'b000001110;
    x_197 = 'b000000001;
    x_198 = 'b111111100;
    x_199 = 'b000100111;
    x_200 = 'b000100011;
    x_201 = 'b000100000;
    x_202 = 'b000011111;
    x_203 = 'b000011001;
    x_204 = 'b000001101;
    x_205 = 'b111111000;
    x_206 = 'b000101100;
    x_207 = 'b000101001;
    x_208 = 'b000100111;
    x_209 = 'b000011101;
    x_210 = 'b000100001;
    x_211 = 'b000011100;
    x_212 = 'b000010010;
    x_213 = 'b111110110;
    x_214 = 'b111101100;
    x_215 = 'b111110010;
    x_216 = 'b111111001;
    x_217 = 'b111111011;
    x_218 = 'b111110011;
    x_219 = 'b111110111;
    x_220 = 'b111110001;
    x_221 = 'b000001110;
    x_222 = 'b111111101;
    x_223 = 'b000001111;
    x_224 = 'b000000111;
    x_225 = 'b000000010;
    x_226 = 'b111111100;
    x_227 = 'b111110110;
    x_228 = 'b111110011;
    x_229 = 'b111100001;
    x_230 = 'b000011100;
    x_231 = 'b111111000;
    x_232 = 'b000101001;
    x_233 = 'b000011011;
    x_234 = 'b000101101;
    x_235 = 'b111110101;
    x_236 = 'b000011110;
    x_237 = 'b000001101;
    x_238 = 'b000101100;
    x_239 = 'b000101101;
    x_240 = 'b000100110;
    x_241 = 'b000110101;
    x_242 = 'b000101000;
    x_243 = 'b000100010;
    x_244 = 'b000100001;
    x_245 = 'b000010101;
    x_246 = 'b000010110;
    x_247 = 'b000110100;
    x_248 = 'b000111001;
    x_249 = 'b000110111;
    x_250 = 'b000100001;
    x_251 = 'b000100000;
    x_252 = 'b001000010;
    x_253 = 'b000111001;
    x_254 = 'b000110001;
    x_255 = 'b000110101;

    h_0 = 'b000010110;
    h_1 = 'b000011011;
    h_2 = 'b000010101;
    h_3 = 'b000010101;
    h_4 = 'b000001110;
    h_5 = 'b000000001;
    h_6 = 'b111111100;
    h_7 = 'b000100111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000010100;
    x_1 = 'b000010101;
    x_2 = 'b000001110;
    x_3 = 'b000001111;
    x_4 = 'b000001001;
    x_5 = 'b000000000;
    x_6 = 'b000001000;
    x_7 = 'b000011110;
    x_8 = 'b000011010;
    x_9 = 'b000010111;
    x_10 = 'b000011001;
    x_11 = 'b000011010;
    x_12 = 'b000010010;
    x_13 = 'b000001101;
    x_14 = 'b000011111;
    x_15 = 'b000011111;
    x_16 = 'b000011110;
    x_17 = 'b000011001;
    x_18 = 'b000100001;
    x_19 = 'b000100000;
    x_20 = 'b000100010;
    x_21 = 'b111111010;
    x_22 = 'b111110000;
    x_23 = 'b111110100;
    x_24 = 'b111111111;
    x_25 = 'b000000000;
    x_26 = 'b111111001;
    x_27 = 'b111111010;
    x_28 = 'b111110010;
    x_29 = 'b000010100;
    x_30 = 'b000000011;
    x_31 = 'b000010100;
    x_32 = 'b000001111;
    x_33 = 'b000001001;
    x_34 = 'b000000011;
    x_35 = 'b111111111;
    x_36 = 'b111111100;
    x_37 = 'b111101001;
    x_38 = 'b000011110;
    x_39 = 'b000001010;
    x_40 = 'b000100100;
    x_41 = 'b000101011;
    x_42 = 'b000101101;
    x_43 = 'b000000110;
    x_44 = 'b000010010;
    x_45 = 'b000011011;
    x_46 = 'b000100111;
    x_47 = 'b000101010;
    x_48 = 'b000100101;
    x_49 = 'b000110011;
    x_50 = 'b000101001;
    x_51 = 'b000100110;
    x_52 = 'b000101001;
    x_53 = 'b000100001;
    x_54 = 'b000100011;
    x_55 = 'b000101111;
    x_56 = 'b000110011;
    x_57 = 'b000110100;
    x_58 = 'b000100101;
    x_59 = 'b000100110;
    x_60 = 'b000111011;
    x_61 = 'b000110101;
    x_62 = 'b000110011;
    x_63 = 'b000110000;
    x_64 = 'b000010100;
    x_65 = 'b000010101;
    x_66 = 'b000001110;
    x_67 = 'b000001111;
    x_68 = 'b000001001;
    x_69 = 'b000000000;
    x_70 = 'b000001000;
    x_71 = 'b000011110;
    x_72 = 'b000011010;
    x_73 = 'b000010111;
    x_74 = 'b000011001;
    x_75 = 'b000011010;
    x_76 = 'b000010010;
    x_77 = 'b000001101;
    x_78 = 'b000011111;
    x_79 = 'b000011111;
    x_80 = 'b000011110;
    x_81 = 'b000011001;
    x_82 = 'b000100001;
    x_83 = 'b000100000;
    x_84 = 'b000100010;
    x_85 = 'b111111010;
    x_86 = 'b111110000;
    x_87 = 'b111110100;
    x_88 = 'b111111111;
    x_89 = 'b000000000;
    x_90 = 'b111111001;
    x_91 = 'b111111010;
    x_92 = 'b111110010;
    x_93 = 'b000010100;
    x_94 = 'b000000011;
    x_95 = 'b000010100;
    x_96 = 'b000001111;
    x_97 = 'b000001001;
    x_98 = 'b000000011;
    x_99 = 'b111111111;
    x_100 = 'b111111100;
    x_101 = 'b111101001;
    x_102 = 'b000011110;
    x_103 = 'b000001010;
    x_104 = 'b000100100;
    x_105 = 'b000101011;
    x_106 = 'b000101101;
    x_107 = 'b000000110;
    x_108 = 'b000010010;
    x_109 = 'b000011011;
    x_110 = 'b000100111;
    x_111 = 'b000101010;
    x_112 = 'b000100101;
    x_113 = 'b000110011;
    x_114 = 'b000101001;
    x_115 = 'b000100110;
    x_116 = 'b000101001;
    x_117 = 'b000100001;
    x_118 = 'b000100011;
    x_119 = 'b000101111;
    x_120 = 'b000110011;
    x_121 = 'b000110100;
    x_122 = 'b000100101;
    x_123 = 'b000100110;
    x_124 = 'b000111011;
    x_125 = 'b000110101;
    x_126 = 'b000110011;
    x_127 = 'b000110000;
    x_128 = 'b000010100;
    x_129 = 'b000010101;
    x_130 = 'b000001110;
    x_131 = 'b000001111;
    x_132 = 'b000001001;
    x_133 = 'b000000000;
    x_134 = 'b000001000;
    x_135 = 'b000011110;
    x_136 = 'b000011010;
    x_137 = 'b000010111;
    x_138 = 'b000011001;
    x_139 = 'b000011010;
    x_140 = 'b000010010;
    x_141 = 'b000001101;
    x_142 = 'b000011111;
    x_143 = 'b000011111;
    x_144 = 'b000011110;
    x_145 = 'b000011001;
    x_146 = 'b000100001;
    x_147 = 'b000100000;
    x_148 = 'b000100010;
    x_149 = 'b111111010;
    x_150 = 'b111110000;
    x_151 = 'b111110100;
    x_152 = 'b111111111;
    x_153 = 'b000000000;
    x_154 = 'b111111001;
    x_155 = 'b111111010;
    x_156 = 'b111110010;
    x_157 = 'b000010100;
    x_158 = 'b000000011;
    x_159 = 'b000010100;
    x_160 = 'b000001111;
    x_161 = 'b000001001;
    x_162 = 'b000000011;
    x_163 = 'b111111111;
    x_164 = 'b111111100;
    x_165 = 'b111101001;
    x_166 = 'b000011110;
    x_167 = 'b000001010;
    x_168 = 'b000100100;
    x_169 = 'b000101011;
    x_170 = 'b000101101;
    x_171 = 'b000000110;
    x_172 = 'b000010010;
    x_173 = 'b000011011;
    x_174 = 'b000100111;
    x_175 = 'b000101010;
    x_176 = 'b000100101;
    x_177 = 'b000110011;
    x_178 = 'b000101001;
    x_179 = 'b000100110;
    x_180 = 'b000101001;
    x_181 = 'b000100001;
    x_182 = 'b000100011;
    x_183 = 'b000101111;
    x_184 = 'b000110011;
    x_185 = 'b000110100;
    x_186 = 'b000100101;
    x_187 = 'b000100110;
    x_188 = 'b000111011;
    x_189 = 'b000110101;
    x_190 = 'b000110011;
    x_191 = 'b000110000;
    x_192 = 'b000010100;
    x_193 = 'b000010101;
    x_194 = 'b000001110;
    x_195 = 'b000001111;
    x_196 = 'b000001001;
    x_197 = 'b000000000;
    x_198 = 'b000001000;
    x_199 = 'b000011110;
    x_200 = 'b000011010;
    x_201 = 'b000010111;
    x_202 = 'b000011001;
    x_203 = 'b000011010;
    x_204 = 'b000010010;
    x_205 = 'b000001101;
    x_206 = 'b000011111;
    x_207 = 'b000011111;
    x_208 = 'b000011110;
    x_209 = 'b000011001;
    x_210 = 'b000100001;
    x_211 = 'b000100000;
    x_212 = 'b000100010;
    x_213 = 'b111111010;
    x_214 = 'b111110000;
    x_215 = 'b111110100;
    x_216 = 'b111111111;
    x_217 = 'b000000000;
    x_218 = 'b111111001;
    x_219 = 'b111111010;
    x_220 = 'b111110010;
    x_221 = 'b000010100;
    x_222 = 'b000000011;
    x_223 = 'b000010100;
    x_224 = 'b000001111;
    x_225 = 'b000001001;
    x_226 = 'b000000011;
    x_227 = 'b111111111;
    x_228 = 'b111111100;
    x_229 = 'b111101001;
    x_230 = 'b000011110;
    x_231 = 'b000001010;
    x_232 = 'b000100100;
    x_233 = 'b000101011;
    x_234 = 'b000101101;
    x_235 = 'b000000110;
    x_236 = 'b000010010;
    x_237 = 'b000011011;
    x_238 = 'b000100111;
    x_239 = 'b000101010;
    x_240 = 'b000100101;
    x_241 = 'b000110011;
    x_242 = 'b000101001;
    x_243 = 'b000100110;
    x_244 = 'b000101001;
    x_245 = 'b000100001;
    x_246 = 'b000100011;
    x_247 = 'b000101111;
    x_248 = 'b000110011;
    x_249 = 'b000110100;
    x_250 = 'b000100101;
    x_251 = 'b000100110;
    x_252 = 'b000111011;
    x_253 = 'b000110101;
    x_254 = 'b000110011;
    x_255 = 'b000110000;

    h_0 = 'b000010100;
    h_1 = 'b000010101;
    h_2 = 'b000001110;
    h_3 = 'b000001111;
    h_4 = 'b000001001;
    h_5 = 'b000000000;
    h_6 = 'b000001000;
    h_7 = 'b000011110;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000011100;
    x_1 = 'b000100000;
    x_2 = 'b000011100;
    x_3 = 'b000011010;
    x_4 = 'b000010011;
    x_5 = 'b000001100;
    x_6 = 'b000010010;
    x_7 = 'b000101001;
    x_8 = 'b000100110;
    x_9 = 'b000100001;
    x_10 = 'b000100001;
    x_11 = 'b000011111;
    x_12 = 'b000011100;
    x_13 = 'b000010000;
    x_14 = 'b000101000;
    x_15 = 'b000100100;
    x_16 = 'b000100001;
    x_17 = 'b000011101;
    x_18 = 'b000100010;
    x_19 = 'b000100010;
    x_20 = 'b000100100;
    x_21 = 'b111111011;
    x_22 = 'b111101111;
    x_23 = 'b111110001;
    x_24 = 'b111111110;
    x_25 = 'b000000001;
    x_26 = 'b111111100;
    x_27 = 'b111111101;
    x_28 = 'b111110001;
    x_29 = 'b000001111;
    x_30 = 'b000000110;
    x_31 = 'b000011011;
    x_32 = 'b000010010;
    x_33 = 'b000001011;
    x_34 = 'b000000110;
    x_35 = 'b000000010;
    x_36 = 'b000000010;
    x_37 = 'b111110011;
    x_38 = 'b000100010;
    x_39 = 'b000000111;
    x_40 = 'b000101010;
    x_41 = 'b000010101;
    x_42 = 'b000011100;
    x_43 = 'b000010110;
    x_44 = 'b000010001;
    x_45 = 'b000011100;
    x_46 = 'b000100011;
    x_47 = 'b000100011;
    x_48 = 'b000011110;
    x_49 = 'b000101001;
    x_50 = 'b000100000;
    x_51 = 'b000011100;
    x_52 = 'b000011110;
    x_53 = 'b000010111;
    x_54 = 'b000011001;
    x_55 = 'b000100001;
    x_56 = 'b000100101;
    x_57 = 'b000100011;
    x_58 = 'b000011000;
    x_59 = 'b000010101;
    x_60 = 'b000101010;
    x_61 = 'b000011111;
    x_62 = 'b000100100;
    x_63 = 'b000010111;
    x_64 = 'b000011100;
    x_65 = 'b000100000;
    x_66 = 'b000011100;
    x_67 = 'b000011010;
    x_68 = 'b000010011;
    x_69 = 'b000001100;
    x_70 = 'b000010010;
    x_71 = 'b000101001;
    x_72 = 'b000100110;
    x_73 = 'b000100001;
    x_74 = 'b000100001;
    x_75 = 'b000011111;
    x_76 = 'b000011100;
    x_77 = 'b000010000;
    x_78 = 'b000101000;
    x_79 = 'b000100100;
    x_80 = 'b000100001;
    x_81 = 'b000011101;
    x_82 = 'b000100010;
    x_83 = 'b000100010;
    x_84 = 'b000100100;
    x_85 = 'b111111011;
    x_86 = 'b111101111;
    x_87 = 'b111110001;
    x_88 = 'b111111110;
    x_89 = 'b000000001;
    x_90 = 'b111111100;
    x_91 = 'b111111101;
    x_92 = 'b111110001;
    x_93 = 'b000001111;
    x_94 = 'b000000110;
    x_95 = 'b000011011;
    x_96 = 'b000010010;
    x_97 = 'b000001011;
    x_98 = 'b000000110;
    x_99 = 'b000000010;
    x_100 = 'b000000010;
    x_101 = 'b111110011;
    x_102 = 'b000100010;
    x_103 = 'b000000111;
    x_104 = 'b000101010;
    x_105 = 'b000010101;
    x_106 = 'b000011100;
    x_107 = 'b000010110;
    x_108 = 'b000010001;
    x_109 = 'b000011100;
    x_110 = 'b000100011;
    x_111 = 'b000100011;
    x_112 = 'b000011110;
    x_113 = 'b000101001;
    x_114 = 'b000100000;
    x_115 = 'b000011100;
    x_116 = 'b000011110;
    x_117 = 'b000010111;
    x_118 = 'b000011001;
    x_119 = 'b000100001;
    x_120 = 'b000100101;
    x_121 = 'b000100011;
    x_122 = 'b000011000;
    x_123 = 'b000010101;
    x_124 = 'b000101010;
    x_125 = 'b000011111;
    x_126 = 'b000100100;
    x_127 = 'b000010111;
    x_128 = 'b000011100;
    x_129 = 'b000100000;
    x_130 = 'b000011100;
    x_131 = 'b000011010;
    x_132 = 'b000010011;
    x_133 = 'b000001100;
    x_134 = 'b000010010;
    x_135 = 'b000101001;
    x_136 = 'b000100110;
    x_137 = 'b000100001;
    x_138 = 'b000100001;
    x_139 = 'b000011111;
    x_140 = 'b000011100;
    x_141 = 'b000010000;
    x_142 = 'b000101000;
    x_143 = 'b000100100;
    x_144 = 'b000100001;
    x_145 = 'b000011101;
    x_146 = 'b000100010;
    x_147 = 'b000100010;
    x_148 = 'b000100100;
    x_149 = 'b111111011;
    x_150 = 'b111101111;
    x_151 = 'b111110001;
    x_152 = 'b111111110;
    x_153 = 'b000000001;
    x_154 = 'b111111100;
    x_155 = 'b111111101;
    x_156 = 'b111110001;
    x_157 = 'b000001111;
    x_158 = 'b000000110;
    x_159 = 'b000011011;
    x_160 = 'b000010010;
    x_161 = 'b000001011;
    x_162 = 'b000000110;
    x_163 = 'b000000010;
    x_164 = 'b000000010;
    x_165 = 'b111110011;
    x_166 = 'b000100010;
    x_167 = 'b000000111;
    x_168 = 'b000101010;
    x_169 = 'b000010101;
    x_170 = 'b000011100;
    x_171 = 'b000010110;
    x_172 = 'b000010001;
    x_173 = 'b000011100;
    x_174 = 'b000100011;
    x_175 = 'b000100011;
    x_176 = 'b000011110;
    x_177 = 'b000101001;
    x_178 = 'b000100000;
    x_179 = 'b000011100;
    x_180 = 'b000011110;
    x_181 = 'b000010111;
    x_182 = 'b000011001;
    x_183 = 'b000100001;
    x_184 = 'b000100101;
    x_185 = 'b000100011;
    x_186 = 'b000011000;
    x_187 = 'b000010101;
    x_188 = 'b000101010;
    x_189 = 'b000011111;
    x_190 = 'b000100100;
    x_191 = 'b000010111;
    x_192 = 'b000011100;
    x_193 = 'b000100000;
    x_194 = 'b000011100;
    x_195 = 'b000011010;
    x_196 = 'b000010011;
    x_197 = 'b000001100;
    x_198 = 'b000010010;
    x_199 = 'b000101001;
    x_200 = 'b000100110;
    x_201 = 'b000100001;
    x_202 = 'b000100001;
    x_203 = 'b000011111;
    x_204 = 'b000011100;
    x_205 = 'b000010000;
    x_206 = 'b000101000;
    x_207 = 'b000100100;
    x_208 = 'b000100001;
    x_209 = 'b000011101;
    x_210 = 'b000100010;
    x_211 = 'b000100010;
    x_212 = 'b000100100;
    x_213 = 'b111111011;
    x_214 = 'b111101111;
    x_215 = 'b111110001;
    x_216 = 'b111111110;
    x_217 = 'b000000001;
    x_218 = 'b111111100;
    x_219 = 'b111111101;
    x_220 = 'b111110001;
    x_221 = 'b000001111;
    x_222 = 'b000000110;
    x_223 = 'b000011011;
    x_224 = 'b000010010;
    x_225 = 'b000001011;
    x_226 = 'b000000110;
    x_227 = 'b000000010;
    x_228 = 'b000000010;
    x_229 = 'b111110011;
    x_230 = 'b000100010;
    x_231 = 'b000000111;
    x_232 = 'b000101010;
    x_233 = 'b000010101;
    x_234 = 'b000011100;
    x_235 = 'b000010110;
    x_236 = 'b000010001;
    x_237 = 'b000011100;
    x_238 = 'b000100011;
    x_239 = 'b000100011;
    x_240 = 'b000011110;
    x_241 = 'b000101001;
    x_242 = 'b000100000;
    x_243 = 'b000011100;
    x_244 = 'b000011110;
    x_245 = 'b000010111;
    x_246 = 'b000011001;
    x_247 = 'b000100001;
    x_248 = 'b000100101;
    x_249 = 'b000100011;
    x_250 = 'b000011000;
    x_251 = 'b000010101;
    x_252 = 'b000101010;
    x_253 = 'b000011111;
    x_254 = 'b000100100;
    x_255 = 'b000010111;

    h_0 = 'b000011100;
    h_1 = 'b000100000;
    h_2 = 'b000011100;
    h_3 = 'b000011010;
    h_4 = 'b000010011;
    h_5 = 'b000001100;
    h_6 = 'b000010010;
    h_7 = 'b000101001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000011010;
    x_1 = 'b000100001;
    x_2 = 'b000011010;
    x_3 = 'b000010111;
    x_4 = 'b000010000;
    x_5 = 'b000001010;
    x_6 = 'b000001110;
    x_7 = 'b000101101;
    x_8 = 'b000100111;
    x_9 = 'b000100011;
    x_10 = 'b000100011;
    x_11 = 'b000011011;
    x_12 = 'b000011010;
    x_13 = 'b000001100;
    x_14 = 'b000110000;
    x_15 = 'b000101000;
    x_16 = 'b000100011;
    x_17 = 'b000011110;
    x_18 = 'b000100010;
    x_19 = 'b000100001;
    x_20 = 'b000100001;
    x_21 = 'b111111011;
    x_22 = 'b111110001;
    x_23 = 'b111110000;
    x_24 = 'b111111110;
    x_25 = 'b000000001;
    x_26 = 'b111111101;
    x_27 = 'b111111111;
    x_28 = 'b111110011;
    x_29 = 'b000001110;
    x_30 = 'b000001011;
    x_31 = 'b000011011;
    x_32 = 'b000010110;
    x_33 = 'b000001101;
    x_34 = 'b000000110;
    x_35 = 'b000000011;
    x_36 = 'b000000000;
    x_37 = 'b111110101;
    x_38 = 'b000101001;
    x_39 = 'b000000101;
    x_40 = 'b000100101;
    x_41 = 'b000001100;
    x_42 = 'b000011111;
    x_43 = 'b000100011;
    x_44 = 'b000010110;
    x_45 = 'b000101011;
    x_46 = 'b000101010;
    x_47 = 'b000101010;
    x_48 = 'b000100100;
    x_49 = 'b000110000;
    x_50 = 'b000101001;
    x_51 = 'b000101000;
    x_52 = 'b000101001;
    x_53 = 'b000100011;
    x_54 = 'b000101000;
    x_55 = 'b000100011;
    x_56 = 'b000101000;
    x_57 = 'b000101010;
    x_58 = 'b000100011;
    x_59 = 'b000100000;
    x_60 = 'b000100000;
    x_61 = 'b000010011;
    x_62 = 'b000011100;
    x_63 = 'b000001101;
    x_64 = 'b000011010;
    x_65 = 'b000100001;
    x_66 = 'b000011010;
    x_67 = 'b000010111;
    x_68 = 'b000010000;
    x_69 = 'b000001010;
    x_70 = 'b000001110;
    x_71 = 'b000101101;
    x_72 = 'b000100111;
    x_73 = 'b000100011;
    x_74 = 'b000100011;
    x_75 = 'b000011011;
    x_76 = 'b000011010;
    x_77 = 'b000001100;
    x_78 = 'b000110000;
    x_79 = 'b000101000;
    x_80 = 'b000100011;
    x_81 = 'b000011110;
    x_82 = 'b000100010;
    x_83 = 'b000100001;
    x_84 = 'b000100001;
    x_85 = 'b111111011;
    x_86 = 'b111110001;
    x_87 = 'b111110000;
    x_88 = 'b111111110;
    x_89 = 'b000000001;
    x_90 = 'b111111101;
    x_91 = 'b111111111;
    x_92 = 'b111110011;
    x_93 = 'b000001110;
    x_94 = 'b000001011;
    x_95 = 'b000011011;
    x_96 = 'b000010110;
    x_97 = 'b000001101;
    x_98 = 'b000000110;
    x_99 = 'b000000011;
    x_100 = 'b000000000;
    x_101 = 'b111110101;
    x_102 = 'b000101001;
    x_103 = 'b000000101;
    x_104 = 'b000100101;
    x_105 = 'b000001100;
    x_106 = 'b000011111;
    x_107 = 'b000100011;
    x_108 = 'b000010110;
    x_109 = 'b000101011;
    x_110 = 'b000101010;
    x_111 = 'b000101010;
    x_112 = 'b000100100;
    x_113 = 'b000110000;
    x_114 = 'b000101001;
    x_115 = 'b000101000;
    x_116 = 'b000101001;
    x_117 = 'b000100011;
    x_118 = 'b000101000;
    x_119 = 'b000100011;
    x_120 = 'b000101000;
    x_121 = 'b000101010;
    x_122 = 'b000100011;
    x_123 = 'b000100000;
    x_124 = 'b000100000;
    x_125 = 'b000010011;
    x_126 = 'b000011100;
    x_127 = 'b000001101;
    x_128 = 'b000011010;
    x_129 = 'b000100001;
    x_130 = 'b000011010;
    x_131 = 'b000010111;
    x_132 = 'b000010000;
    x_133 = 'b000001010;
    x_134 = 'b000001110;
    x_135 = 'b000101101;
    x_136 = 'b000100111;
    x_137 = 'b000100011;
    x_138 = 'b000100011;
    x_139 = 'b000011011;
    x_140 = 'b000011010;
    x_141 = 'b000001100;
    x_142 = 'b000110000;
    x_143 = 'b000101000;
    x_144 = 'b000100011;
    x_145 = 'b000011110;
    x_146 = 'b000100010;
    x_147 = 'b000100001;
    x_148 = 'b000100001;
    x_149 = 'b111111011;
    x_150 = 'b111110001;
    x_151 = 'b111110000;
    x_152 = 'b111111110;
    x_153 = 'b000000001;
    x_154 = 'b111111101;
    x_155 = 'b111111111;
    x_156 = 'b111110011;
    x_157 = 'b000001110;
    x_158 = 'b000001011;
    x_159 = 'b000011011;
    x_160 = 'b000010110;
    x_161 = 'b000001101;
    x_162 = 'b000000110;
    x_163 = 'b000000011;
    x_164 = 'b000000000;
    x_165 = 'b111110101;
    x_166 = 'b000101001;
    x_167 = 'b000000101;
    x_168 = 'b000100101;
    x_169 = 'b000001100;
    x_170 = 'b000011111;
    x_171 = 'b000100011;
    x_172 = 'b000010110;
    x_173 = 'b000101011;
    x_174 = 'b000101010;
    x_175 = 'b000101010;
    x_176 = 'b000100100;
    x_177 = 'b000110000;
    x_178 = 'b000101001;
    x_179 = 'b000101000;
    x_180 = 'b000101001;
    x_181 = 'b000100011;
    x_182 = 'b000101000;
    x_183 = 'b000100011;
    x_184 = 'b000101000;
    x_185 = 'b000101010;
    x_186 = 'b000100011;
    x_187 = 'b000100000;
    x_188 = 'b000100000;
    x_189 = 'b000010011;
    x_190 = 'b000011100;
    x_191 = 'b000001101;
    x_192 = 'b000011010;
    x_193 = 'b000100001;
    x_194 = 'b000011010;
    x_195 = 'b000010111;
    x_196 = 'b000010000;
    x_197 = 'b000001010;
    x_198 = 'b000001110;
    x_199 = 'b000101101;
    x_200 = 'b000100111;
    x_201 = 'b000100011;
    x_202 = 'b000100011;
    x_203 = 'b000011011;
    x_204 = 'b000011010;
    x_205 = 'b000001100;
    x_206 = 'b000110000;
    x_207 = 'b000101000;
    x_208 = 'b000100011;
    x_209 = 'b000011110;
    x_210 = 'b000100010;
    x_211 = 'b000100001;
    x_212 = 'b000100001;
    x_213 = 'b111111011;
    x_214 = 'b111110001;
    x_215 = 'b111110000;
    x_216 = 'b111111110;
    x_217 = 'b000000001;
    x_218 = 'b111111101;
    x_219 = 'b111111111;
    x_220 = 'b111110011;
    x_221 = 'b000001110;
    x_222 = 'b000001011;
    x_223 = 'b000011011;
    x_224 = 'b000010110;
    x_225 = 'b000001101;
    x_226 = 'b000000110;
    x_227 = 'b000000011;
    x_228 = 'b000000000;
    x_229 = 'b111110101;
    x_230 = 'b000101001;
    x_231 = 'b000000101;
    x_232 = 'b000100101;
    x_233 = 'b000001100;
    x_234 = 'b000011111;
    x_235 = 'b000100011;
    x_236 = 'b000010110;
    x_237 = 'b000101011;
    x_238 = 'b000101010;
    x_239 = 'b000101010;
    x_240 = 'b000100100;
    x_241 = 'b000110000;
    x_242 = 'b000101001;
    x_243 = 'b000101000;
    x_244 = 'b000101001;
    x_245 = 'b000100011;
    x_246 = 'b000101000;
    x_247 = 'b000100011;
    x_248 = 'b000101000;
    x_249 = 'b000101010;
    x_250 = 'b000100011;
    x_251 = 'b000100000;
    x_252 = 'b000100000;
    x_253 = 'b000010011;
    x_254 = 'b000011100;
    x_255 = 'b000001101;

    h_0 = 'b000011010;
    h_1 = 'b000100001;
    h_2 = 'b000011010;
    h_3 = 'b000010111;
    h_4 = 'b000010000;
    h_5 = 'b000001010;
    h_6 = 'b000001110;
    h_7 = 'b000101101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000100110;
    x_1 = 'b000101100;
    x_2 = 'b000100011;
    x_3 = 'b000100100;
    x_4 = 'b000011010;
    x_5 = 'b000001110;
    x_6 = 'b000001101;
    x_7 = 'b000110100;
    x_8 = 'b000101101;
    x_9 = 'b000110001;
    x_10 = 'b000110000;
    x_11 = 'b000101011;
    x_12 = 'b000100010;
    x_13 = 'b000010001;
    x_14 = 'b000101011;
    x_15 = 'b000101101;
    x_16 = 'b000101101;
    x_17 = 'b000101010;
    x_18 = 'b000110000;
    x_19 = 'b000101101;
    x_20 = 'b000100111;
    x_21 = 'b111111011;
    x_22 = 'b111110011;
    x_23 = 'b111110011;
    x_24 = 'b111111110;
    x_25 = 'b000000001;
    x_26 = 'b000000010;
    x_27 = 'b000000000;
    x_28 = 'b111110101;
    x_29 = 'b000010111;
    x_30 = 'b000000011;
    x_31 = 'b000011010;
    x_32 = 'b000011000;
    x_33 = 'b000010000;
    x_34 = 'b000001000;
    x_35 = 'b000000010;
    x_36 = 'b111111101;
    x_37 = 'b111101110;
    x_38 = 'b000011011;
    x_39 = 'b000000011;
    x_40 = 'b000001001;
    x_41 = 'b000010100;
    x_42 = 'b000101110;
    x_43 = 'b000100000;
    x_44 = 'b000010010;
    x_45 = 'b000100110;
    x_46 = 'b000100001;
    x_47 = 'b000100010;
    x_48 = 'b000011111;
    x_49 = 'b000101001;
    x_50 = 'b000101000;
    x_51 = 'b000101001;
    x_52 = 'b000101001;
    x_53 = 'b000100001;
    x_54 = 'b000100010;
    x_55 = 'b000011011;
    x_56 = 'b000100100;
    x_57 = 'b000101000;
    x_58 = 'b000100101;
    x_59 = 'b000100001;
    x_60 = 'b000011100;
    x_61 = 'b000010011;
    x_62 = 'b000011110;
    x_63 = 'b000010011;
    x_64 = 'b000100110;
    x_65 = 'b000101100;
    x_66 = 'b000100011;
    x_67 = 'b000100100;
    x_68 = 'b000011010;
    x_69 = 'b000001110;
    x_70 = 'b000001101;
    x_71 = 'b000110100;
    x_72 = 'b000101101;
    x_73 = 'b000110001;
    x_74 = 'b000110000;
    x_75 = 'b000101011;
    x_76 = 'b000100010;
    x_77 = 'b000010001;
    x_78 = 'b000101011;
    x_79 = 'b000101101;
    x_80 = 'b000101101;
    x_81 = 'b000101010;
    x_82 = 'b000110000;
    x_83 = 'b000101101;
    x_84 = 'b000100111;
    x_85 = 'b111111011;
    x_86 = 'b111110011;
    x_87 = 'b111110011;
    x_88 = 'b111111110;
    x_89 = 'b000000001;
    x_90 = 'b000000010;
    x_91 = 'b000000000;
    x_92 = 'b111110101;
    x_93 = 'b000010111;
    x_94 = 'b000000011;
    x_95 = 'b000011010;
    x_96 = 'b000011000;
    x_97 = 'b000010000;
    x_98 = 'b000001000;
    x_99 = 'b000000010;
    x_100 = 'b111111101;
    x_101 = 'b111101110;
    x_102 = 'b000011011;
    x_103 = 'b000000011;
    x_104 = 'b000001001;
    x_105 = 'b000010100;
    x_106 = 'b000101110;
    x_107 = 'b000100000;
    x_108 = 'b000010010;
    x_109 = 'b000100110;
    x_110 = 'b000100001;
    x_111 = 'b000100010;
    x_112 = 'b000011111;
    x_113 = 'b000101001;
    x_114 = 'b000101000;
    x_115 = 'b000101001;
    x_116 = 'b000101001;
    x_117 = 'b000100001;
    x_118 = 'b000100010;
    x_119 = 'b000011011;
    x_120 = 'b000100100;
    x_121 = 'b000101000;
    x_122 = 'b000100101;
    x_123 = 'b000100001;
    x_124 = 'b000011100;
    x_125 = 'b000010011;
    x_126 = 'b000011110;
    x_127 = 'b000010011;
    x_128 = 'b000100110;
    x_129 = 'b000101100;
    x_130 = 'b000100011;
    x_131 = 'b000100100;
    x_132 = 'b000011010;
    x_133 = 'b000001110;
    x_134 = 'b000001101;
    x_135 = 'b000110100;
    x_136 = 'b000101101;
    x_137 = 'b000110001;
    x_138 = 'b000110000;
    x_139 = 'b000101011;
    x_140 = 'b000100010;
    x_141 = 'b000010001;
    x_142 = 'b000101011;
    x_143 = 'b000101101;
    x_144 = 'b000101101;
    x_145 = 'b000101010;
    x_146 = 'b000110000;
    x_147 = 'b000101101;
    x_148 = 'b000100111;
    x_149 = 'b111111011;
    x_150 = 'b111110011;
    x_151 = 'b111110011;
    x_152 = 'b111111110;
    x_153 = 'b000000001;
    x_154 = 'b000000010;
    x_155 = 'b000000000;
    x_156 = 'b111110101;
    x_157 = 'b000010111;
    x_158 = 'b000000011;
    x_159 = 'b000011010;
    x_160 = 'b000011000;
    x_161 = 'b000010000;
    x_162 = 'b000001000;
    x_163 = 'b000000010;
    x_164 = 'b111111101;
    x_165 = 'b111101110;
    x_166 = 'b000011011;
    x_167 = 'b000000011;
    x_168 = 'b000001001;
    x_169 = 'b000010100;
    x_170 = 'b000101110;
    x_171 = 'b000100000;
    x_172 = 'b000010010;
    x_173 = 'b000100110;
    x_174 = 'b000100001;
    x_175 = 'b000100010;
    x_176 = 'b000011111;
    x_177 = 'b000101001;
    x_178 = 'b000101000;
    x_179 = 'b000101001;
    x_180 = 'b000101001;
    x_181 = 'b000100001;
    x_182 = 'b000100010;
    x_183 = 'b000011011;
    x_184 = 'b000100100;
    x_185 = 'b000101000;
    x_186 = 'b000100101;
    x_187 = 'b000100001;
    x_188 = 'b000011100;
    x_189 = 'b000010011;
    x_190 = 'b000011110;
    x_191 = 'b000010011;
    x_192 = 'b000100110;
    x_193 = 'b000101100;
    x_194 = 'b000100011;
    x_195 = 'b000100100;
    x_196 = 'b000011010;
    x_197 = 'b000001110;
    x_198 = 'b000001101;
    x_199 = 'b000110100;
    x_200 = 'b000101101;
    x_201 = 'b000110001;
    x_202 = 'b000110000;
    x_203 = 'b000101011;
    x_204 = 'b000100010;
    x_205 = 'b000010001;
    x_206 = 'b000101011;
    x_207 = 'b000101101;
    x_208 = 'b000101101;
    x_209 = 'b000101010;
    x_210 = 'b000110000;
    x_211 = 'b000101101;
    x_212 = 'b000100111;
    x_213 = 'b111111011;
    x_214 = 'b111110011;
    x_215 = 'b111110011;
    x_216 = 'b111111110;
    x_217 = 'b000000001;
    x_218 = 'b000000010;
    x_219 = 'b000000000;
    x_220 = 'b111110101;
    x_221 = 'b000010111;
    x_222 = 'b000000011;
    x_223 = 'b000011010;
    x_224 = 'b000011000;
    x_225 = 'b000010000;
    x_226 = 'b000001000;
    x_227 = 'b000000010;
    x_228 = 'b111111101;
    x_229 = 'b111101110;
    x_230 = 'b000011011;
    x_231 = 'b000000011;
    x_232 = 'b000001001;
    x_233 = 'b000010100;
    x_234 = 'b000101110;
    x_235 = 'b000100000;
    x_236 = 'b000010010;
    x_237 = 'b000100110;
    x_238 = 'b000100001;
    x_239 = 'b000100010;
    x_240 = 'b000011111;
    x_241 = 'b000101001;
    x_242 = 'b000101000;
    x_243 = 'b000101001;
    x_244 = 'b000101001;
    x_245 = 'b000100001;
    x_246 = 'b000100010;
    x_247 = 'b000011011;
    x_248 = 'b000100100;
    x_249 = 'b000101000;
    x_250 = 'b000100101;
    x_251 = 'b000100001;
    x_252 = 'b000011100;
    x_253 = 'b000010011;
    x_254 = 'b000011110;
    x_255 = 'b000010011;

    h_0 = 'b000100110;
    h_1 = 'b000101100;
    h_2 = 'b000100011;
    h_3 = 'b000100100;
    h_4 = 'b000011010;
    h_5 = 'b000001110;
    h_6 = 'b000001101;
    h_7 = 'b000110100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000010101;
    x_1 = 'b000011100;
    x_2 = 'b000011001;
    x_3 = 'b000100000;
    x_4 = 'b000011001;
    x_5 = 'b000001100;
    x_6 = 'b000001111;
    x_7 = 'b000010111;
    x_8 = 'b000100000;
    x_9 = 'b000100100;
    x_10 = 'b000100110;
    x_11 = 'b000100010;
    x_12 = 'b000100001;
    x_13 = 'b000010000;
    x_14 = 'b000011101;
    x_15 = 'b000100010;
    x_16 = 'b000100100;
    x_17 = 'b000100001;
    x_18 = 'b000101011;
    x_19 = 'b000101000;
    x_20 = 'b000100011;
    x_21 = 'b111111010;
    x_22 = 'b111110010;
    x_23 = 'b111110011;
    x_24 = 'b111111100;
    x_25 = 'b111111110;
    x_26 = 'b111111111;
    x_27 = 'b000000000;
    x_28 = 'b111110100;
    x_29 = 'b000010011;
    x_30 = 'b111111111;
    x_31 = 'b000011001;
    x_32 = 'b000010000;
    x_33 = 'b000001011;
    x_34 = 'b000000110;
    x_35 = 'b111111111;
    x_36 = 'b111111111;
    x_37 = 'b111110100;
    x_38 = 'b000010111;
    x_39 = 'b000001000;
    x_40 = 'b000011100;
    x_41 = 'b000100000;
    x_42 = 'b000110001;
    x_43 = 'b111110101;
    x_44 = 'b000011010;
    x_45 = 'b000100111;
    x_46 = 'b000011011;
    x_47 = 'b000100010;
    x_48 = 'b000011111;
    x_49 = 'b000101010;
    x_50 = 'b000101001;
    x_51 = 'b000101111;
    x_52 = 'b000101101;
    x_53 = 'b000100111;
    x_54 = 'b000101000;
    x_55 = 'b000011101;
    x_56 = 'b000100111;
    x_57 = 'b000110000;
    x_58 = 'b000110000;
    x_59 = 'b000101101;
    x_60 = 'b000011110;
    x_61 = 'b000011101;
    x_62 = 'b000101011;
    x_63 = 'b000100011;
    x_64 = 'b000010101;
    x_65 = 'b000011100;
    x_66 = 'b000011001;
    x_67 = 'b000100000;
    x_68 = 'b000011001;
    x_69 = 'b000001100;
    x_70 = 'b000001111;
    x_71 = 'b000010111;
    x_72 = 'b000100000;
    x_73 = 'b000100100;
    x_74 = 'b000100110;
    x_75 = 'b000100010;
    x_76 = 'b000100001;
    x_77 = 'b000010000;
    x_78 = 'b000011101;
    x_79 = 'b000100010;
    x_80 = 'b000100100;
    x_81 = 'b000100001;
    x_82 = 'b000101011;
    x_83 = 'b000101000;
    x_84 = 'b000100011;
    x_85 = 'b111111010;
    x_86 = 'b111110010;
    x_87 = 'b111110011;
    x_88 = 'b111111100;
    x_89 = 'b111111110;
    x_90 = 'b111111111;
    x_91 = 'b000000000;
    x_92 = 'b111110100;
    x_93 = 'b000010011;
    x_94 = 'b111111111;
    x_95 = 'b000011001;
    x_96 = 'b000010000;
    x_97 = 'b000001011;
    x_98 = 'b000000110;
    x_99 = 'b111111111;
    x_100 = 'b111111111;
    x_101 = 'b111110100;
    x_102 = 'b000010111;
    x_103 = 'b000001000;
    x_104 = 'b000011100;
    x_105 = 'b000100000;
    x_106 = 'b000110001;
    x_107 = 'b111110101;
    x_108 = 'b000011010;
    x_109 = 'b000100111;
    x_110 = 'b000011011;
    x_111 = 'b000100010;
    x_112 = 'b000011111;
    x_113 = 'b000101010;
    x_114 = 'b000101001;
    x_115 = 'b000101111;
    x_116 = 'b000101101;
    x_117 = 'b000100111;
    x_118 = 'b000101000;
    x_119 = 'b000011101;
    x_120 = 'b000100111;
    x_121 = 'b000110000;
    x_122 = 'b000110000;
    x_123 = 'b000101101;
    x_124 = 'b000011110;
    x_125 = 'b000011101;
    x_126 = 'b000101011;
    x_127 = 'b000100011;
    x_128 = 'b000010101;
    x_129 = 'b000011100;
    x_130 = 'b000011001;
    x_131 = 'b000100000;
    x_132 = 'b000011001;
    x_133 = 'b000001100;
    x_134 = 'b000001111;
    x_135 = 'b000010111;
    x_136 = 'b000100000;
    x_137 = 'b000100100;
    x_138 = 'b000100110;
    x_139 = 'b000100010;
    x_140 = 'b000100001;
    x_141 = 'b000010000;
    x_142 = 'b000011101;
    x_143 = 'b000100010;
    x_144 = 'b000100100;
    x_145 = 'b000100001;
    x_146 = 'b000101011;
    x_147 = 'b000101000;
    x_148 = 'b000100011;
    x_149 = 'b111111010;
    x_150 = 'b111110010;
    x_151 = 'b111110011;
    x_152 = 'b111111100;
    x_153 = 'b111111110;
    x_154 = 'b111111111;
    x_155 = 'b000000000;
    x_156 = 'b111110100;
    x_157 = 'b000010011;
    x_158 = 'b111111111;
    x_159 = 'b000011001;
    x_160 = 'b000010000;
    x_161 = 'b000001011;
    x_162 = 'b000000110;
    x_163 = 'b111111111;
    x_164 = 'b111111111;
    x_165 = 'b111110100;
    x_166 = 'b000010111;
    x_167 = 'b000001000;
    x_168 = 'b000011100;
    x_169 = 'b000100000;
    x_170 = 'b000110001;
    x_171 = 'b111110101;
    x_172 = 'b000011010;
    x_173 = 'b000100111;
    x_174 = 'b000011011;
    x_175 = 'b000100010;
    x_176 = 'b000011111;
    x_177 = 'b000101010;
    x_178 = 'b000101001;
    x_179 = 'b000101111;
    x_180 = 'b000101101;
    x_181 = 'b000100111;
    x_182 = 'b000101000;
    x_183 = 'b000011101;
    x_184 = 'b000100111;
    x_185 = 'b000110000;
    x_186 = 'b000110000;
    x_187 = 'b000101101;
    x_188 = 'b000011110;
    x_189 = 'b000011101;
    x_190 = 'b000101011;
    x_191 = 'b000100011;
    x_192 = 'b000010101;
    x_193 = 'b000011100;
    x_194 = 'b000011001;
    x_195 = 'b000100000;
    x_196 = 'b000011001;
    x_197 = 'b000001100;
    x_198 = 'b000001111;
    x_199 = 'b000010111;
    x_200 = 'b000100000;
    x_201 = 'b000100100;
    x_202 = 'b000100110;
    x_203 = 'b000100010;
    x_204 = 'b000100001;
    x_205 = 'b000010000;
    x_206 = 'b000011101;
    x_207 = 'b000100010;
    x_208 = 'b000100100;
    x_209 = 'b000100001;
    x_210 = 'b000101011;
    x_211 = 'b000101000;
    x_212 = 'b000100011;
    x_213 = 'b111111010;
    x_214 = 'b111110010;
    x_215 = 'b111110011;
    x_216 = 'b111111100;
    x_217 = 'b111111110;
    x_218 = 'b111111111;
    x_219 = 'b000000000;
    x_220 = 'b111110100;
    x_221 = 'b000010011;
    x_222 = 'b111111111;
    x_223 = 'b000011001;
    x_224 = 'b000010000;
    x_225 = 'b000001011;
    x_226 = 'b000000110;
    x_227 = 'b111111111;
    x_228 = 'b111111111;
    x_229 = 'b111110100;
    x_230 = 'b000010111;
    x_231 = 'b000001000;
    x_232 = 'b000011100;
    x_233 = 'b000100000;
    x_234 = 'b000110001;
    x_235 = 'b111110101;
    x_236 = 'b000011010;
    x_237 = 'b000100111;
    x_238 = 'b000011011;
    x_239 = 'b000100010;
    x_240 = 'b000011111;
    x_241 = 'b000101010;
    x_242 = 'b000101001;
    x_243 = 'b000101111;
    x_244 = 'b000101101;
    x_245 = 'b000100111;
    x_246 = 'b000101000;
    x_247 = 'b000011101;
    x_248 = 'b000100111;
    x_249 = 'b000110000;
    x_250 = 'b000110000;
    x_251 = 'b000101101;
    x_252 = 'b000011110;
    x_253 = 'b000011101;
    x_254 = 'b000101011;
    x_255 = 'b000100011;

    h_0 = 'b000010101;
    h_1 = 'b000011100;
    h_2 = 'b000011001;
    h_3 = 'b000100000;
    h_4 = 'b000011001;
    h_5 = 'b000001100;
    h_6 = 'b000001111;
    h_7 = 'b000010111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111100111;
    x_1 = 'b111011000;
    x_2 = 'b111000111;
    x_3 = 'b110111000;
    x_4 = 'b110111100;
    x_5 = 'b110111000;
    x_6 = 'b111000110;
    x_7 = 'b111101111;
    x_8 = 'b111000110;
    x_9 = 'b111000010;
    x_10 = 'b110111101;
    x_11 = 'b110110101;
    x_12 = 'b111000000;
    x_13 = 'b110110111;
    x_14 = 'b111010010;
    x_15 = 'b111001100;
    x_16 = 'b111000100;
    x_17 = 'b111000000;
    x_18 = 'b111001011;
    x_19 = 'b111001111;
    x_20 = 'b111001011;
    x_21 = 'b111101011;
    x_22 = 'b111011010;
    x_23 = 'b111011001;
    x_24 = 'b111111001;
    x_25 = 'b111110111;
    x_26 = 'b111000010;
    x_27 = 'b110111111;
    x_28 = 'b111010100;
    x_29 = 'b111101110;
    x_30 = 'b111100101;
    x_31 = 'b110111101;
    x_32 = 'b111000001;
    x_33 = 'b110111001;
    x_34 = 'b110110110;
    x_35 = 'b111000000;
    x_36 = 'b110111010;
    x_37 = 'b111101000;
    x_38 = 'b111011110;
    x_39 = 'b110110101;
    x_40 = 'b111001101;
    x_41 = 'b110110110;
    x_42 = 'b111010110;
    x_43 = 'b111100011;
    x_44 = 'b111011010;
    x_45 = 'b111100001;
    x_46 = 'b111011001;
    x_47 = 'b111010101;
    x_48 = 'b111010010;
    x_49 = 'b111001111;
    x_50 = 'b111001001;
    x_51 = 'b111011010;
    x_52 = 'b111100000;
    x_53 = 'b111101010;
    x_54 = 'b111100000;
    x_55 = 'b111110100;
    x_56 = 'b111100010;
    x_57 = 'b111100101;
    x_58 = 'b111110010;
    x_59 = 'b111110100;
    x_60 = 'b000000111;
    x_61 = 'b111110110;
    x_62 = 'b000000100;
    x_63 = 'b000001001;
    x_64 = 'b111100111;
    x_65 = 'b111011000;
    x_66 = 'b111000111;
    x_67 = 'b110111000;
    x_68 = 'b110111100;
    x_69 = 'b110111000;
    x_70 = 'b111000110;
    x_71 = 'b111101111;
    x_72 = 'b111000110;
    x_73 = 'b111000010;
    x_74 = 'b110111101;
    x_75 = 'b110110101;
    x_76 = 'b111000000;
    x_77 = 'b110110111;
    x_78 = 'b111010010;
    x_79 = 'b111001100;
    x_80 = 'b111000100;
    x_81 = 'b111000000;
    x_82 = 'b111001011;
    x_83 = 'b111001111;
    x_84 = 'b111001011;
    x_85 = 'b111101011;
    x_86 = 'b111011010;
    x_87 = 'b111011001;
    x_88 = 'b111111001;
    x_89 = 'b111110111;
    x_90 = 'b111000010;
    x_91 = 'b110111111;
    x_92 = 'b111010100;
    x_93 = 'b111101110;
    x_94 = 'b111100101;
    x_95 = 'b110111101;
    x_96 = 'b111000001;
    x_97 = 'b110111001;
    x_98 = 'b110110110;
    x_99 = 'b111000000;
    x_100 = 'b110111010;
    x_101 = 'b111101000;
    x_102 = 'b111011110;
    x_103 = 'b110110101;
    x_104 = 'b111001101;
    x_105 = 'b110110110;
    x_106 = 'b111010110;
    x_107 = 'b111100011;
    x_108 = 'b111011010;
    x_109 = 'b111100001;
    x_110 = 'b111011001;
    x_111 = 'b111010101;
    x_112 = 'b111010010;
    x_113 = 'b111001111;
    x_114 = 'b111001001;
    x_115 = 'b111011010;
    x_116 = 'b111100000;
    x_117 = 'b111101010;
    x_118 = 'b111100000;
    x_119 = 'b111110100;
    x_120 = 'b111100010;
    x_121 = 'b111100101;
    x_122 = 'b111110010;
    x_123 = 'b111110100;
    x_124 = 'b000000111;
    x_125 = 'b111110110;
    x_126 = 'b000000100;
    x_127 = 'b000001001;
    x_128 = 'b111100111;
    x_129 = 'b111011000;
    x_130 = 'b111000111;
    x_131 = 'b110111000;
    x_132 = 'b110111100;
    x_133 = 'b110111000;
    x_134 = 'b111000110;
    x_135 = 'b111101111;
    x_136 = 'b111000110;
    x_137 = 'b111000010;
    x_138 = 'b110111101;
    x_139 = 'b110110101;
    x_140 = 'b111000000;
    x_141 = 'b110110111;
    x_142 = 'b111010010;
    x_143 = 'b111001100;
    x_144 = 'b111000100;
    x_145 = 'b111000000;
    x_146 = 'b111001011;
    x_147 = 'b111001111;
    x_148 = 'b111001011;
    x_149 = 'b111101011;
    x_150 = 'b111011010;
    x_151 = 'b111011001;
    x_152 = 'b111111001;
    x_153 = 'b111110111;
    x_154 = 'b111000010;
    x_155 = 'b110111111;
    x_156 = 'b111010100;
    x_157 = 'b111101110;
    x_158 = 'b111100101;
    x_159 = 'b110111101;
    x_160 = 'b111000001;
    x_161 = 'b110111001;
    x_162 = 'b110110110;
    x_163 = 'b111000000;
    x_164 = 'b110111010;
    x_165 = 'b111101000;
    x_166 = 'b111011110;
    x_167 = 'b110110101;
    x_168 = 'b111001101;
    x_169 = 'b110110110;
    x_170 = 'b111010110;
    x_171 = 'b111100011;
    x_172 = 'b111011010;
    x_173 = 'b111100001;
    x_174 = 'b111011001;
    x_175 = 'b111010101;
    x_176 = 'b111010010;
    x_177 = 'b111001111;
    x_178 = 'b111001001;
    x_179 = 'b111011010;
    x_180 = 'b111100000;
    x_181 = 'b111101010;
    x_182 = 'b111100000;
    x_183 = 'b111110100;
    x_184 = 'b111100010;
    x_185 = 'b111100101;
    x_186 = 'b111110010;
    x_187 = 'b111110100;
    x_188 = 'b000000111;
    x_189 = 'b111110110;
    x_190 = 'b000000100;
    x_191 = 'b000001001;
    x_192 = 'b111100111;
    x_193 = 'b111011000;
    x_194 = 'b111000111;
    x_195 = 'b110111000;
    x_196 = 'b110111100;
    x_197 = 'b110111000;
    x_198 = 'b111000110;
    x_199 = 'b111101111;
    x_200 = 'b111000110;
    x_201 = 'b111000010;
    x_202 = 'b110111101;
    x_203 = 'b110110101;
    x_204 = 'b111000000;
    x_205 = 'b110110111;
    x_206 = 'b111010010;
    x_207 = 'b111001100;
    x_208 = 'b111000100;
    x_209 = 'b111000000;
    x_210 = 'b111001011;
    x_211 = 'b111001111;
    x_212 = 'b111001011;
    x_213 = 'b111101011;
    x_214 = 'b111011010;
    x_215 = 'b111011001;
    x_216 = 'b111111001;
    x_217 = 'b111110111;
    x_218 = 'b111000010;
    x_219 = 'b110111111;
    x_220 = 'b111010100;
    x_221 = 'b111101110;
    x_222 = 'b111100101;
    x_223 = 'b110111101;
    x_224 = 'b111000001;
    x_225 = 'b110111001;
    x_226 = 'b110110110;
    x_227 = 'b111000000;
    x_228 = 'b110111010;
    x_229 = 'b111101000;
    x_230 = 'b111011110;
    x_231 = 'b110110101;
    x_232 = 'b111001101;
    x_233 = 'b110110110;
    x_234 = 'b111010110;
    x_235 = 'b111100011;
    x_236 = 'b111011010;
    x_237 = 'b111100001;
    x_238 = 'b111011001;
    x_239 = 'b111010101;
    x_240 = 'b111010010;
    x_241 = 'b111001111;
    x_242 = 'b111001001;
    x_243 = 'b111011010;
    x_244 = 'b111100000;
    x_245 = 'b111101010;
    x_246 = 'b111100000;
    x_247 = 'b111110100;
    x_248 = 'b111100010;
    x_249 = 'b111100101;
    x_250 = 'b111110010;
    x_251 = 'b111110100;
    x_252 = 'b000000111;
    x_253 = 'b111110110;
    x_254 = 'b000000100;
    x_255 = 'b000001001;

    h_0 = 'b111100111;
    h_1 = 'b111011000;
    h_2 = 'b111000111;
    h_3 = 'b110111000;
    h_4 = 'b110111100;
    h_5 = 'b110111000;
    h_6 = 'b111000110;
    h_7 = 'b111101111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111010111;
    x_1 = 'b111001010;
    x_2 = 'b110110101;
    x_3 = 'b110100100;
    x_4 = 'b110100100;
    x_5 = 'b110011100;
    x_6 = 'b110110011;
    x_7 = 'b111100000;
    x_8 = 'b110111001;
    x_9 = 'b110110100;
    x_10 = 'b110101110;
    x_11 = 'b110101001;
    x_12 = 'b110101001;
    x_13 = 'b110101011;
    x_14 = 'b111001001;
    x_15 = 'b111000001;
    x_16 = 'b110111010;
    x_17 = 'b110110110;
    x_18 = 'b110111110;
    x_19 = 'b110111111;
    x_20 = 'b110111110;
    x_21 = 'b111100110;
    x_22 = 'b111010111;
    x_23 = 'b111010111;
    x_24 = 'b111110111;
    x_25 = 'b111110110;
    x_26 = 'b110111001;
    x_27 = 'b110110111;
    x_28 = 'b111010010;
    x_29 = 'b111101110;
    x_30 = 'b111100100;
    x_31 = 'b110110011;
    x_32 = 'b110111000;
    x_33 = 'b110101110;
    x_34 = 'b110101011;
    x_35 = 'b110110101;
    x_36 = 'b110110000;
    x_37 = 'b111100101;
    x_38 = 'b111100000;
    x_39 = 'b110110001;
    x_40 = 'b111010001;
    x_41 = 'b110101000;
    x_42 = 'b111101110;
    x_43 = 'b111000011;
    x_44 = 'b111100100;
    x_45 = 'b111011101;
    x_46 = 'b111100010;
    x_47 = 'b111011001;
    x_48 = 'b111010101;
    x_49 = 'b111010101;
    x_50 = 'b111001111;
    x_51 = 'b111011111;
    x_52 = 'b111100010;
    x_53 = 'b111101010;
    x_54 = 'b111100011;
    x_55 = 'b111110111;
    x_56 = 'b111100110;
    x_57 = 'b111110000;
    x_58 = 'b111110011;
    x_59 = 'b111110010;
    x_60 = 'b111111100;
    x_61 = 'b111101111;
    x_62 = 'b111111001;
    x_63 = 'b111110011;
    x_64 = 'b111010111;
    x_65 = 'b111001010;
    x_66 = 'b110110101;
    x_67 = 'b110100100;
    x_68 = 'b110100100;
    x_69 = 'b110011100;
    x_70 = 'b110110011;
    x_71 = 'b111100000;
    x_72 = 'b110111001;
    x_73 = 'b110110100;
    x_74 = 'b110101110;
    x_75 = 'b110101001;
    x_76 = 'b110101001;
    x_77 = 'b110101011;
    x_78 = 'b111001001;
    x_79 = 'b111000001;
    x_80 = 'b110111010;
    x_81 = 'b110110110;
    x_82 = 'b110111110;
    x_83 = 'b110111111;
    x_84 = 'b110111110;
    x_85 = 'b111100110;
    x_86 = 'b111010111;
    x_87 = 'b111010111;
    x_88 = 'b111110111;
    x_89 = 'b111110110;
    x_90 = 'b110111001;
    x_91 = 'b110110111;
    x_92 = 'b111010010;
    x_93 = 'b111101110;
    x_94 = 'b111100100;
    x_95 = 'b110110011;
    x_96 = 'b110111000;
    x_97 = 'b110101110;
    x_98 = 'b110101011;
    x_99 = 'b110110101;
    x_100 = 'b110110000;
    x_101 = 'b111100101;
    x_102 = 'b111100000;
    x_103 = 'b110110001;
    x_104 = 'b111010001;
    x_105 = 'b110101000;
    x_106 = 'b111101110;
    x_107 = 'b111000011;
    x_108 = 'b111100100;
    x_109 = 'b111011101;
    x_110 = 'b111100010;
    x_111 = 'b111011001;
    x_112 = 'b111010101;
    x_113 = 'b111010101;
    x_114 = 'b111001111;
    x_115 = 'b111011111;
    x_116 = 'b111100010;
    x_117 = 'b111101010;
    x_118 = 'b111100011;
    x_119 = 'b111110111;
    x_120 = 'b111100110;
    x_121 = 'b111110000;
    x_122 = 'b111110011;
    x_123 = 'b111110010;
    x_124 = 'b111111100;
    x_125 = 'b111101111;
    x_126 = 'b111111001;
    x_127 = 'b111110011;
    x_128 = 'b111010111;
    x_129 = 'b111001010;
    x_130 = 'b110110101;
    x_131 = 'b110100100;
    x_132 = 'b110100100;
    x_133 = 'b110011100;
    x_134 = 'b110110011;
    x_135 = 'b111100000;
    x_136 = 'b110111001;
    x_137 = 'b110110100;
    x_138 = 'b110101110;
    x_139 = 'b110101001;
    x_140 = 'b110101001;
    x_141 = 'b110101011;
    x_142 = 'b111001001;
    x_143 = 'b111000001;
    x_144 = 'b110111010;
    x_145 = 'b110110110;
    x_146 = 'b110111110;
    x_147 = 'b110111111;
    x_148 = 'b110111110;
    x_149 = 'b111100110;
    x_150 = 'b111010111;
    x_151 = 'b111010111;
    x_152 = 'b111110111;
    x_153 = 'b111110110;
    x_154 = 'b110111001;
    x_155 = 'b110110111;
    x_156 = 'b111010010;
    x_157 = 'b111101110;
    x_158 = 'b111100100;
    x_159 = 'b110110011;
    x_160 = 'b110111000;
    x_161 = 'b110101110;
    x_162 = 'b110101011;
    x_163 = 'b110110101;
    x_164 = 'b110110000;
    x_165 = 'b111100101;
    x_166 = 'b111100000;
    x_167 = 'b110110001;
    x_168 = 'b111010001;
    x_169 = 'b110101000;
    x_170 = 'b111101110;
    x_171 = 'b111000011;
    x_172 = 'b111100100;
    x_173 = 'b111011101;
    x_174 = 'b111100010;
    x_175 = 'b111011001;
    x_176 = 'b111010101;
    x_177 = 'b111010101;
    x_178 = 'b111001111;
    x_179 = 'b111011111;
    x_180 = 'b111100010;
    x_181 = 'b111101010;
    x_182 = 'b111100011;
    x_183 = 'b111110111;
    x_184 = 'b111100110;
    x_185 = 'b111110000;
    x_186 = 'b111110011;
    x_187 = 'b111110010;
    x_188 = 'b111111100;
    x_189 = 'b111101111;
    x_190 = 'b111111001;
    x_191 = 'b111110011;
    x_192 = 'b111010111;
    x_193 = 'b111001010;
    x_194 = 'b110110101;
    x_195 = 'b110100100;
    x_196 = 'b110100100;
    x_197 = 'b110011100;
    x_198 = 'b110110011;
    x_199 = 'b111100000;
    x_200 = 'b110111001;
    x_201 = 'b110110100;
    x_202 = 'b110101110;
    x_203 = 'b110101001;
    x_204 = 'b110101001;
    x_205 = 'b110101011;
    x_206 = 'b111001001;
    x_207 = 'b111000001;
    x_208 = 'b110111010;
    x_209 = 'b110110110;
    x_210 = 'b110111110;
    x_211 = 'b110111111;
    x_212 = 'b110111110;
    x_213 = 'b111100110;
    x_214 = 'b111010111;
    x_215 = 'b111010111;
    x_216 = 'b111110111;
    x_217 = 'b111110110;
    x_218 = 'b110111001;
    x_219 = 'b110110111;
    x_220 = 'b111010010;
    x_221 = 'b111101110;
    x_222 = 'b111100100;
    x_223 = 'b110110011;
    x_224 = 'b110111000;
    x_225 = 'b110101110;
    x_226 = 'b110101011;
    x_227 = 'b110110101;
    x_228 = 'b110110000;
    x_229 = 'b111100101;
    x_230 = 'b111100000;
    x_231 = 'b110110001;
    x_232 = 'b111010001;
    x_233 = 'b110101000;
    x_234 = 'b111101110;
    x_235 = 'b111000011;
    x_236 = 'b111100100;
    x_237 = 'b111011101;
    x_238 = 'b111100010;
    x_239 = 'b111011001;
    x_240 = 'b111010101;
    x_241 = 'b111010101;
    x_242 = 'b111001111;
    x_243 = 'b111011111;
    x_244 = 'b111100010;
    x_245 = 'b111101010;
    x_246 = 'b111100011;
    x_247 = 'b111110111;
    x_248 = 'b111100110;
    x_249 = 'b111110000;
    x_250 = 'b111110011;
    x_251 = 'b111110010;
    x_252 = 'b111111100;
    x_253 = 'b111101111;
    x_254 = 'b111111001;
    x_255 = 'b111110011;

    h_0 = 'b111010111;
    h_1 = 'b111001010;
    h_2 = 'b110110101;
    h_3 = 'b110100100;
    h_4 = 'b110100100;
    h_5 = 'b110011100;
    h_6 = 'b110110011;
    h_7 = 'b111100000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111011001;
    x_1 = 'b111001001;
    x_2 = 'b110111001;
    x_3 = 'b110101010;
    x_4 = 'b110101001;
    x_5 = 'b110100110;
    x_6 = 'b110111010;
    x_7 = 'b111100101;
    x_8 = 'b111000100;
    x_9 = 'b110111111;
    x_10 = 'b110111100;
    x_11 = 'b110110111;
    x_12 = 'b110110000;
    x_13 = 'b110110010;
    x_14 = 'b111011000;
    x_15 = 'b111001111;
    x_16 = 'b111001010;
    x_17 = 'b111000110;
    x_18 = 'b111001100;
    x_19 = 'b111001011;
    x_20 = 'b111000101;
    x_21 = 'b111101010;
    x_22 = 'b111011011;
    x_23 = 'b111011011;
    x_24 = 'b111111100;
    x_25 = 'b111111011;
    x_26 = 'b111000010;
    x_27 = 'b110111111;
    x_28 = 'b111010101;
    x_29 = 'b111110110;
    x_30 = 'b111101101;
    x_31 = 'b111000001;
    x_32 = 'b111000100;
    x_33 = 'b110111001;
    x_34 = 'b110111000;
    x_35 = 'b111000011;
    x_36 = 'b110111101;
    x_37 = 'b111110011;
    x_38 = 'b111110011;
    x_39 = 'b111000111;
    x_40 = 'b111110111;
    x_41 = 'b111000001;
    x_42 = 'b111110101;
    x_43 = 'b111001101;
    x_44 = 'b111110111;
    x_45 = 'b111110100;
    x_46 = 'b111110010;
    x_47 = 'b111101010;
    x_48 = 'b111100111;
    x_49 = 'b111101010;
    x_50 = 'b111100111;
    x_51 = 'b111110010;
    x_52 = 'b111110010;
    x_53 = 'b111110111;
    x_54 = 'b111110010;
    x_55 = 'b111111010;
    x_56 = 'b111101110;
    x_57 = 'b000000000;
    x_58 = 'b111111101;
    x_59 = 'b111110101;
    x_60 = 'b111111000;
    x_61 = 'b111110001;
    x_62 = 'b111111001;
    x_63 = 'b111101111;
    x_64 = 'b111011001;
    x_65 = 'b111001001;
    x_66 = 'b110111001;
    x_67 = 'b110101010;
    x_68 = 'b110101001;
    x_69 = 'b110100110;
    x_70 = 'b110111010;
    x_71 = 'b111100101;
    x_72 = 'b111000100;
    x_73 = 'b110111111;
    x_74 = 'b110111100;
    x_75 = 'b110110111;
    x_76 = 'b110110000;
    x_77 = 'b110110010;
    x_78 = 'b111011000;
    x_79 = 'b111001111;
    x_80 = 'b111001010;
    x_81 = 'b111000110;
    x_82 = 'b111001100;
    x_83 = 'b111001011;
    x_84 = 'b111000101;
    x_85 = 'b111101010;
    x_86 = 'b111011011;
    x_87 = 'b111011011;
    x_88 = 'b111111100;
    x_89 = 'b111111011;
    x_90 = 'b111000010;
    x_91 = 'b110111111;
    x_92 = 'b111010101;
    x_93 = 'b111110110;
    x_94 = 'b111101101;
    x_95 = 'b111000001;
    x_96 = 'b111000100;
    x_97 = 'b110111001;
    x_98 = 'b110111000;
    x_99 = 'b111000011;
    x_100 = 'b110111101;
    x_101 = 'b111110011;
    x_102 = 'b111110011;
    x_103 = 'b111000111;
    x_104 = 'b111110111;
    x_105 = 'b111000001;
    x_106 = 'b111110101;
    x_107 = 'b111001101;
    x_108 = 'b111110111;
    x_109 = 'b111110100;
    x_110 = 'b111110010;
    x_111 = 'b111101010;
    x_112 = 'b111100111;
    x_113 = 'b111101010;
    x_114 = 'b111100111;
    x_115 = 'b111110010;
    x_116 = 'b111110010;
    x_117 = 'b111110111;
    x_118 = 'b111110010;
    x_119 = 'b111111010;
    x_120 = 'b111101110;
    x_121 = 'b000000000;
    x_122 = 'b111111101;
    x_123 = 'b111110101;
    x_124 = 'b111111000;
    x_125 = 'b111110001;
    x_126 = 'b111111001;
    x_127 = 'b111101111;
    x_128 = 'b111011001;
    x_129 = 'b111001001;
    x_130 = 'b110111001;
    x_131 = 'b110101010;
    x_132 = 'b110101001;
    x_133 = 'b110100110;
    x_134 = 'b110111010;
    x_135 = 'b111100101;
    x_136 = 'b111000100;
    x_137 = 'b110111111;
    x_138 = 'b110111100;
    x_139 = 'b110110111;
    x_140 = 'b110110000;
    x_141 = 'b110110010;
    x_142 = 'b111011000;
    x_143 = 'b111001111;
    x_144 = 'b111001010;
    x_145 = 'b111000110;
    x_146 = 'b111001100;
    x_147 = 'b111001011;
    x_148 = 'b111000101;
    x_149 = 'b111101010;
    x_150 = 'b111011011;
    x_151 = 'b111011011;
    x_152 = 'b111111100;
    x_153 = 'b111111011;
    x_154 = 'b111000010;
    x_155 = 'b110111111;
    x_156 = 'b111010101;
    x_157 = 'b111110110;
    x_158 = 'b111101101;
    x_159 = 'b111000001;
    x_160 = 'b111000100;
    x_161 = 'b110111001;
    x_162 = 'b110111000;
    x_163 = 'b111000011;
    x_164 = 'b110111101;
    x_165 = 'b111110011;
    x_166 = 'b111110011;
    x_167 = 'b111000111;
    x_168 = 'b111110111;
    x_169 = 'b111000001;
    x_170 = 'b111110101;
    x_171 = 'b111001101;
    x_172 = 'b111110111;
    x_173 = 'b111110100;
    x_174 = 'b111110010;
    x_175 = 'b111101010;
    x_176 = 'b111100111;
    x_177 = 'b111101010;
    x_178 = 'b111100111;
    x_179 = 'b111110010;
    x_180 = 'b111110010;
    x_181 = 'b111110111;
    x_182 = 'b111110010;
    x_183 = 'b111111010;
    x_184 = 'b111101110;
    x_185 = 'b000000000;
    x_186 = 'b111111101;
    x_187 = 'b111110101;
    x_188 = 'b111111000;
    x_189 = 'b111110001;
    x_190 = 'b111111001;
    x_191 = 'b111101111;
    x_192 = 'b111011001;
    x_193 = 'b111001001;
    x_194 = 'b110111001;
    x_195 = 'b110101010;
    x_196 = 'b110101001;
    x_197 = 'b110100110;
    x_198 = 'b110111010;
    x_199 = 'b111100101;
    x_200 = 'b111000100;
    x_201 = 'b110111111;
    x_202 = 'b110111100;
    x_203 = 'b110110111;
    x_204 = 'b110110000;
    x_205 = 'b110110010;
    x_206 = 'b111011000;
    x_207 = 'b111001111;
    x_208 = 'b111001010;
    x_209 = 'b111000110;
    x_210 = 'b111001100;
    x_211 = 'b111001011;
    x_212 = 'b111000101;
    x_213 = 'b111101010;
    x_214 = 'b111011011;
    x_215 = 'b111011011;
    x_216 = 'b111111100;
    x_217 = 'b111111011;
    x_218 = 'b111000010;
    x_219 = 'b110111111;
    x_220 = 'b111010101;
    x_221 = 'b111110110;
    x_222 = 'b111101101;
    x_223 = 'b111000001;
    x_224 = 'b111000100;
    x_225 = 'b110111001;
    x_226 = 'b110111000;
    x_227 = 'b111000011;
    x_228 = 'b110111101;
    x_229 = 'b111110011;
    x_230 = 'b111110011;
    x_231 = 'b111000111;
    x_232 = 'b111110111;
    x_233 = 'b111000001;
    x_234 = 'b111110101;
    x_235 = 'b111001101;
    x_236 = 'b111110111;
    x_237 = 'b111110100;
    x_238 = 'b111110010;
    x_239 = 'b111101010;
    x_240 = 'b111100111;
    x_241 = 'b111101010;
    x_242 = 'b111100111;
    x_243 = 'b111110010;
    x_244 = 'b111110010;
    x_245 = 'b111110111;
    x_246 = 'b111110010;
    x_247 = 'b111111010;
    x_248 = 'b111101110;
    x_249 = 'b000000000;
    x_250 = 'b111111101;
    x_251 = 'b111110101;
    x_252 = 'b111111000;
    x_253 = 'b111110001;
    x_254 = 'b111111001;
    x_255 = 'b111101111;

    h_0 = 'b111011001;
    h_1 = 'b111001001;
    h_2 = 'b110111001;
    h_3 = 'b110101010;
    h_4 = 'b110101001;
    h_5 = 'b110100110;
    h_6 = 'b110111010;
    h_7 = 'b111100101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111101101;
    x_1 = 'b111100001;
    x_2 = 'b111010000;
    x_3 = 'b111000000;
    x_4 = 'b111000000;
    x_5 = 'b110111110;
    x_6 = 'b111010110;
    x_7 = 'b000000110;
    x_8 = 'b111011111;
    x_9 = 'b111011110;
    x_10 = 'b111011010;
    x_11 = 'b111001100;
    x_12 = 'b111001011;
    x_13 = 'b111001001;
    x_14 = 'b111110110;
    x_15 = 'b111101011;
    x_16 = 'b111100101;
    x_17 = 'b111100011;
    x_18 = 'b111100101;
    x_19 = 'b111100010;
    x_20 = 'b111010111;
    x_21 = 'b111110000;
    x_22 = 'b111100010;
    x_23 = 'b111100001;
    x_24 = 'b000000011;
    x_25 = 'b000000010;
    x_26 = 'b111001010;
    x_27 = 'b111001000;
    x_28 = 'b111011011;
    x_29 = 'b111111111;
    x_30 = 'b111110101;
    x_31 = 'b111001011;
    x_32 = 'b111010011;
    x_33 = 'b111001000;
    x_34 = 'b111000101;
    x_35 = 'b111010001;
    x_36 = 'b111001110;
    x_37 = 'b111111110;
    x_38 = 'b000000010;
    x_39 = 'b111010110;
    x_40 = 'b111111000;
    x_41 = 'b111100000;
    x_42 = 'b111110111;
    x_43 = 'b000000000;
    x_44 = 'b111111110;
    x_45 = 'b111111000;
    x_46 = 'b111101101;
    x_47 = 'b111101110;
    x_48 = 'b111101101;
    x_49 = 'b111110000;
    x_50 = 'b111110011;
    x_51 = 'b111111000;
    x_52 = 'b111110111;
    x_53 = 'b111111000;
    x_54 = 'b111101111;
    x_55 = 'b111110100;
    x_56 = 'b111101011;
    x_57 = 'b000000001;
    x_58 = 'b111111001;
    x_59 = 'b111101010;
    x_60 = 'b111110101;
    x_61 = 'b111110001;
    x_62 = 'b111111011;
    x_63 = 'b111101110;
    x_64 = 'b111101101;
    x_65 = 'b111100001;
    x_66 = 'b111010000;
    x_67 = 'b111000000;
    x_68 = 'b111000000;
    x_69 = 'b110111110;
    x_70 = 'b111010110;
    x_71 = 'b000000110;
    x_72 = 'b111011111;
    x_73 = 'b111011110;
    x_74 = 'b111011010;
    x_75 = 'b111001100;
    x_76 = 'b111001011;
    x_77 = 'b111001001;
    x_78 = 'b111110110;
    x_79 = 'b111101011;
    x_80 = 'b111100101;
    x_81 = 'b111100011;
    x_82 = 'b111100101;
    x_83 = 'b111100010;
    x_84 = 'b111010111;
    x_85 = 'b111110000;
    x_86 = 'b111100010;
    x_87 = 'b111100001;
    x_88 = 'b000000011;
    x_89 = 'b000000010;
    x_90 = 'b111001010;
    x_91 = 'b111001000;
    x_92 = 'b111011011;
    x_93 = 'b111111111;
    x_94 = 'b111110101;
    x_95 = 'b111001011;
    x_96 = 'b111010011;
    x_97 = 'b111001000;
    x_98 = 'b111000101;
    x_99 = 'b111010001;
    x_100 = 'b111001110;
    x_101 = 'b111111110;
    x_102 = 'b000000010;
    x_103 = 'b111010110;
    x_104 = 'b111111000;
    x_105 = 'b111100000;
    x_106 = 'b111110111;
    x_107 = 'b000000000;
    x_108 = 'b111111110;
    x_109 = 'b111111000;
    x_110 = 'b111101101;
    x_111 = 'b111101110;
    x_112 = 'b111101101;
    x_113 = 'b111110000;
    x_114 = 'b111110011;
    x_115 = 'b111111000;
    x_116 = 'b111110111;
    x_117 = 'b111111000;
    x_118 = 'b111101111;
    x_119 = 'b111110100;
    x_120 = 'b111101011;
    x_121 = 'b000000001;
    x_122 = 'b111111001;
    x_123 = 'b111101010;
    x_124 = 'b111110101;
    x_125 = 'b111110001;
    x_126 = 'b111111011;
    x_127 = 'b111101110;
    x_128 = 'b111101101;
    x_129 = 'b111100001;
    x_130 = 'b111010000;
    x_131 = 'b111000000;
    x_132 = 'b111000000;
    x_133 = 'b110111110;
    x_134 = 'b111010110;
    x_135 = 'b000000110;
    x_136 = 'b111011111;
    x_137 = 'b111011110;
    x_138 = 'b111011010;
    x_139 = 'b111001100;
    x_140 = 'b111001011;
    x_141 = 'b111001001;
    x_142 = 'b111110110;
    x_143 = 'b111101011;
    x_144 = 'b111100101;
    x_145 = 'b111100011;
    x_146 = 'b111100101;
    x_147 = 'b111100010;
    x_148 = 'b111010111;
    x_149 = 'b111110000;
    x_150 = 'b111100010;
    x_151 = 'b111100001;
    x_152 = 'b000000011;
    x_153 = 'b000000010;
    x_154 = 'b111001010;
    x_155 = 'b111001000;
    x_156 = 'b111011011;
    x_157 = 'b111111111;
    x_158 = 'b111110101;
    x_159 = 'b111001011;
    x_160 = 'b111010011;
    x_161 = 'b111001000;
    x_162 = 'b111000101;
    x_163 = 'b111010001;
    x_164 = 'b111001110;
    x_165 = 'b111111110;
    x_166 = 'b000000010;
    x_167 = 'b111010110;
    x_168 = 'b111111000;
    x_169 = 'b111100000;
    x_170 = 'b111110111;
    x_171 = 'b000000000;
    x_172 = 'b111111110;
    x_173 = 'b111111000;
    x_174 = 'b111101101;
    x_175 = 'b111101110;
    x_176 = 'b111101101;
    x_177 = 'b111110000;
    x_178 = 'b111110011;
    x_179 = 'b111111000;
    x_180 = 'b111110111;
    x_181 = 'b111111000;
    x_182 = 'b111101111;
    x_183 = 'b111110100;
    x_184 = 'b111101011;
    x_185 = 'b000000001;
    x_186 = 'b111111001;
    x_187 = 'b111101010;
    x_188 = 'b111110101;
    x_189 = 'b111110001;
    x_190 = 'b111111011;
    x_191 = 'b111101110;
    x_192 = 'b111101101;
    x_193 = 'b111100001;
    x_194 = 'b111010000;
    x_195 = 'b111000000;
    x_196 = 'b111000000;
    x_197 = 'b110111110;
    x_198 = 'b111010110;
    x_199 = 'b000000110;
    x_200 = 'b111011111;
    x_201 = 'b111011110;
    x_202 = 'b111011010;
    x_203 = 'b111001100;
    x_204 = 'b111001011;
    x_205 = 'b111001001;
    x_206 = 'b111110110;
    x_207 = 'b111101011;
    x_208 = 'b111100101;
    x_209 = 'b111100011;
    x_210 = 'b111100101;
    x_211 = 'b111100010;
    x_212 = 'b111010111;
    x_213 = 'b111110000;
    x_214 = 'b111100010;
    x_215 = 'b111100001;
    x_216 = 'b000000011;
    x_217 = 'b000000010;
    x_218 = 'b111001010;
    x_219 = 'b111001000;
    x_220 = 'b111011011;
    x_221 = 'b111111111;
    x_222 = 'b111110101;
    x_223 = 'b111001011;
    x_224 = 'b111010011;
    x_225 = 'b111001000;
    x_226 = 'b111000101;
    x_227 = 'b111010001;
    x_228 = 'b111001110;
    x_229 = 'b111111110;
    x_230 = 'b000000010;
    x_231 = 'b111010110;
    x_232 = 'b111111000;
    x_233 = 'b111100000;
    x_234 = 'b111110111;
    x_235 = 'b000000000;
    x_236 = 'b111111110;
    x_237 = 'b111111000;
    x_238 = 'b111101101;
    x_239 = 'b111101110;
    x_240 = 'b111101101;
    x_241 = 'b111110000;
    x_242 = 'b111110011;
    x_243 = 'b111111000;
    x_244 = 'b111110111;
    x_245 = 'b111111000;
    x_246 = 'b111101111;
    x_247 = 'b111110100;
    x_248 = 'b111101011;
    x_249 = 'b000000001;
    x_250 = 'b111111001;
    x_251 = 'b111101010;
    x_252 = 'b111110101;
    x_253 = 'b111110001;
    x_254 = 'b111111011;
    x_255 = 'b111101110;

    h_0 = 'b111101101;
    h_1 = 'b111100001;
    h_2 = 'b111010000;
    h_3 = 'b111000000;
    h_4 = 'b111000000;
    h_5 = 'b110111110;
    h_6 = 'b111010110;
    h_7 = 'b000000110;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111111101;
    x_1 = 'b111110000;
    x_2 = 'b111100001;
    x_3 = 'b111010110;
    x_4 = 'b111010110;
    x_5 = 'b111010010;
    x_6 = 'b111101001;
    x_7 = 'b000001101;
    x_8 = 'b111100110;
    x_9 = 'b111101100;
    x_10 = 'b111101100;
    x_11 = 'b111011011;
    x_12 = 'b111011101;
    x_13 = 'b111011001;
    x_14 = 'b111101110;
    x_15 = 'b111101101;
    x_16 = 'b111101101;
    x_17 = 'b111101100;
    x_18 = 'b111101101;
    x_19 = 'b111101001;
    x_20 = 'b111011111;
    x_21 = 'b111110100;
    x_22 = 'b111101000;
    x_23 = 'b111101001;
    x_24 = 'b000000110;
    x_25 = 'b000000101;
    x_26 = 'b111010100;
    x_27 = 'b111010011;
    x_28 = 'b111100101;
    x_29 = 'b000000010;
    x_30 = 'b111111110;
    x_31 = 'b111011001;
    x_32 = 'b111011100;
    x_33 = 'b111010100;
    x_34 = 'b111010001;
    x_35 = 'b111011100;
    x_36 = 'b111011100;
    x_37 = 'b000000111;
    x_38 = 'b000000001;
    x_39 = 'b111100001;
    x_40 = 'b111110011;
    x_41 = 'b111011101;
    x_42 = 'b000001111;
    x_43 = 'b111111011;
    x_44 = 'b000000101;
    x_45 = 'b111101111;
    x_46 = 'b111101101;
    x_47 = 'b111101010;
    x_48 = 'b111101001;
    x_49 = 'b111101110;
    x_50 = 'b111110011;
    x_51 = 'b111110110;
    x_52 = 'b111110011;
    x_53 = 'b111110011;
    x_54 = 'b111100000;
    x_55 = 'b111101100;
    x_56 = 'b111100011;
    x_57 = 'b111111010;
    x_58 = 'b111101101;
    x_59 = 'b111011110;
    x_60 = 'b111101101;
    x_61 = 'b111101001;
    x_62 = 'b111110001;
    x_63 = 'b111100111;
    x_64 = 'b111111101;
    x_65 = 'b111110000;
    x_66 = 'b111100001;
    x_67 = 'b111010110;
    x_68 = 'b111010110;
    x_69 = 'b111010010;
    x_70 = 'b111101001;
    x_71 = 'b000001101;
    x_72 = 'b111100110;
    x_73 = 'b111101100;
    x_74 = 'b111101100;
    x_75 = 'b111011011;
    x_76 = 'b111011101;
    x_77 = 'b111011001;
    x_78 = 'b111101110;
    x_79 = 'b111101101;
    x_80 = 'b111101101;
    x_81 = 'b111101100;
    x_82 = 'b111101101;
    x_83 = 'b111101001;
    x_84 = 'b111011111;
    x_85 = 'b111110100;
    x_86 = 'b111101000;
    x_87 = 'b111101001;
    x_88 = 'b000000110;
    x_89 = 'b000000101;
    x_90 = 'b111010100;
    x_91 = 'b111010011;
    x_92 = 'b111100101;
    x_93 = 'b000000010;
    x_94 = 'b111111110;
    x_95 = 'b111011001;
    x_96 = 'b111011100;
    x_97 = 'b111010100;
    x_98 = 'b111010001;
    x_99 = 'b111011100;
    x_100 = 'b111011100;
    x_101 = 'b000000111;
    x_102 = 'b000000001;
    x_103 = 'b111100001;
    x_104 = 'b111110011;
    x_105 = 'b111011101;
    x_106 = 'b000001111;
    x_107 = 'b111111011;
    x_108 = 'b000000101;
    x_109 = 'b111101111;
    x_110 = 'b111101101;
    x_111 = 'b111101010;
    x_112 = 'b111101001;
    x_113 = 'b111101110;
    x_114 = 'b111110011;
    x_115 = 'b111110110;
    x_116 = 'b111110011;
    x_117 = 'b111110011;
    x_118 = 'b111100000;
    x_119 = 'b111101100;
    x_120 = 'b111100011;
    x_121 = 'b111111010;
    x_122 = 'b111101101;
    x_123 = 'b111011110;
    x_124 = 'b111101101;
    x_125 = 'b111101001;
    x_126 = 'b111110001;
    x_127 = 'b111100111;
    x_128 = 'b111111101;
    x_129 = 'b111110000;
    x_130 = 'b111100001;
    x_131 = 'b111010110;
    x_132 = 'b111010110;
    x_133 = 'b111010010;
    x_134 = 'b111101001;
    x_135 = 'b000001101;
    x_136 = 'b111100110;
    x_137 = 'b111101100;
    x_138 = 'b111101100;
    x_139 = 'b111011011;
    x_140 = 'b111011101;
    x_141 = 'b111011001;
    x_142 = 'b111101110;
    x_143 = 'b111101101;
    x_144 = 'b111101101;
    x_145 = 'b111101100;
    x_146 = 'b111101101;
    x_147 = 'b111101001;
    x_148 = 'b111011111;
    x_149 = 'b111110100;
    x_150 = 'b111101000;
    x_151 = 'b111101001;
    x_152 = 'b000000110;
    x_153 = 'b000000101;
    x_154 = 'b111010100;
    x_155 = 'b111010011;
    x_156 = 'b111100101;
    x_157 = 'b000000010;
    x_158 = 'b111111110;
    x_159 = 'b111011001;
    x_160 = 'b111011100;
    x_161 = 'b111010100;
    x_162 = 'b111010001;
    x_163 = 'b111011100;
    x_164 = 'b111011100;
    x_165 = 'b000000111;
    x_166 = 'b000000001;
    x_167 = 'b111100001;
    x_168 = 'b111110011;
    x_169 = 'b111011101;
    x_170 = 'b000001111;
    x_171 = 'b111111011;
    x_172 = 'b000000101;
    x_173 = 'b111101111;
    x_174 = 'b111101101;
    x_175 = 'b111101010;
    x_176 = 'b111101001;
    x_177 = 'b111101110;
    x_178 = 'b111110011;
    x_179 = 'b111110110;
    x_180 = 'b111110011;
    x_181 = 'b111110011;
    x_182 = 'b111100000;
    x_183 = 'b111101100;
    x_184 = 'b111100011;
    x_185 = 'b111111010;
    x_186 = 'b111101101;
    x_187 = 'b111011110;
    x_188 = 'b111101101;
    x_189 = 'b111101001;
    x_190 = 'b111110001;
    x_191 = 'b111100111;
    x_192 = 'b111111101;
    x_193 = 'b111110000;
    x_194 = 'b111100001;
    x_195 = 'b111010110;
    x_196 = 'b111010110;
    x_197 = 'b111010010;
    x_198 = 'b111101001;
    x_199 = 'b000001101;
    x_200 = 'b111100110;
    x_201 = 'b111101100;
    x_202 = 'b111101100;
    x_203 = 'b111011011;
    x_204 = 'b111011101;
    x_205 = 'b111011001;
    x_206 = 'b111101110;
    x_207 = 'b111101101;
    x_208 = 'b111101101;
    x_209 = 'b111101100;
    x_210 = 'b111101101;
    x_211 = 'b111101001;
    x_212 = 'b111011111;
    x_213 = 'b111110100;
    x_214 = 'b111101000;
    x_215 = 'b111101001;
    x_216 = 'b000000110;
    x_217 = 'b000000101;
    x_218 = 'b111010100;
    x_219 = 'b111010011;
    x_220 = 'b111100101;
    x_221 = 'b000000010;
    x_222 = 'b111111110;
    x_223 = 'b111011001;
    x_224 = 'b111011100;
    x_225 = 'b111010100;
    x_226 = 'b111010001;
    x_227 = 'b111011100;
    x_228 = 'b111011100;
    x_229 = 'b000000111;
    x_230 = 'b000000001;
    x_231 = 'b111100001;
    x_232 = 'b111110011;
    x_233 = 'b111011101;
    x_234 = 'b000001111;
    x_235 = 'b111111011;
    x_236 = 'b000000101;
    x_237 = 'b111101111;
    x_238 = 'b111101101;
    x_239 = 'b111101010;
    x_240 = 'b111101001;
    x_241 = 'b111101110;
    x_242 = 'b111110011;
    x_243 = 'b111110110;
    x_244 = 'b111110011;
    x_245 = 'b111110011;
    x_246 = 'b111100000;
    x_247 = 'b111101100;
    x_248 = 'b111100011;
    x_249 = 'b111111010;
    x_250 = 'b111101101;
    x_251 = 'b111011110;
    x_252 = 'b111101101;
    x_253 = 'b111101001;
    x_254 = 'b111110001;
    x_255 = 'b111100111;

    h_0 = 'b111111101;
    h_1 = 'b111110000;
    h_2 = 'b111100001;
    h_3 = 'b111010110;
    h_4 = 'b111010110;
    h_5 = 'b111010010;
    h_6 = 'b111101001;
    h_7 = 'b000001101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111111011;
    x_1 = 'b111101111;
    x_2 = 'b111100010;
    x_3 = 'b111011010;
    x_4 = 'b111011001;
    x_5 = 'b111010100;
    x_6 = 'b111100110;
    x_7 = 'b000001000;
    x_8 = 'b111100100;
    x_9 = 'b111101000;
    x_10 = 'b111100110;
    x_11 = 'b111010110;
    x_12 = 'b111011011;
    x_13 = 'b111011100;
    x_14 = 'b111101101;
    x_15 = 'b111101001;
    x_16 = 'b111101001;
    x_17 = 'b111100101;
    x_18 = 'b111100101;
    x_19 = 'b111100001;
    x_20 = 'b111011000;
    x_21 = 'b111110101;
    x_22 = 'b111101001;
    x_23 = 'b111101100;
    x_24 = 'b000000110;
    x_25 = 'b000000101;
    x_26 = 'b111010100;
    x_27 = 'b111010111;
    x_28 = 'b111101000;
    x_29 = 'b000000011;
    x_30 = 'b111111111;
    x_31 = 'b111011010;
    x_32 = 'b111011011;
    x_33 = 'b111010010;
    x_34 = 'b111010001;
    x_35 = 'b111011101;
    x_36 = 'b111011100;
    x_37 = 'b000001101;
    x_38 = 'b111111111;
    x_39 = 'b111100010;
    x_40 = 'b000001011;
    x_41 = 'b111011000;
    x_42 = 'b000001001;
    x_43 = 'b111001011;
    x_44 = 'b000010100;
    x_45 = 'b111011001;
    x_46 = 'b111110001;
    x_47 = 'b111101011;
    x_48 = 'b111100111;
    x_49 = 'b111101000;
    x_50 = 'b111100111;
    x_51 = 'b111100101;
    x_52 = 'b111100001;
    x_53 = 'b111100000;
    x_54 = 'b111010001;
    x_55 = 'b111100110;
    x_56 = 'b111011101;
    x_57 = 'b111101110;
    x_58 = 'b111011000;
    x_59 = 'b111001111;
    x_60 = 'b111100010;
    x_61 = 'b111011010;
    x_62 = 'b111011011;
    x_63 = 'b111011110;
    x_64 = 'b111111011;
    x_65 = 'b111101111;
    x_66 = 'b111100010;
    x_67 = 'b111011010;
    x_68 = 'b111011001;
    x_69 = 'b111010100;
    x_70 = 'b111100110;
    x_71 = 'b000001000;
    x_72 = 'b111100100;
    x_73 = 'b111101000;
    x_74 = 'b111100110;
    x_75 = 'b111010110;
    x_76 = 'b111011011;
    x_77 = 'b111011100;
    x_78 = 'b111101101;
    x_79 = 'b111101001;
    x_80 = 'b111101001;
    x_81 = 'b111100101;
    x_82 = 'b111100101;
    x_83 = 'b111100001;
    x_84 = 'b111011000;
    x_85 = 'b111110101;
    x_86 = 'b111101001;
    x_87 = 'b111101100;
    x_88 = 'b000000110;
    x_89 = 'b000000101;
    x_90 = 'b111010100;
    x_91 = 'b111010111;
    x_92 = 'b111101000;
    x_93 = 'b000000011;
    x_94 = 'b111111111;
    x_95 = 'b111011010;
    x_96 = 'b111011011;
    x_97 = 'b111010010;
    x_98 = 'b111010001;
    x_99 = 'b111011101;
    x_100 = 'b111011100;
    x_101 = 'b000001101;
    x_102 = 'b111111111;
    x_103 = 'b111100010;
    x_104 = 'b000001011;
    x_105 = 'b111011000;
    x_106 = 'b000001001;
    x_107 = 'b111001011;
    x_108 = 'b000010100;
    x_109 = 'b111011001;
    x_110 = 'b111110001;
    x_111 = 'b111101011;
    x_112 = 'b111100111;
    x_113 = 'b111101000;
    x_114 = 'b111100111;
    x_115 = 'b111100101;
    x_116 = 'b111100001;
    x_117 = 'b111100000;
    x_118 = 'b111010001;
    x_119 = 'b111100110;
    x_120 = 'b111011101;
    x_121 = 'b111101110;
    x_122 = 'b111011000;
    x_123 = 'b111001111;
    x_124 = 'b111100010;
    x_125 = 'b111011010;
    x_126 = 'b111011011;
    x_127 = 'b111011110;
    x_128 = 'b111111011;
    x_129 = 'b111101111;
    x_130 = 'b111100010;
    x_131 = 'b111011010;
    x_132 = 'b111011001;
    x_133 = 'b111010100;
    x_134 = 'b111100110;
    x_135 = 'b000001000;
    x_136 = 'b111100100;
    x_137 = 'b111101000;
    x_138 = 'b111100110;
    x_139 = 'b111010110;
    x_140 = 'b111011011;
    x_141 = 'b111011100;
    x_142 = 'b111101101;
    x_143 = 'b111101001;
    x_144 = 'b111101001;
    x_145 = 'b111100101;
    x_146 = 'b111100101;
    x_147 = 'b111100001;
    x_148 = 'b111011000;
    x_149 = 'b111110101;
    x_150 = 'b111101001;
    x_151 = 'b111101100;
    x_152 = 'b000000110;
    x_153 = 'b000000101;
    x_154 = 'b111010100;
    x_155 = 'b111010111;
    x_156 = 'b111101000;
    x_157 = 'b000000011;
    x_158 = 'b111111111;
    x_159 = 'b111011010;
    x_160 = 'b111011011;
    x_161 = 'b111010010;
    x_162 = 'b111010001;
    x_163 = 'b111011101;
    x_164 = 'b111011100;
    x_165 = 'b000001101;
    x_166 = 'b111111111;
    x_167 = 'b111100010;
    x_168 = 'b000001011;
    x_169 = 'b111011000;
    x_170 = 'b000001001;
    x_171 = 'b111001011;
    x_172 = 'b000010100;
    x_173 = 'b111011001;
    x_174 = 'b111110001;
    x_175 = 'b111101011;
    x_176 = 'b111100111;
    x_177 = 'b111101000;
    x_178 = 'b111100111;
    x_179 = 'b111100101;
    x_180 = 'b111100001;
    x_181 = 'b111100000;
    x_182 = 'b111010001;
    x_183 = 'b111100110;
    x_184 = 'b111011101;
    x_185 = 'b111101110;
    x_186 = 'b111011000;
    x_187 = 'b111001111;
    x_188 = 'b111100010;
    x_189 = 'b111011010;
    x_190 = 'b111011011;
    x_191 = 'b111011110;
    x_192 = 'b111111011;
    x_193 = 'b111101111;
    x_194 = 'b111100010;
    x_195 = 'b111011010;
    x_196 = 'b111011001;
    x_197 = 'b111010100;
    x_198 = 'b111100110;
    x_199 = 'b000001000;
    x_200 = 'b111100100;
    x_201 = 'b111101000;
    x_202 = 'b111100110;
    x_203 = 'b111010110;
    x_204 = 'b111011011;
    x_205 = 'b111011100;
    x_206 = 'b111101101;
    x_207 = 'b111101001;
    x_208 = 'b111101001;
    x_209 = 'b111100101;
    x_210 = 'b111100101;
    x_211 = 'b111100001;
    x_212 = 'b111011000;
    x_213 = 'b111110101;
    x_214 = 'b111101001;
    x_215 = 'b111101100;
    x_216 = 'b000000110;
    x_217 = 'b000000101;
    x_218 = 'b111010100;
    x_219 = 'b111010111;
    x_220 = 'b111101000;
    x_221 = 'b000000011;
    x_222 = 'b111111111;
    x_223 = 'b111011010;
    x_224 = 'b111011011;
    x_225 = 'b111010010;
    x_226 = 'b111010001;
    x_227 = 'b111011101;
    x_228 = 'b111011100;
    x_229 = 'b000001101;
    x_230 = 'b111111111;
    x_231 = 'b111100010;
    x_232 = 'b000001011;
    x_233 = 'b111011000;
    x_234 = 'b000001001;
    x_235 = 'b111001011;
    x_236 = 'b000010100;
    x_237 = 'b111011001;
    x_238 = 'b111110001;
    x_239 = 'b111101011;
    x_240 = 'b111100111;
    x_241 = 'b111101000;
    x_242 = 'b111100111;
    x_243 = 'b111100101;
    x_244 = 'b111100001;
    x_245 = 'b111100000;
    x_246 = 'b111010001;
    x_247 = 'b111100110;
    x_248 = 'b111011101;
    x_249 = 'b111101110;
    x_250 = 'b111011000;
    x_251 = 'b111001111;
    x_252 = 'b111100010;
    x_253 = 'b111011010;
    x_254 = 'b111011011;
    x_255 = 'b111011110;

    h_0 = 'b111111011;
    h_1 = 'b111101111;
    h_2 = 'b111100010;
    h_3 = 'b111011010;
    h_4 = 'b111011001;
    h_5 = 'b111010100;
    h_6 = 'b111100110;
    h_7 = 'b000001000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111111010;
    x_1 = 'b111101100;
    x_2 = 'b111011100;
    x_3 = 'b111010001;
    x_4 = 'b111010001;
    x_5 = 'b111001101;
    x_6 = 'b111011101;
    x_7 = 'b000000111;
    x_8 = 'b111100110;
    x_9 = 'b111100010;
    x_10 = 'b111011100;
    x_11 = 'b111001010;
    x_12 = 'b111010100;
    x_13 = 'b111010000;
    x_14 = 'b111111000;
    x_15 = 'b111101000;
    x_16 = 'b111100010;
    x_17 = 'b111011010;
    x_18 = 'b111011011;
    x_19 = 'b111010111;
    x_20 = 'b111001111;
    x_21 = 'b111110100;
    x_22 = 'b111100111;
    x_23 = 'b111100111;
    x_24 = 'b000000110;
    x_25 = 'b000000101;
    x_26 = 'b111010000;
    x_27 = 'b111010001;
    x_28 = 'b111100011;
    x_29 = 'b000000100;
    x_30 = 'b111111010;
    x_31 = 'b111010010;
    x_32 = 'b111010111;
    x_33 = 'b111001100;
    x_34 = 'b111001010;
    x_35 = 'b111010111;
    x_36 = 'b111010001;
    x_37 = 'b000000001;
    x_38 = 'b000001001;
    x_39 = 'b111001110;
    x_40 = 'b000010110;
    x_41 = 'b110100110;
    x_42 = 'b000010001;
    x_43 = 'b111110111;
    x_44 = 'b000010011;
    x_45 = 'b111100100;
    x_46 = 'b111101111;
    x_47 = 'b111101001;
    x_48 = 'b111100011;
    x_49 = 'b111100000;
    x_50 = 'b111011101;
    x_51 = 'b111011000;
    x_52 = 'b111011000;
    x_53 = 'b111011100;
    x_54 = 'b111010111;
    x_55 = 'b111100010;
    x_56 = 'b111011010;
    x_57 = 'b111100011;
    x_58 = 'b111010000;
    x_59 = 'b111001111;
    x_60 = 'b111011001;
    x_61 = 'b111001111;
    x_62 = 'b111001001;
    x_63 = 'b111011010;
    x_64 = 'b111111010;
    x_65 = 'b111101100;
    x_66 = 'b111011100;
    x_67 = 'b111010001;
    x_68 = 'b111010001;
    x_69 = 'b111001101;
    x_70 = 'b111011101;
    x_71 = 'b000000111;
    x_72 = 'b111100110;
    x_73 = 'b111100010;
    x_74 = 'b111011100;
    x_75 = 'b111001010;
    x_76 = 'b111010100;
    x_77 = 'b111010000;
    x_78 = 'b111111000;
    x_79 = 'b111101000;
    x_80 = 'b111100010;
    x_81 = 'b111011010;
    x_82 = 'b111011011;
    x_83 = 'b111010111;
    x_84 = 'b111001111;
    x_85 = 'b111110100;
    x_86 = 'b111100111;
    x_87 = 'b111100111;
    x_88 = 'b000000110;
    x_89 = 'b000000101;
    x_90 = 'b111010000;
    x_91 = 'b111010001;
    x_92 = 'b111100011;
    x_93 = 'b000000100;
    x_94 = 'b111111010;
    x_95 = 'b111010010;
    x_96 = 'b111010111;
    x_97 = 'b111001100;
    x_98 = 'b111001010;
    x_99 = 'b111010111;
    x_100 = 'b111010001;
    x_101 = 'b000000001;
    x_102 = 'b000001001;
    x_103 = 'b111001110;
    x_104 = 'b000010110;
    x_105 = 'b110100110;
    x_106 = 'b000010001;
    x_107 = 'b111110111;
    x_108 = 'b000010011;
    x_109 = 'b111100100;
    x_110 = 'b111101111;
    x_111 = 'b111101001;
    x_112 = 'b111100011;
    x_113 = 'b111100000;
    x_114 = 'b111011101;
    x_115 = 'b111011000;
    x_116 = 'b111011000;
    x_117 = 'b111011100;
    x_118 = 'b111010111;
    x_119 = 'b111100010;
    x_120 = 'b111011010;
    x_121 = 'b111100011;
    x_122 = 'b111010000;
    x_123 = 'b111001111;
    x_124 = 'b111011001;
    x_125 = 'b111001111;
    x_126 = 'b111001001;
    x_127 = 'b111011010;
    x_128 = 'b111111010;
    x_129 = 'b111101100;
    x_130 = 'b111011100;
    x_131 = 'b111010001;
    x_132 = 'b111010001;
    x_133 = 'b111001101;
    x_134 = 'b111011101;
    x_135 = 'b000000111;
    x_136 = 'b111100110;
    x_137 = 'b111100010;
    x_138 = 'b111011100;
    x_139 = 'b111001010;
    x_140 = 'b111010100;
    x_141 = 'b111010000;
    x_142 = 'b111111000;
    x_143 = 'b111101000;
    x_144 = 'b111100010;
    x_145 = 'b111011010;
    x_146 = 'b111011011;
    x_147 = 'b111010111;
    x_148 = 'b111001111;
    x_149 = 'b111110100;
    x_150 = 'b111100111;
    x_151 = 'b111100111;
    x_152 = 'b000000110;
    x_153 = 'b000000101;
    x_154 = 'b111010000;
    x_155 = 'b111010001;
    x_156 = 'b111100011;
    x_157 = 'b000000100;
    x_158 = 'b111111010;
    x_159 = 'b111010010;
    x_160 = 'b111010111;
    x_161 = 'b111001100;
    x_162 = 'b111001010;
    x_163 = 'b111010111;
    x_164 = 'b111010001;
    x_165 = 'b000000001;
    x_166 = 'b000001001;
    x_167 = 'b111001110;
    x_168 = 'b000010110;
    x_169 = 'b110100110;
    x_170 = 'b000010001;
    x_171 = 'b111110111;
    x_172 = 'b000010011;
    x_173 = 'b111100100;
    x_174 = 'b111101111;
    x_175 = 'b111101001;
    x_176 = 'b111100011;
    x_177 = 'b111100000;
    x_178 = 'b111011101;
    x_179 = 'b111011000;
    x_180 = 'b111011000;
    x_181 = 'b111011100;
    x_182 = 'b111010111;
    x_183 = 'b111100010;
    x_184 = 'b111011010;
    x_185 = 'b111100011;
    x_186 = 'b111010000;
    x_187 = 'b111001111;
    x_188 = 'b111011001;
    x_189 = 'b111001111;
    x_190 = 'b111001001;
    x_191 = 'b111011010;
    x_192 = 'b111111010;
    x_193 = 'b111101100;
    x_194 = 'b111011100;
    x_195 = 'b111010001;
    x_196 = 'b111010001;
    x_197 = 'b111001101;
    x_198 = 'b111011101;
    x_199 = 'b000000111;
    x_200 = 'b111100110;
    x_201 = 'b111100010;
    x_202 = 'b111011100;
    x_203 = 'b111001010;
    x_204 = 'b111010100;
    x_205 = 'b111010000;
    x_206 = 'b111111000;
    x_207 = 'b111101000;
    x_208 = 'b111100010;
    x_209 = 'b111011010;
    x_210 = 'b111011011;
    x_211 = 'b111010111;
    x_212 = 'b111001111;
    x_213 = 'b111110100;
    x_214 = 'b111100111;
    x_215 = 'b111100111;
    x_216 = 'b000000110;
    x_217 = 'b000000101;
    x_218 = 'b111010000;
    x_219 = 'b111010001;
    x_220 = 'b111100011;
    x_221 = 'b000000100;
    x_222 = 'b111111010;
    x_223 = 'b111010010;
    x_224 = 'b111010111;
    x_225 = 'b111001100;
    x_226 = 'b111001010;
    x_227 = 'b111010111;
    x_228 = 'b111010001;
    x_229 = 'b000000001;
    x_230 = 'b000001001;
    x_231 = 'b111001110;
    x_232 = 'b000010110;
    x_233 = 'b110100110;
    x_234 = 'b000010001;
    x_235 = 'b111110111;
    x_236 = 'b000010011;
    x_237 = 'b111100100;
    x_238 = 'b111101111;
    x_239 = 'b111101001;
    x_240 = 'b111100011;
    x_241 = 'b111100000;
    x_242 = 'b111011101;
    x_243 = 'b111011000;
    x_244 = 'b111011000;
    x_245 = 'b111011100;
    x_246 = 'b111010111;
    x_247 = 'b111100010;
    x_248 = 'b111011010;
    x_249 = 'b111100011;
    x_250 = 'b111010000;
    x_251 = 'b111001111;
    x_252 = 'b111011001;
    x_253 = 'b111001111;
    x_254 = 'b111001001;
    x_255 = 'b111011010;

    h_0 = 'b111111010;
    h_1 = 'b111101100;
    h_2 = 'b111011100;
    h_3 = 'b111010001;
    h_4 = 'b111010001;
    h_5 = 'b111001101;
    h_6 = 'b111011101;
    h_7 = 'b000000111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111110111;
    x_1 = 'b111100111;
    x_2 = 'b111010110;
    x_3 = 'b111001110;
    x_4 = 'b111001101;
    x_5 = 'b111001010;
    x_6 = 'b111010011;
    x_7 = 'b000000001;
    x_8 = 'b111100000;
    x_9 = 'b111011011;
    x_10 = 'b111011000;
    x_11 = 'b111001001;
    x_12 = 'b111010000;
    x_13 = 'b111000000;
    x_14 = 'b111110010;
    x_15 = 'b111100011;
    x_16 = 'b111011100;
    x_17 = 'b111010100;
    x_18 = 'b111011000;
    x_19 = 'b111010100;
    x_20 = 'b111001101;
    x_21 = 'b111110000;
    x_22 = 'b111100011;
    x_23 = 'b111100010;
    x_24 = 'b000000100;
    x_25 = 'b000000100;
    x_26 = 'b111001110;
    x_27 = 'b111001101;
    x_28 = 'b111100001;
    x_29 = 'b000000100;
    x_30 = 'b111111011;
    x_31 = 'b111010001;
    x_32 = 'b111010001;
    x_33 = 'b111001001;
    x_34 = 'b111000111;
    x_35 = 'b111010011;
    x_36 = 'b111001110;
    x_37 = 'b111111010;
    x_38 = 'b000000001;
    x_39 = 'b111001011;
    x_40 = 'b000001001;
    x_41 = 'b111000100;
    x_42 = 'b000001100;
    x_43 = 'b111110101;
    x_44 = 'b000000101;
    x_45 = 'b111110010;
    x_46 = 'b111110101;
    x_47 = 'b111101010;
    x_48 = 'b111100010;
    x_49 = 'b111011110;
    x_50 = 'b111011100;
    x_51 = 'b111011011;
    x_52 = 'b111011111;
    x_53 = 'b111100111;
    x_54 = 'b111101001;
    x_55 = 'b111100011;
    x_56 = 'b111011100;
    x_57 = 'b111100110;
    x_58 = 'b111100001;
    x_59 = 'b111100110;
    x_60 = 'b111010111;
    x_61 = 'b111010001;
    x_62 = 'b111001011;
    x_63 = 'b111100011;
    x_64 = 'b111110111;
    x_65 = 'b111100111;
    x_66 = 'b111010110;
    x_67 = 'b111001110;
    x_68 = 'b111001101;
    x_69 = 'b111001010;
    x_70 = 'b111010011;
    x_71 = 'b000000001;
    x_72 = 'b111100000;
    x_73 = 'b111011011;
    x_74 = 'b111011000;
    x_75 = 'b111001001;
    x_76 = 'b111010000;
    x_77 = 'b111000000;
    x_78 = 'b111110010;
    x_79 = 'b111100011;
    x_80 = 'b111011100;
    x_81 = 'b111010100;
    x_82 = 'b111011000;
    x_83 = 'b111010100;
    x_84 = 'b111001101;
    x_85 = 'b111110000;
    x_86 = 'b111100011;
    x_87 = 'b111100010;
    x_88 = 'b000000100;
    x_89 = 'b000000100;
    x_90 = 'b111001110;
    x_91 = 'b111001101;
    x_92 = 'b111100001;
    x_93 = 'b000000100;
    x_94 = 'b111111011;
    x_95 = 'b111010001;
    x_96 = 'b111010001;
    x_97 = 'b111001001;
    x_98 = 'b111000111;
    x_99 = 'b111010011;
    x_100 = 'b111001110;
    x_101 = 'b111111010;
    x_102 = 'b000000001;
    x_103 = 'b111001011;
    x_104 = 'b000001001;
    x_105 = 'b111000100;
    x_106 = 'b000001100;
    x_107 = 'b111110101;
    x_108 = 'b000000101;
    x_109 = 'b111110010;
    x_110 = 'b111110101;
    x_111 = 'b111101010;
    x_112 = 'b111100010;
    x_113 = 'b111011110;
    x_114 = 'b111011100;
    x_115 = 'b111011011;
    x_116 = 'b111011111;
    x_117 = 'b111100111;
    x_118 = 'b111101001;
    x_119 = 'b111100011;
    x_120 = 'b111011100;
    x_121 = 'b111100110;
    x_122 = 'b111100001;
    x_123 = 'b111100110;
    x_124 = 'b111010111;
    x_125 = 'b111010001;
    x_126 = 'b111001011;
    x_127 = 'b111100011;
    x_128 = 'b111110111;
    x_129 = 'b111100111;
    x_130 = 'b111010110;
    x_131 = 'b111001110;
    x_132 = 'b111001101;
    x_133 = 'b111001010;
    x_134 = 'b111010011;
    x_135 = 'b000000001;
    x_136 = 'b111100000;
    x_137 = 'b111011011;
    x_138 = 'b111011000;
    x_139 = 'b111001001;
    x_140 = 'b111010000;
    x_141 = 'b111000000;
    x_142 = 'b111110010;
    x_143 = 'b111100011;
    x_144 = 'b111011100;
    x_145 = 'b111010100;
    x_146 = 'b111011000;
    x_147 = 'b111010100;
    x_148 = 'b111001101;
    x_149 = 'b111110000;
    x_150 = 'b111100011;
    x_151 = 'b111100010;
    x_152 = 'b000000100;
    x_153 = 'b000000100;
    x_154 = 'b111001110;
    x_155 = 'b111001101;
    x_156 = 'b111100001;
    x_157 = 'b000000100;
    x_158 = 'b111111011;
    x_159 = 'b111010001;
    x_160 = 'b111010001;
    x_161 = 'b111001001;
    x_162 = 'b111000111;
    x_163 = 'b111010011;
    x_164 = 'b111001110;
    x_165 = 'b111111010;
    x_166 = 'b000000001;
    x_167 = 'b111001011;
    x_168 = 'b000001001;
    x_169 = 'b111000100;
    x_170 = 'b000001100;
    x_171 = 'b111110101;
    x_172 = 'b000000101;
    x_173 = 'b111110010;
    x_174 = 'b111110101;
    x_175 = 'b111101010;
    x_176 = 'b111100010;
    x_177 = 'b111011110;
    x_178 = 'b111011100;
    x_179 = 'b111011011;
    x_180 = 'b111011111;
    x_181 = 'b111100111;
    x_182 = 'b111101001;
    x_183 = 'b111100011;
    x_184 = 'b111011100;
    x_185 = 'b111100110;
    x_186 = 'b111100001;
    x_187 = 'b111100110;
    x_188 = 'b111010111;
    x_189 = 'b111010001;
    x_190 = 'b111001011;
    x_191 = 'b111100011;
    x_192 = 'b111110111;
    x_193 = 'b111100111;
    x_194 = 'b111010110;
    x_195 = 'b111001110;
    x_196 = 'b111001101;
    x_197 = 'b111001010;
    x_198 = 'b111010011;
    x_199 = 'b000000001;
    x_200 = 'b111100000;
    x_201 = 'b111011011;
    x_202 = 'b111011000;
    x_203 = 'b111001001;
    x_204 = 'b111010000;
    x_205 = 'b111000000;
    x_206 = 'b111110010;
    x_207 = 'b111100011;
    x_208 = 'b111011100;
    x_209 = 'b111010100;
    x_210 = 'b111011000;
    x_211 = 'b111010100;
    x_212 = 'b111001101;
    x_213 = 'b111110000;
    x_214 = 'b111100011;
    x_215 = 'b111100010;
    x_216 = 'b000000100;
    x_217 = 'b000000100;
    x_218 = 'b111001110;
    x_219 = 'b111001101;
    x_220 = 'b111100001;
    x_221 = 'b000000100;
    x_222 = 'b111111011;
    x_223 = 'b111010001;
    x_224 = 'b111010001;
    x_225 = 'b111001001;
    x_226 = 'b111000111;
    x_227 = 'b111010011;
    x_228 = 'b111001110;
    x_229 = 'b111111010;
    x_230 = 'b000000001;
    x_231 = 'b111001011;
    x_232 = 'b000001001;
    x_233 = 'b111000100;
    x_234 = 'b000001100;
    x_235 = 'b111110101;
    x_236 = 'b000000101;
    x_237 = 'b111110010;
    x_238 = 'b111110101;
    x_239 = 'b111101010;
    x_240 = 'b111100010;
    x_241 = 'b111011110;
    x_242 = 'b111011100;
    x_243 = 'b111011011;
    x_244 = 'b111011111;
    x_245 = 'b111100111;
    x_246 = 'b111101001;
    x_247 = 'b111100011;
    x_248 = 'b111011100;
    x_249 = 'b111100110;
    x_250 = 'b111100001;
    x_251 = 'b111100110;
    x_252 = 'b111010111;
    x_253 = 'b111010001;
    x_254 = 'b111001011;
    x_255 = 'b111100011;

    h_0 = 'b111110111;
    h_1 = 'b111100111;
    h_2 = 'b111010110;
    h_3 = 'b111001110;
    h_4 = 'b111001101;
    h_5 = 'b111001010;
    h_6 = 'b111010011;
    h_7 = 'b000000001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111110110;
    x_1 = 'b111011111;
    x_2 = 'b111010000;
    x_3 = 'b111000111;
    x_4 = 'b111001000;
    x_5 = 'b111001010;
    x_6 = 'b111011001;
    x_7 = 'b000000000;
    x_8 = 'b111011010;
    x_9 = 'b111011000;
    x_10 = 'b111010101;
    x_11 = 'b111001001;
    x_12 = 'b111010010;
    x_13 = 'b111001100;
    x_14 = 'b111110001;
    x_15 = 'b111100100;
    x_16 = 'b111011100;
    x_17 = 'b111010101;
    x_18 = 'b111011011;
    x_19 = 'b111011001;
    x_20 = 'b111010011;
    x_21 = 'b111101100;
    x_22 = 'b111100001;
    x_23 = 'b111100000;
    x_24 = 'b000000001;
    x_25 = 'b000000000;
    x_26 = 'b111001100;
    x_27 = 'b111001100;
    x_28 = 'b111011111;
    x_29 = 'b000000011;
    x_30 = 'b111110110;
    x_31 = 'b111001111;
    x_32 = 'b111001101;
    x_33 = 'b111001000;
    x_34 = 'b111000111;
    x_35 = 'b111010010;
    x_36 = 'b111010011;
    x_37 = 'b111111001;
    x_38 = 'b111111011;
    x_39 = 'b111011001;
    x_40 = 'b111111101;
    x_41 = 'b111011111;
    x_42 = 'b111110101;
    x_43 = 'b111011101;
    x_44 = 'b000000010;
    x_45 = 'b111101001;
    x_46 = 'b111110011;
    x_47 = 'b111110000;
    x_48 = 'b111100111;
    x_49 = 'b111101001;
    x_50 = 'b111100011;
    x_51 = 'b111101100;
    x_52 = 'b111110000;
    x_53 = 'b111111011;
    x_54 = 'b111111100;
    x_55 = 'b111110000;
    x_56 = 'b111101010;
    x_57 = 'b111110101;
    x_58 = 'b111111111;
    x_59 = 'b000001100;
    x_60 = 'b111100100;
    x_61 = 'b111100110;
    x_62 = 'b111101001;
    x_63 = 'b111111001;
    x_64 = 'b111110110;
    x_65 = 'b111011111;
    x_66 = 'b111010000;
    x_67 = 'b111000111;
    x_68 = 'b111001000;
    x_69 = 'b111001010;
    x_70 = 'b111011001;
    x_71 = 'b000000000;
    x_72 = 'b111011010;
    x_73 = 'b111011000;
    x_74 = 'b111010101;
    x_75 = 'b111001001;
    x_76 = 'b111010010;
    x_77 = 'b111001100;
    x_78 = 'b111110001;
    x_79 = 'b111100100;
    x_80 = 'b111011100;
    x_81 = 'b111010101;
    x_82 = 'b111011011;
    x_83 = 'b111011001;
    x_84 = 'b111010011;
    x_85 = 'b111101100;
    x_86 = 'b111100001;
    x_87 = 'b111100000;
    x_88 = 'b000000001;
    x_89 = 'b000000000;
    x_90 = 'b111001100;
    x_91 = 'b111001100;
    x_92 = 'b111011111;
    x_93 = 'b000000011;
    x_94 = 'b111110110;
    x_95 = 'b111001111;
    x_96 = 'b111001101;
    x_97 = 'b111001000;
    x_98 = 'b111000111;
    x_99 = 'b111010010;
    x_100 = 'b111010011;
    x_101 = 'b111111001;
    x_102 = 'b111111011;
    x_103 = 'b111011001;
    x_104 = 'b111111101;
    x_105 = 'b111011111;
    x_106 = 'b111110101;
    x_107 = 'b111011101;
    x_108 = 'b000000010;
    x_109 = 'b111101001;
    x_110 = 'b111110011;
    x_111 = 'b111110000;
    x_112 = 'b111100111;
    x_113 = 'b111101001;
    x_114 = 'b111100011;
    x_115 = 'b111101100;
    x_116 = 'b111110000;
    x_117 = 'b111111011;
    x_118 = 'b111111100;
    x_119 = 'b111110000;
    x_120 = 'b111101010;
    x_121 = 'b111110101;
    x_122 = 'b111111111;
    x_123 = 'b000001100;
    x_124 = 'b111100100;
    x_125 = 'b111100110;
    x_126 = 'b111101001;
    x_127 = 'b111111001;
    x_128 = 'b111110110;
    x_129 = 'b111011111;
    x_130 = 'b111010000;
    x_131 = 'b111000111;
    x_132 = 'b111001000;
    x_133 = 'b111001010;
    x_134 = 'b111011001;
    x_135 = 'b000000000;
    x_136 = 'b111011010;
    x_137 = 'b111011000;
    x_138 = 'b111010101;
    x_139 = 'b111001001;
    x_140 = 'b111010010;
    x_141 = 'b111001100;
    x_142 = 'b111110001;
    x_143 = 'b111100100;
    x_144 = 'b111011100;
    x_145 = 'b111010101;
    x_146 = 'b111011011;
    x_147 = 'b111011001;
    x_148 = 'b111010011;
    x_149 = 'b111101100;
    x_150 = 'b111100001;
    x_151 = 'b111100000;
    x_152 = 'b000000001;
    x_153 = 'b000000000;
    x_154 = 'b111001100;
    x_155 = 'b111001100;
    x_156 = 'b111011111;
    x_157 = 'b000000011;
    x_158 = 'b111110110;
    x_159 = 'b111001111;
    x_160 = 'b111001101;
    x_161 = 'b111001000;
    x_162 = 'b111000111;
    x_163 = 'b111010010;
    x_164 = 'b111010011;
    x_165 = 'b111111001;
    x_166 = 'b111111011;
    x_167 = 'b111011001;
    x_168 = 'b111111101;
    x_169 = 'b111011111;
    x_170 = 'b111110101;
    x_171 = 'b111011101;
    x_172 = 'b000000010;
    x_173 = 'b111101001;
    x_174 = 'b111110011;
    x_175 = 'b111110000;
    x_176 = 'b111100111;
    x_177 = 'b111101001;
    x_178 = 'b111100011;
    x_179 = 'b111101100;
    x_180 = 'b111110000;
    x_181 = 'b111111011;
    x_182 = 'b111111100;
    x_183 = 'b111110000;
    x_184 = 'b111101010;
    x_185 = 'b111110101;
    x_186 = 'b111111111;
    x_187 = 'b000001100;
    x_188 = 'b111100100;
    x_189 = 'b111100110;
    x_190 = 'b111101001;
    x_191 = 'b111111001;
    x_192 = 'b111110110;
    x_193 = 'b111011111;
    x_194 = 'b111010000;
    x_195 = 'b111000111;
    x_196 = 'b111001000;
    x_197 = 'b111001010;
    x_198 = 'b111011001;
    x_199 = 'b000000000;
    x_200 = 'b111011010;
    x_201 = 'b111011000;
    x_202 = 'b111010101;
    x_203 = 'b111001001;
    x_204 = 'b111010010;
    x_205 = 'b111001100;
    x_206 = 'b111110001;
    x_207 = 'b111100100;
    x_208 = 'b111011100;
    x_209 = 'b111010101;
    x_210 = 'b111011011;
    x_211 = 'b111011001;
    x_212 = 'b111010011;
    x_213 = 'b111101100;
    x_214 = 'b111100001;
    x_215 = 'b111100000;
    x_216 = 'b000000001;
    x_217 = 'b000000000;
    x_218 = 'b111001100;
    x_219 = 'b111001100;
    x_220 = 'b111011111;
    x_221 = 'b000000011;
    x_222 = 'b111110110;
    x_223 = 'b111001111;
    x_224 = 'b111001101;
    x_225 = 'b111001000;
    x_226 = 'b111000111;
    x_227 = 'b111010010;
    x_228 = 'b111010011;
    x_229 = 'b111111001;
    x_230 = 'b111111011;
    x_231 = 'b111011001;
    x_232 = 'b111111101;
    x_233 = 'b111011111;
    x_234 = 'b111110101;
    x_235 = 'b111011101;
    x_236 = 'b000000010;
    x_237 = 'b111101001;
    x_238 = 'b111110011;
    x_239 = 'b111110000;
    x_240 = 'b111100111;
    x_241 = 'b111101001;
    x_242 = 'b111100011;
    x_243 = 'b111101100;
    x_244 = 'b111110000;
    x_245 = 'b111111011;
    x_246 = 'b111111100;
    x_247 = 'b111110000;
    x_248 = 'b111101010;
    x_249 = 'b111110101;
    x_250 = 'b111111111;
    x_251 = 'b000001100;
    x_252 = 'b111100100;
    x_253 = 'b111100110;
    x_254 = 'b111101001;
    x_255 = 'b111111001;

    h_0 = 'b111110110;
    h_1 = 'b111011111;
    h_2 = 'b111010000;
    h_3 = 'b111000111;
    h_4 = 'b111001000;
    h_5 = 'b111001010;
    h_6 = 'b111011001;
    h_7 = 'b000000000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111101111;
    x_1 = 'b111011011;
    x_2 = 'b111001101;
    x_3 = 'b111000011;
    x_4 = 'b111001000;
    x_5 = 'b111001001;
    x_6 = 'b111011000;
    x_7 = 'b111111011;
    x_8 = 'b111011010;
    x_9 = 'b111011000;
    x_10 = 'b111010111;
    x_11 = 'b111001011;
    x_12 = 'b111010101;
    x_13 = 'b111010000;
    x_14 = 'b111110000;
    x_15 = 'b111101000;
    x_16 = 'b111100010;
    x_17 = 'b111010111;
    x_18 = 'b111100011;
    x_19 = 'b111100001;
    x_20 = 'b111011010;
    x_21 = 'b111101010;
    x_22 = 'b111011100;
    x_23 = 'b111011011;
    x_24 = 'b111111011;
    x_25 = 'b111111011;
    x_26 = 'b111000101;
    x_27 = 'b111000101;
    x_28 = 'b111011001;
    x_29 = 'b111110111;
    x_30 = 'b111101110;
    x_31 = 'b111000111;
    x_32 = 'b111001000;
    x_33 = 'b111000010;
    x_34 = 'b111000010;
    x_35 = 'b111001011;
    x_36 = 'b111001010;
    x_37 = 'b111101110;
    x_38 = 'b111111010;
    x_39 = 'b111001011;
    x_40 = 'b111110011;
    x_41 = 'b110110111;
    x_42 = 'b111111000;
    x_43 = 'b111101010;
    x_44 = 'b000000001;
    x_45 = 'b111111010;
    x_46 = 'b111110010;
    x_47 = 'b111110101;
    x_48 = 'b111110000;
    x_49 = 'b111110010;
    x_50 = 'b111101010;
    x_51 = 'b111111101;
    x_52 = 'b000000010;
    x_53 = 'b000010010;
    x_54 = 'b000011001;
    x_55 = 'b111111110;
    x_56 = 'b111110111;
    x_57 = 'b000000011;
    x_58 = 'b000011111;
    x_59 = 'b000110100;
    x_60 = 'b111111001;
    x_61 = 'b000000111;
    x_62 = 'b000011000;
    x_63 = 'b000010100;
    x_64 = 'b111101111;
    x_65 = 'b111011011;
    x_66 = 'b111001101;
    x_67 = 'b111000011;
    x_68 = 'b111001000;
    x_69 = 'b111001001;
    x_70 = 'b111011000;
    x_71 = 'b111111011;
    x_72 = 'b111011010;
    x_73 = 'b111011000;
    x_74 = 'b111010111;
    x_75 = 'b111001011;
    x_76 = 'b111010101;
    x_77 = 'b111010000;
    x_78 = 'b111110000;
    x_79 = 'b111101000;
    x_80 = 'b111100010;
    x_81 = 'b111010111;
    x_82 = 'b111100011;
    x_83 = 'b111100001;
    x_84 = 'b111011010;
    x_85 = 'b111101010;
    x_86 = 'b111011100;
    x_87 = 'b111011011;
    x_88 = 'b111111011;
    x_89 = 'b111111011;
    x_90 = 'b111000101;
    x_91 = 'b111000101;
    x_92 = 'b111011001;
    x_93 = 'b111110111;
    x_94 = 'b111101110;
    x_95 = 'b111000111;
    x_96 = 'b111001000;
    x_97 = 'b111000010;
    x_98 = 'b111000010;
    x_99 = 'b111001011;
    x_100 = 'b111001010;
    x_101 = 'b111101110;
    x_102 = 'b111111010;
    x_103 = 'b111001011;
    x_104 = 'b111110011;
    x_105 = 'b110110111;
    x_106 = 'b111111000;
    x_107 = 'b111101010;
    x_108 = 'b000000001;
    x_109 = 'b111111010;
    x_110 = 'b111110010;
    x_111 = 'b111110101;
    x_112 = 'b111110000;
    x_113 = 'b111110010;
    x_114 = 'b111101010;
    x_115 = 'b111111101;
    x_116 = 'b000000010;
    x_117 = 'b000010010;
    x_118 = 'b000011001;
    x_119 = 'b111111110;
    x_120 = 'b111110111;
    x_121 = 'b000000011;
    x_122 = 'b000011111;
    x_123 = 'b000110100;
    x_124 = 'b111111001;
    x_125 = 'b000000111;
    x_126 = 'b000011000;
    x_127 = 'b000010100;
    x_128 = 'b111101111;
    x_129 = 'b111011011;
    x_130 = 'b111001101;
    x_131 = 'b111000011;
    x_132 = 'b111001000;
    x_133 = 'b111001001;
    x_134 = 'b111011000;
    x_135 = 'b111111011;
    x_136 = 'b111011010;
    x_137 = 'b111011000;
    x_138 = 'b111010111;
    x_139 = 'b111001011;
    x_140 = 'b111010101;
    x_141 = 'b111010000;
    x_142 = 'b111110000;
    x_143 = 'b111101000;
    x_144 = 'b111100010;
    x_145 = 'b111010111;
    x_146 = 'b111100011;
    x_147 = 'b111100001;
    x_148 = 'b111011010;
    x_149 = 'b111101010;
    x_150 = 'b111011100;
    x_151 = 'b111011011;
    x_152 = 'b111111011;
    x_153 = 'b111111011;
    x_154 = 'b111000101;
    x_155 = 'b111000101;
    x_156 = 'b111011001;
    x_157 = 'b111110111;
    x_158 = 'b111101110;
    x_159 = 'b111000111;
    x_160 = 'b111001000;
    x_161 = 'b111000010;
    x_162 = 'b111000010;
    x_163 = 'b111001011;
    x_164 = 'b111001010;
    x_165 = 'b111101110;
    x_166 = 'b111111010;
    x_167 = 'b111001011;
    x_168 = 'b111110011;
    x_169 = 'b110110111;
    x_170 = 'b111111000;
    x_171 = 'b111101010;
    x_172 = 'b000000001;
    x_173 = 'b111111010;
    x_174 = 'b111110010;
    x_175 = 'b111110101;
    x_176 = 'b111110000;
    x_177 = 'b111110010;
    x_178 = 'b111101010;
    x_179 = 'b111111101;
    x_180 = 'b000000010;
    x_181 = 'b000010010;
    x_182 = 'b000011001;
    x_183 = 'b111111110;
    x_184 = 'b111110111;
    x_185 = 'b000000011;
    x_186 = 'b000011111;
    x_187 = 'b000110100;
    x_188 = 'b111111001;
    x_189 = 'b000000111;
    x_190 = 'b000011000;
    x_191 = 'b000010100;
    x_192 = 'b111101111;
    x_193 = 'b111011011;
    x_194 = 'b111001101;
    x_195 = 'b111000011;
    x_196 = 'b111001000;
    x_197 = 'b111001001;
    x_198 = 'b111011000;
    x_199 = 'b111111011;
    x_200 = 'b111011010;
    x_201 = 'b111011000;
    x_202 = 'b111010111;
    x_203 = 'b111001011;
    x_204 = 'b111010101;
    x_205 = 'b111010000;
    x_206 = 'b111110000;
    x_207 = 'b111101000;
    x_208 = 'b111100010;
    x_209 = 'b111010111;
    x_210 = 'b111100011;
    x_211 = 'b111100001;
    x_212 = 'b111011010;
    x_213 = 'b111101010;
    x_214 = 'b111011100;
    x_215 = 'b111011011;
    x_216 = 'b111111011;
    x_217 = 'b111111011;
    x_218 = 'b111000101;
    x_219 = 'b111000101;
    x_220 = 'b111011001;
    x_221 = 'b111110111;
    x_222 = 'b111101110;
    x_223 = 'b111000111;
    x_224 = 'b111001000;
    x_225 = 'b111000010;
    x_226 = 'b111000010;
    x_227 = 'b111001011;
    x_228 = 'b111001010;
    x_229 = 'b111101110;
    x_230 = 'b111111010;
    x_231 = 'b111001011;
    x_232 = 'b111110011;
    x_233 = 'b110110111;
    x_234 = 'b111111000;
    x_235 = 'b111101010;
    x_236 = 'b000000001;
    x_237 = 'b111111010;
    x_238 = 'b111110010;
    x_239 = 'b111110101;
    x_240 = 'b111110000;
    x_241 = 'b111110010;
    x_242 = 'b111101010;
    x_243 = 'b111111101;
    x_244 = 'b000000010;
    x_245 = 'b000010010;
    x_246 = 'b000011001;
    x_247 = 'b111111110;
    x_248 = 'b111110111;
    x_249 = 'b000000011;
    x_250 = 'b000011111;
    x_251 = 'b000110100;
    x_252 = 'b111111001;
    x_253 = 'b000000111;
    x_254 = 'b000011000;
    x_255 = 'b000010100;

    h_0 = 'b111101111;
    h_1 = 'b111011011;
    h_2 = 'b111001101;
    h_3 = 'b111000011;
    h_4 = 'b111001000;
    h_5 = 'b111001001;
    h_6 = 'b111011000;
    h_7 = 'b111111011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111101110;
    x_1 = 'b111100000;
    x_2 = 'b111001101;
    x_3 = 'b111000011;
    x_4 = 'b111000110;
    x_5 = 'b111000101;
    x_6 = 'b111001101;
    x_7 = 'b111111010;
    x_8 = 'b111011111;
    x_9 = 'b111011011;
    x_10 = 'b111011010;
    x_11 = 'b111001110;
    x_12 = 'b111010011;
    x_13 = 'b111000101;
    x_14 = 'b111110100;
    x_15 = 'b111101100;
    x_16 = 'b111100111;
    x_17 = 'b111011010;
    x_18 = 'b111100111;
    x_19 = 'b111100111;
    x_20 = 'b111100000;
    x_21 = 'b111101111;
    x_22 = 'b111100001;
    x_23 = 'b111100001;
    x_24 = 'b000000001;
    x_25 = 'b000000000;
    x_26 = 'b111001101;
    x_27 = 'b111001011;
    x_28 = 'b111011101;
    x_29 = 'b000000000;
    x_30 = 'b111110101;
    x_31 = 'b111010000;
    x_32 = 'b111010001;
    x_33 = 'b111000111;
    x_34 = 'b111000110;
    x_35 = 'b111010010;
    x_36 = 'b111001010;
    x_37 = 'b111101011;
    x_38 = 'b000000100;
    x_39 = 'b111000110;
    x_40 = 'b000000101;
    x_41 = 'b110111000;
    x_42 = 'b000010101;
    x_43 = 'b111100001;
    x_44 = 'b000010101;
    x_45 = 'b000010000;
    x_46 = 'b000000011;
    x_47 = 'b000000001;
    x_48 = 'b111111001;
    x_49 = 'b111110100;
    x_50 = 'b111101011;
    x_51 = 'b000000001;
    x_52 = 'b000001010;
    x_53 = 'b000011110;
    x_54 = 'b000101000;
    x_55 = 'b000001111;
    x_56 = 'b000000010;
    x_57 = 'b000000011;
    x_58 = 'b000101001;
    x_59 = 'b001000100;
    x_60 = 'b000001110;
    x_61 = 'b000100000;
    x_62 = 'b000111101;
    x_63 = 'b000101001;
    x_64 = 'b111101110;
    x_65 = 'b111100000;
    x_66 = 'b111001101;
    x_67 = 'b111000011;
    x_68 = 'b111000110;
    x_69 = 'b111000101;
    x_70 = 'b111001101;
    x_71 = 'b111111010;
    x_72 = 'b111011111;
    x_73 = 'b111011011;
    x_74 = 'b111011010;
    x_75 = 'b111001110;
    x_76 = 'b111010011;
    x_77 = 'b111000101;
    x_78 = 'b111110100;
    x_79 = 'b111101100;
    x_80 = 'b111100111;
    x_81 = 'b111011010;
    x_82 = 'b111100111;
    x_83 = 'b111100111;
    x_84 = 'b111100000;
    x_85 = 'b111101111;
    x_86 = 'b111100001;
    x_87 = 'b111100001;
    x_88 = 'b000000001;
    x_89 = 'b000000000;
    x_90 = 'b111001101;
    x_91 = 'b111001011;
    x_92 = 'b111011101;
    x_93 = 'b000000000;
    x_94 = 'b111110101;
    x_95 = 'b111010000;
    x_96 = 'b111010001;
    x_97 = 'b111000111;
    x_98 = 'b111000110;
    x_99 = 'b111010010;
    x_100 = 'b111001010;
    x_101 = 'b111101011;
    x_102 = 'b000000100;
    x_103 = 'b111000110;
    x_104 = 'b000000101;
    x_105 = 'b110111000;
    x_106 = 'b000010101;
    x_107 = 'b111100001;
    x_108 = 'b000010101;
    x_109 = 'b000010000;
    x_110 = 'b000000011;
    x_111 = 'b000000001;
    x_112 = 'b111111001;
    x_113 = 'b111110100;
    x_114 = 'b111101011;
    x_115 = 'b000000001;
    x_116 = 'b000001010;
    x_117 = 'b000011110;
    x_118 = 'b000101000;
    x_119 = 'b000001111;
    x_120 = 'b000000010;
    x_121 = 'b000000011;
    x_122 = 'b000101001;
    x_123 = 'b001000100;
    x_124 = 'b000001110;
    x_125 = 'b000100000;
    x_126 = 'b000111101;
    x_127 = 'b000101001;
    x_128 = 'b111101110;
    x_129 = 'b111100000;
    x_130 = 'b111001101;
    x_131 = 'b111000011;
    x_132 = 'b111000110;
    x_133 = 'b111000101;
    x_134 = 'b111001101;
    x_135 = 'b111111010;
    x_136 = 'b111011111;
    x_137 = 'b111011011;
    x_138 = 'b111011010;
    x_139 = 'b111001110;
    x_140 = 'b111010011;
    x_141 = 'b111000101;
    x_142 = 'b111110100;
    x_143 = 'b111101100;
    x_144 = 'b111100111;
    x_145 = 'b111011010;
    x_146 = 'b111100111;
    x_147 = 'b111100111;
    x_148 = 'b111100000;
    x_149 = 'b111101111;
    x_150 = 'b111100001;
    x_151 = 'b111100001;
    x_152 = 'b000000001;
    x_153 = 'b000000000;
    x_154 = 'b111001101;
    x_155 = 'b111001011;
    x_156 = 'b111011101;
    x_157 = 'b000000000;
    x_158 = 'b111110101;
    x_159 = 'b111010000;
    x_160 = 'b111010001;
    x_161 = 'b111000111;
    x_162 = 'b111000110;
    x_163 = 'b111010010;
    x_164 = 'b111001010;
    x_165 = 'b111101011;
    x_166 = 'b000000100;
    x_167 = 'b111000110;
    x_168 = 'b000000101;
    x_169 = 'b110111000;
    x_170 = 'b000010101;
    x_171 = 'b111100001;
    x_172 = 'b000010101;
    x_173 = 'b000010000;
    x_174 = 'b000000011;
    x_175 = 'b000000001;
    x_176 = 'b111111001;
    x_177 = 'b111110100;
    x_178 = 'b111101011;
    x_179 = 'b000000001;
    x_180 = 'b000001010;
    x_181 = 'b000011110;
    x_182 = 'b000101000;
    x_183 = 'b000001111;
    x_184 = 'b000000010;
    x_185 = 'b000000011;
    x_186 = 'b000101001;
    x_187 = 'b001000100;
    x_188 = 'b000001110;
    x_189 = 'b000100000;
    x_190 = 'b000111101;
    x_191 = 'b000101001;
    x_192 = 'b111101110;
    x_193 = 'b111100000;
    x_194 = 'b111001101;
    x_195 = 'b111000011;
    x_196 = 'b111000110;
    x_197 = 'b111000101;
    x_198 = 'b111001101;
    x_199 = 'b111111010;
    x_200 = 'b111011111;
    x_201 = 'b111011011;
    x_202 = 'b111011010;
    x_203 = 'b111001110;
    x_204 = 'b111010011;
    x_205 = 'b111000101;
    x_206 = 'b111110100;
    x_207 = 'b111101100;
    x_208 = 'b111100111;
    x_209 = 'b111011010;
    x_210 = 'b111100111;
    x_211 = 'b111100111;
    x_212 = 'b111100000;
    x_213 = 'b111101111;
    x_214 = 'b111100001;
    x_215 = 'b111100001;
    x_216 = 'b000000001;
    x_217 = 'b000000000;
    x_218 = 'b111001101;
    x_219 = 'b111001011;
    x_220 = 'b111011101;
    x_221 = 'b000000000;
    x_222 = 'b111110101;
    x_223 = 'b111010000;
    x_224 = 'b111010001;
    x_225 = 'b111000111;
    x_226 = 'b111000110;
    x_227 = 'b111010010;
    x_228 = 'b111001010;
    x_229 = 'b111101011;
    x_230 = 'b000000100;
    x_231 = 'b111000110;
    x_232 = 'b000000101;
    x_233 = 'b110111000;
    x_234 = 'b000010101;
    x_235 = 'b111100001;
    x_236 = 'b000010101;
    x_237 = 'b000010000;
    x_238 = 'b000000011;
    x_239 = 'b000000001;
    x_240 = 'b111111001;
    x_241 = 'b111110100;
    x_242 = 'b111101011;
    x_243 = 'b000000001;
    x_244 = 'b000001010;
    x_245 = 'b000011110;
    x_246 = 'b000101000;
    x_247 = 'b000001111;
    x_248 = 'b000000010;
    x_249 = 'b000000011;
    x_250 = 'b000101001;
    x_251 = 'b001000100;
    x_252 = 'b000001110;
    x_253 = 'b000100000;
    x_254 = 'b000111101;
    x_255 = 'b000101001;

    h_0 = 'b111101110;
    h_1 = 'b111100000;
    h_2 = 'b111001101;
    h_3 = 'b111000011;
    h_4 = 'b111000110;
    h_5 = 'b111000101;
    h_6 = 'b111001101;
    h_7 = 'b111111010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111111101;
    x_1 = 'b111110000;
    x_2 = 'b111011010;
    x_3 = 'b111001111;
    x_4 = 'b111001011;
    x_5 = 'b111001001;
    x_6 = 'b111010010;
    x_7 = 'b000001000;
    x_8 = 'b111101010;
    x_9 = 'b111100010;
    x_10 = 'b111011111;
    x_11 = 'b111010001;
    x_12 = 'b111011001;
    x_13 = 'b111001111;
    x_14 = 'b000000000;
    x_15 = 'b111110000;
    x_16 = 'b111101001;
    x_17 = 'b111011101;
    x_18 = 'b111101001;
    x_19 = 'b111101100;
    x_20 = 'b111101010;
    x_21 = 'b111110001;
    x_22 = 'b111100000;
    x_23 = 'b111011111;
    x_24 = 'b000000100;
    x_25 = 'b000000010;
    x_26 = 'b111010000;
    x_27 = 'b111001000;
    x_28 = 'b111011000;
    x_29 = 'b000000101;
    x_30 = 'b111111011;
    x_31 = 'b111001110;
    x_32 = 'b111010111;
    x_33 = 'b111001100;
    x_34 = 'b111000110;
    x_35 = 'b111010010;
    x_36 = 'b111000100;
    x_37 = 'b111101000;
    x_38 = 'b000000110;
    x_39 = 'b111000111;
    x_40 = 'b000010011;
    x_41 = 'b111001001;
    x_42 = 'b000010010;
    x_43 = 'b111011111;
    x_44 = 'b000010110;
    x_45 = 'b111111100;
    x_46 = 'b000001010;
    x_47 = 'b000000011;
    x_48 = 'b111111000;
    x_49 = 'b111110010;
    x_50 = 'b111101000;
    x_51 = 'b000000001;
    x_52 = 'b000001011;
    x_53 = 'b000011110;
    x_54 = 'b000100101;
    x_55 = 'b000010101;
    x_56 = 'b000000100;
    x_57 = 'b000000010;
    x_58 = 'b000101011;
    x_59 = 'b001000111;
    x_60 = 'b000011011;
    x_61 = 'b000100111;
    x_62 = 'b001001010;
    x_63 = 'b000101011;
    x_64 = 'b111111101;
    x_65 = 'b111110000;
    x_66 = 'b111011010;
    x_67 = 'b111001111;
    x_68 = 'b111001011;
    x_69 = 'b111001001;
    x_70 = 'b111010010;
    x_71 = 'b000001000;
    x_72 = 'b111101010;
    x_73 = 'b111100010;
    x_74 = 'b111011111;
    x_75 = 'b111010001;
    x_76 = 'b111011001;
    x_77 = 'b111001111;
    x_78 = 'b000000000;
    x_79 = 'b111110000;
    x_80 = 'b111101001;
    x_81 = 'b111011101;
    x_82 = 'b111101001;
    x_83 = 'b111101100;
    x_84 = 'b111101010;
    x_85 = 'b111110001;
    x_86 = 'b111100000;
    x_87 = 'b111011111;
    x_88 = 'b000000100;
    x_89 = 'b000000010;
    x_90 = 'b111010000;
    x_91 = 'b111001000;
    x_92 = 'b111011000;
    x_93 = 'b000000101;
    x_94 = 'b111111011;
    x_95 = 'b111001110;
    x_96 = 'b111010111;
    x_97 = 'b111001100;
    x_98 = 'b111000110;
    x_99 = 'b111010010;
    x_100 = 'b111000100;
    x_101 = 'b111101000;
    x_102 = 'b000000110;
    x_103 = 'b111000111;
    x_104 = 'b000010011;
    x_105 = 'b111001001;
    x_106 = 'b000010010;
    x_107 = 'b111011111;
    x_108 = 'b000010110;
    x_109 = 'b111111100;
    x_110 = 'b000001010;
    x_111 = 'b000000011;
    x_112 = 'b111111000;
    x_113 = 'b111110010;
    x_114 = 'b111101000;
    x_115 = 'b000000001;
    x_116 = 'b000001011;
    x_117 = 'b000011110;
    x_118 = 'b000100101;
    x_119 = 'b000010101;
    x_120 = 'b000000100;
    x_121 = 'b000000010;
    x_122 = 'b000101011;
    x_123 = 'b001000111;
    x_124 = 'b000011011;
    x_125 = 'b000100111;
    x_126 = 'b001001010;
    x_127 = 'b000101011;
    x_128 = 'b111111101;
    x_129 = 'b111110000;
    x_130 = 'b111011010;
    x_131 = 'b111001111;
    x_132 = 'b111001011;
    x_133 = 'b111001001;
    x_134 = 'b111010010;
    x_135 = 'b000001000;
    x_136 = 'b111101010;
    x_137 = 'b111100010;
    x_138 = 'b111011111;
    x_139 = 'b111010001;
    x_140 = 'b111011001;
    x_141 = 'b111001111;
    x_142 = 'b000000000;
    x_143 = 'b111110000;
    x_144 = 'b111101001;
    x_145 = 'b111011101;
    x_146 = 'b111101001;
    x_147 = 'b111101100;
    x_148 = 'b111101010;
    x_149 = 'b111110001;
    x_150 = 'b111100000;
    x_151 = 'b111011111;
    x_152 = 'b000000100;
    x_153 = 'b000000010;
    x_154 = 'b111010000;
    x_155 = 'b111001000;
    x_156 = 'b111011000;
    x_157 = 'b000000101;
    x_158 = 'b111111011;
    x_159 = 'b111001110;
    x_160 = 'b111010111;
    x_161 = 'b111001100;
    x_162 = 'b111000110;
    x_163 = 'b111010010;
    x_164 = 'b111000100;
    x_165 = 'b111101000;
    x_166 = 'b000000110;
    x_167 = 'b111000111;
    x_168 = 'b000010011;
    x_169 = 'b111001001;
    x_170 = 'b000010010;
    x_171 = 'b111011111;
    x_172 = 'b000010110;
    x_173 = 'b111111100;
    x_174 = 'b000001010;
    x_175 = 'b000000011;
    x_176 = 'b111111000;
    x_177 = 'b111110010;
    x_178 = 'b111101000;
    x_179 = 'b000000001;
    x_180 = 'b000001011;
    x_181 = 'b000011110;
    x_182 = 'b000100101;
    x_183 = 'b000010101;
    x_184 = 'b000000100;
    x_185 = 'b000000010;
    x_186 = 'b000101011;
    x_187 = 'b001000111;
    x_188 = 'b000011011;
    x_189 = 'b000100111;
    x_190 = 'b001001010;
    x_191 = 'b000101011;
    x_192 = 'b111111101;
    x_193 = 'b111110000;
    x_194 = 'b111011010;
    x_195 = 'b111001111;
    x_196 = 'b111001011;
    x_197 = 'b111001001;
    x_198 = 'b111010010;
    x_199 = 'b000001000;
    x_200 = 'b111101010;
    x_201 = 'b111100010;
    x_202 = 'b111011111;
    x_203 = 'b111010001;
    x_204 = 'b111011001;
    x_205 = 'b111001111;
    x_206 = 'b000000000;
    x_207 = 'b111110000;
    x_208 = 'b111101001;
    x_209 = 'b111011101;
    x_210 = 'b111101001;
    x_211 = 'b111101100;
    x_212 = 'b111101010;
    x_213 = 'b111110001;
    x_214 = 'b111100000;
    x_215 = 'b111011111;
    x_216 = 'b000000100;
    x_217 = 'b000000010;
    x_218 = 'b111010000;
    x_219 = 'b111001000;
    x_220 = 'b111011000;
    x_221 = 'b000000101;
    x_222 = 'b111111011;
    x_223 = 'b111001110;
    x_224 = 'b111010111;
    x_225 = 'b111001100;
    x_226 = 'b111000110;
    x_227 = 'b111010010;
    x_228 = 'b111000100;
    x_229 = 'b111101000;
    x_230 = 'b000000110;
    x_231 = 'b111000111;
    x_232 = 'b000010011;
    x_233 = 'b111001001;
    x_234 = 'b000010010;
    x_235 = 'b111011111;
    x_236 = 'b000010110;
    x_237 = 'b111111100;
    x_238 = 'b000001010;
    x_239 = 'b000000011;
    x_240 = 'b111111000;
    x_241 = 'b111110010;
    x_242 = 'b111101000;
    x_243 = 'b000000001;
    x_244 = 'b000001011;
    x_245 = 'b000011110;
    x_246 = 'b000100101;
    x_247 = 'b000010101;
    x_248 = 'b000000100;
    x_249 = 'b000000010;
    x_250 = 'b000101011;
    x_251 = 'b001000111;
    x_252 = 'b000011011;
    x_253 = 'b000100111;
    x_254 = 'b001001010;
    x_255 = 'b000101011;

    h_0 = 'b111111101;
    h_1 = 'b111110000;
    h_2 = 'b111011010;
    h_3 = 'b111001111;
    h_4 = 'b111001011;
    h_5 = 'b111001001;
    h_6 = 'b111010010;
    h_7 = 'b000001000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111111101;
    x_1 = 'b111101011;
    x_2 = 'b111010111;
    x_3 = 'b111001010;
    x_4 = 'b111000101;
    x_5 = 'b111000010;
    x_6 = 'b111001000;
    x_7 = 'b000000110;
    x_8 = 'b111100110;
    x_9 = 'b111100000;
    x_10 = 'b111011111;
    x_11 = 'b111001101;
    x_12 = 'b111010111;
    x_13 = 'b111010000;
    x_14 = 'b000000001;
    x_15 = 'b111101101;
    x_16 = 'b111101000;
    x_17 = 'b111011111;
    x_18 = 'b111101101;
    x_19 = 'b111110000;
    x_20 = 'b111110000;
    x_21 = 'b111101000;
    x_22 = 'b111010110;
    x_23 = 'b111010100;
    x_24 = 'b111111101;
    x_25 = 'b111111011;
    x_26 = 'b111000101;
    x_27 = 'b110111011;
    x_28 = 'b111001110;
    x_29 = 'b000001010;
    x_30 = 'b111110010;
    x_31 = 'b111000111;
    x_32 = 'b111001111;
    x_33 = 'b111000011;
    x_34 = 'b110111011;
    x_35 = 'b111000110;
    x_36 = 'b110111100;
    x_37 = 'b111100111;
    x_38 = 'b000001100;
    x_39 = 'b110111111;
    x_40 = 'b000010101;
    x_41 = 'b111000110;
    x_42 = 'b000001110;
    x_43 = 'b000010000;
    x_44 = 'b000100000;
    x_45 = 'b000001110;
    x_46 = 'b000011011;
    x_47 = 'b000010010;
    x_48 = 'b000000100;
    x_49 = 'b111111111;
    x_50 = 'b111110110;
    x_51 = 'b000001111;
    x_52 = 'b000011000;
    x_53 = 'b000101100;
    x_54 = 'b000110011;
    x_55 = 'b000101001;
    x_56 = 'b000010110;
    x_57 = 'b000001111;
    x_58 = 'b000110101;
    x_59 = 'b001001011;
    x_60 = 'b000100110;
    x_61 = 'b000101000;
    x_62 = 'b001001001;
    x_63 = 'b000101101;
    x_64 = 'b111111101;
    x_65 = 'b111101011;
    x_66 = 'b111010111;
    x_67 = 'b111001010;
    x_68 = 'b111000101;
    x_69 = 'b111000010;
    x_70 = 'b111001000;
    x_71 = 'b000000110;
    x_72 = 'b111100110;
    x_73 = 'b111100000;
    x_74 = 'b111011111;
    x_75 = 'b111001101;
    x_76 = 'b111010111;
    x_77 = 'b111010000;
    x_78 = 'b000000001;
    x_79 = 'b111101101;
    x_80 = 'b111101000;
    x_81 = 'b111011111;
    x_82 = 'b111101101;
    x_83 = 'b111110000;
    x_84 = 'b111110000;
    x_85 = 'b111101000;
    x_86 = 'b111010110;
    x_87 = 'b111010100;
    x_88 = 'b111111101;
    x_89 = 'b111111011;
    x_90 = 'b111000101;
    x_91 = 'b110111011;
    x_92 = 'b111001110;
    x_93 = 'b000001010;
    x_94 = 'b111110010;
    x_95 = 'b111000111;
    x_96 = 'b111001111;
    x_97 = 'b111000011;
    x_98 = 'b110111011;
    x_99 = 'b111000110;
    x_100 = 'b110111100;
    x_101 = 'b111100111;
    x_102 = 'b000001100;
    x_103 = 'b110111111;
    x_104 = 'b000010101;
    x_105 = 'b111000110;
    x_106 = 'b000001110;
    x_107 = 'b000010000;
    x_108 = 'b000100000;
    x_109 = 'b000001110;
    x_110 = 'b000011011;
    x_111 = 'b000010010;
    x_112 = 'b000000100;
    x_113 = 'b111111111;
    x_114 = 'b111110110;
    x_115 = 'b000001111;
    x_116 = 'b000011000;
    x_117 = 'b000101100;
    x_118 = 'b000110011;
    x_119 = 'b000101001;
    x_120 = 'b000010110;
    x_121 = 'b000001111;
    x_122 = 'b000110101;
    x_123 = 'b001001011;
    x_124 = 'b000100110;
    x_125 = 'b000101000;
    x_126 = 'b001001001;
    x_127 = 'b000101101;
    x_128 = 'b111111101;
    x_129 = 'b111101011;
    x_130 = 'b111010111;
    x_131 = 'b111001010;
    x_132 = 'b111000101;
    x_133 = 'b111000010;
    x_134 = 'b111001000;
    x_135 = 'b000000110;
    x_136 = 'b111100110;
    x_137 = 'b111100000;
    x_138 = 'b111011111;
    x_139 = 'b111001101;
    x_140 = 'b111010111;
    x_141 = 'b111010000;
    x_142 = 'b000000001;
    x_143 = 'b111101101;
    x_144 = 'b111101000;
    x_145 = 'b111011111;
    x_146 = 'b111101101;
    x_147 = 'b111110000;
    x_148 = 'b111110000;
    x_149 = 'b111101000;
    x_150 = 'b111010110;
    x_151 = 'b111010100;
    x_152 = 'b111111101;
    x_153 = 'b111111011;
    x_154 = 'b111000101;
    x_155 = 'b110111011;
    x_156 = 'b111001110;
    x_157 = 'b000001010;
    x_158 = 'b111110010;
    x_159 = 'b111000111;
    x_160 = 'b111001111;
    x_161 = 'b111000011;
    x_162 = 'b110111011;
    x_163 = 'b111000110;
    x_164 = 'b110111100;
    x_165 = 'b111100111;
    x_166 = 'b000001100;
    x_167 = 'b110111111;
    x_168 = 'b000010101;
    x_169 = 'b111000110;
    x_170 = 'b000001110;
    x_171 = 'b000010000;
    x_172 = 'b000100000;
    x_173 = 'b000001110;
    x_174 = 'b000011011;
    x_175 = 'b000010010;
    x_176 = 'b000000100;
    x_177 = 'b111111111;
    x_178 = 'b111110110;
    x_179 = 'b000001111;
    x_180 = 'b000011000;
    x_181 = 'b000101100;
    x_182 = 'b000110011;
    x_183 = 'b000101001;
    x_184 = 'b000010110;
    x_185 = 'b000001111;
    x_186 = 'b000110101;
    x_187 = 'b001001011;
    x_188 = 'b000100110;
    x_189 = 'b000101000;
    x_190 = 'b001001001;
    x_191 = 'b000101101;
    x_192 = 'b111111101;
    x_193 = 'b111101011;
    x_194 = 'b111010111;
    x_195 = 'b111001010;
    x_196 = 'b111000101;
    x_197 = 'b111000010;
    x_198 = 'b111001000;
    x_199 = 'b000000110;
    x_200 = 'b111100110;
    x_201 = 'b111100000;
    x_202 = 'b111011111;
    x_203 = 'b111001101;
    x_204 = 'b111010111;
    x_205 = 'b111010000;
    x_206 = 'b000000001;
    x_207 = 'b111101101;
    x_208 = 'b111101000;
    x_209 = 'b111011111;
    x_210 = 'b111101101;
    x_211 = 'b111110000;
    x_212 = 'b111110000;
    x_213 = 'b111101000;
    x_214 = 'b111010110;
    x_215 = 'b111010100;
    x_216 = 'b111111101;
    x_217 = 'b111111011;
    x_218 = 'b111000101;
    x_219 = 'b110111011;
    x_220 = 'b111001110;
    x_221 = 'b000001010;
    x_222 = 'b111110010;
    x_223 = 'b111000111;
    x_224 = 'b111001111;
    x_225 = 'b111000011;
    x_226 = 'b110111011;
    x_227 = 'b111000110;
    x_228 = 'b110111100;
    x_229 = 'b111100111;
    x_230 = 'b000001100;
    x_231 = 'b110111111;
    x_232 = 'b000010101;
    x_233 = 'b111000110;
    x_234 = 'b000001110;
    x_235 = 'b000010000;
    x_236 = 'b000100000;
    x_237 = 'b000001110;
    x_238 = 'b000011011;
    x_239 = 'b000010010;
    x_240 = 'b000000100;
    x_241 = 'b111111111;
    x_242 = 'b111110110;
    x_243 = 'b000001111;
    x_244 = 'b000011000;
    x_245 = 'b000101100;
    x_246 = 'b000110011;
    x_247 = 'b000101001;
    x_248 = 'b000010110;
    x_249 = 'b000001111;
    x_250 = 'b000110101;
    x_251 = 'b001001011;
    x_252 = 'b000100110;
    x_253 = 'b000101000;
    x_254 = 'b001001001;
    x_255 = 'b000101101;

    h_0 = 'b111111101;
    h_1 = 'b111101011;
    h_2 = 'b111010111;
    h_3 = 'b111001010;
    h_4 = 'b111000101;
    h_5 = 'b111000010;
    h_6 = 'b111001000;
    h_7 = 'b000000110;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000000101;
    x_1 = 'b111110010;
    x_2 = 'b111011100;
    x_3 = 'b111000110;
    x_4 = 'b111000100;
    x_5 = 'b111000010;
    x_6 = 'b111001111;
    x_7 = 'b000010101;
    x_8 = 'b111110011;
    x_9 = 'b111101101;
    x_10 = 'b111101010;
    x_11 = 'b111010100;
    x_12 = 'b111011011;
    x_13 = 'b111011101;
    x_14 = 'b000010011;
    x_15 = 'b000000010;
    x_16 = 'b111111010;
    x_17 = 'b111101110;
    x_18 = 'b111111010;
    x_19 = 'b111111100;
    x_20 = 'b111111110;
    x_21 = 'b111101011;
    x_22 = 'b111011000;
    x_23 = 'b111011000;
    x_24 = 'b111111111;
    x_25 = 'b111111101;
    x_26 = 'b111000110;
    x_27 = 'b110111100;
    x_28 = 'b111010011;
    x_29 = 'b000001001;
    x_30 = 'b111110110;
    x_31 = 'b111000111;
    x_32 = 'b111010010;
    x_33 = 'b111000010;
    x_34 = 'b110111010;
    x_35 = 'b111000110;
    x_36 = 'b111000000;
    x_37 = 'b111110000;
    x_38 = 'b000010001;
    x_39 = 'b111001001;
    x_40 = 'b000001111;
    x_41 = 'b111001001;
    x_42 = 'b000100100;
    x_43 = 'b111110110;
    x_44 = 'b000110110;
    x_45 = 'b000011011;
    x_46 = 'b000110101;
    x_47 = 'b000100010;
    x_48 = 'b000001111;
    x_49 = 'b000001010;
    x_50 = 'b111111111;
    x_51 = 'b000010001;
    x_52 = 'b000010110;
    x_53 = 'b000101000;
    x_54 = 'b000101110;
    x_55 = 'b000111000;
    x_56 = 'b000100001;
    x_57 = 'b000010101;
    x_58 = 'b000101111;
    x_59 = 'b001000001;
    x_60 = 'b000110010;
    x_61 = 'b000101011;
    x_62 = 'b001000011;
    x_63 = 'b000111000;
    x_64 = 'b000000101;
    x_65 = 'b111110010;
    x_66 = 'b111011100;
    x_67 = 'b111000110;
    x_68 = 'b111000100;
    x_69 = 'b111000010;
    x_70 = 'b111001111;
    x_71 = 'b000010101;
    x_72 = 'b111110011;
    x_73 = 'b111101101;
    x_74 = 'b111101010;
    x_75 = 'b111010100;
    x_76 = 'b111011011;
    x_77 = 'b111011101;
    x_78 = 'b000010011;
    x_79 = 'b000000010;
    x_80 = 'b111111010;
    x_81 = 'b111101110;
    x_82 = 'b111111010;
    x_83 = 'b111111100;
    x_84 = 'b111111110;
    x_85 = 'b111101011;
    x_86 = 'b111011000;
    x_87 = 'b111011000;
    x_88 = 'b111111111;
    x_89 = 'b111111101;
    x_90 = 'b111000110;
    x_91 = 'b110111100;
    x_92 = 'b111010011;
    x_93 = 'b000001001;
    x_94 = 'b111110110;
    x_95 = 'b111000111;
    x_96 = 'b111010010;
    x_97 = 'b111000010;
    x_98 = 'b110111010;
    x_99 = 'b111000110;
    x_100 = 'b111000000;
    x_101 = 'b111110000;
    x_102 = 'b000010001;
    x_103 = 'b111001001;
    x_104 = 'b000001111;
    x_105 = 'b111001001;
    x_106 = 'b000100100;
    x_107 = 'b111110110;
    x_108 = 'b000110110;
    x_109 = 'b000011011;
    x_110 = 'b000110101;
    x_111 = 'b000100010;
    x_112 = 'b000001111;
    x_113 = 'b000001010;
    x_114 = 'b111111111;
    x_115 = 'b000010001;
    x_116 = 'b000010110;
    x_117 = 'b000101000;
    x_118 = 'b000101110;
    x_119 = 'b000111000;
    x_120 = 'b000100001;
    x_121 = 'b000010101;
    x_122 = 'b000101111;
    x_123 = 'b001000001;
    x_124 = 'b000110010;
    x_125 = 'b000101011;
    x_126 = 'b001000011;
    x_127 = 'b000111000;
    x_128 = 'b000000101;
    x_129 = 'b111110010;
    x_130 = 'b111011100;
    x_131 = 'b111000110;
    x_132 = 'b111000100;
    x_133 = 'b111000010;
    x_134 = 'b111001111;
    x_135 = 'b000010101;
    x_136 = 'b111110011;
    x_137 = 'b111101101;
    x_138 = 'b111101010;
    x_139 = 'b111010100;
    x_140 = 'b111011011;
    x_141 = 'b111011101;
    x_142 = 'b000010011;
    x_143 = 'b000000010;
    x_144 = 'b111111010;
    x_145 = 'b111101110;
    x_146 = 'b111111010;
    x_147 = 'b111111100;
    x_148 = 'b111111110;
    x_149 = 'b111101011;
    x_150 = 'b111011000;
    x_151 = 'b111011000;
    x_152 = 'b111111111;
    x_153 = 'b111111101;
    x_154 = 'b111000110;
    x_155 = 'b110111100;
    x_156 = 'b111010011;
    x_157 = 'b000001001;
    x_158 = 'b111110110;
    x_159 = 'b111000111;
    x_160 = 'b111010010;
    x_161 = 'b111000010;
    x_162 = 'b110111010;
    x_163 = 'b111000110;
    x_164 = 'b111000000;
    x_165 = 'b111110000;
    x_166 = 'b000010001;
    x_167 = 'b111001001;
    x_168 = 'b000001111;
    x_169 = 'b111001001;
    x_170 = 'b000100100;
    x_171 = 'b111110110;
    x_172 = 'b000110110;
    x_173 = 'b000011011;
    x_174 = 'b000110101;
    x_175 = 'b000100010;
    x_176 = 'b000001111;
    x_177 = 'b000001010;
    x_178 = 'b111111111;
    x_179 = 'b000010001;
    x_180 = 'b000010110;
    x_181 = 'b000101000;
    x_182 = 'b000101110;
    x_183 = 'b000111000;
    x_184 = 'b000100001;
    x_185 = 'b000010101;
    x_186 = 'b000101111;
    x_187 = 'b001000001;
    x_188 = 'b000110010;
    x_189 = 'b000101011;
    x_190 = 'b001000011;
    x_191 = 'b000111000;
    x_192 = 'b000000101;
    x_193 = 'b111110010;
    x_194 = 'b111011100;
    x_195 = 'b111000110;
    x_196 = 'b111000100;
    x_197 = 'b111000010;
    x_198 = 'b111001111;
    x_199 = 'b000010101;
    x_200 = 'b111110011;
    x_201 = 'b111101101;
    x_202 = 'b111101010;
    x_203 = 'b111010100;
    x_204 = 'b111011011;
    x_205 = 'b111011101;
    x_206 = 'b000010011;
    x_207 = 'b000000010;
    x_208 = 'b111111010;
    x_209 = 'b111101110;
    x_210 = 'b111111010;
    x_211 = 'b111111100;
    x_212 = 'b111111110;
    x_213 = 'b111101011;
    x_214 = 'b111011000;
    x_215 = 'b111011000;
    x_216 = 'b111111111;
    x_217 = 'b111111101;
    x_218 = 'b111000110;
    x_219 = 'b110111100;
    x_220 = 'b111010011;
    x_221 = 'b000001001;
    x_222 = 'b111110110;
    x_223 = 'b111000111;
    x_224 = 'b111010010;
    x_225 = 'b111000010;
    x_226 = 'b110111010;
    x_227 = 'b111000110;
    x_228 = 'b111000000;
    x_229 = 'b111110000;
    x_230 = 'b000010001;
    x_231 = 'b111001001;
    x_232 = 'b000001111;
    x_233 = 'b111001001;
    x_234 = 'b000100100;
    x_235 = 'b111110110;
    x_236 = 'b000110110;
    x_237 = 'b000011011;
    x_238 = 'b000110101;
    x_239 = 'b000100010;
    x_240 = 'b000001111;
    x_241 = 'b000001010;
    x_242 = 'b111111111;
    x_243 = 'b000010001;
    x_244 = 'b000010110;
    x_245 = 'b000101000;
    x_246 = 'b000101110;
    x_247 = 'b000111000;
    x_248 = 'b000100001;
    x_249 = 'b000010101;
    x_250 = 'b000101111;
    x_251 = 'b001000001;
    x_252 = 'b000110010;
    x_253 = 'b000101011;
    x_254 = 'b001000011;
    x_255 = 'b000111000;

    h_0 = 'b000000101;
    h_1 = 'b111110010;
    h_2 = 'b111011100;
    h_3 = 'b111000110;
    h_4 = 'b111000100;
    h_5 = 'b111000010;
    h_6 = 'b111001111;
    h_7 = 'b000010101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000000001;
    x_1 = 'b111110111;
    x_2 = 'b111100001;
    x_3 = 'b111001011;
    x_4 = 'b111000001;
    x_5 = 'b110111010;
    x_6 = 'b111001010;
    x_7 = 'b000010100;
    x_8 = 'b111110101;
    x_9 = 'b111110010;
    x_10 = 'b111101011;
    x_11 = 'b111001100;
    x_12 = 'b111001011;
    x_13 = 'b111010000;
    x_14 = 'b000011100;
    x_15 = 'b000000101;
    x_16 = 'b111111100;
    x_17 = 'b111101111;
    x_18 = 'b111110101;
    x_19 = 'b111110001;
    x_20 = 'b111101101;
    x_21 = 'b111101111;
    x_22 = 'b111011100;
    x_23 = 'b111011011;
    x_24 = 'b000000100;
    x_25 = 'b000000010;
    x_26 = 'b111001010;
    x_27 = 'b110111110;
    x_28 = 'b111001111;
    x_29 = 'b000001111;
    x_30 = 'b111111010;
    x_31 = 'b111001010;
    x_32 = 'b111011001;
    x_33 = 'b111001010;
    x_34 = 'b111000000;
    x_35 = 'b111001011;
    x_36 = 'b111000001;
    x_37 = 'b111110000;
    x_38 = 'b000010010;
    x_39 = 'b111001010;
    x_40 = 'b000011011;
    x_41 = 'b111011100;
    x_42 = 'b000101100;
    x_43 = 'b111101011;
    x_44 = 'b000110110;
    x_45 = 'b000000101;
    x_46 = 'b000110000;
    x_47 = 'b000100001;
    x_48 = 'b000001101;
    x_49 = 'b000001001;
    x_50 = 'b111111011;
    x_51 = 'b000000111;
    x_52 = 'b000001011;
    x_53 = 'b000010111;
    x_54 = 'b000011100;
    x_55 = 'b000110111;
    x_56 = 'b000100000;
    x_57 = 'b000010001;
    x_58 = 'b000011110;
    x_59 = 'b000100011;
    x_60 = 'b000110110;
    x_61 = 'b000100011;
    x_62 = 'b000110100;
    x_63 = 'b000110100;
    x_64 = 'b000000001;
    x_65 = 'b111110111;
    x_66 = 'b111100001;
    x_67 = 'b111001011;
    x_68 = 'b111000001;
    x_69 = 'b110111010;
    x_70 = 'b111001010;
    x_71 = 'b000010100;
    x_72 = 'b111110101;
    x_73 = 'b111110010;
    x_74 = 'b111101011;
    x_75 = 'b111001100;
    x_76 = 'b111001011;
    x_77 = 'b111010000;
    x_78 = 'b000011100;
    x_79 = 'b000000101;
    x_80 = 'b111111100;
    x_81 = 'b111101111;
    x_82 = 'b111110101;
    x_83 = 'b111110001;
    x_84 = 'b111101101;
    x_85 = 'b111101111;
    x_86 = 'b111011100;
    x_87 = 'b111011011;
    x_88 = 'b000000100;
    x_89 = 'b000000010;
    x_90 = 'b111001010;
    x_91 = 'b110111110;
    x_92 = 'b111001111;
    x_93 = 'b000001111;
    x_94 = 'b111111010;
    x_95 = 'b111001010;
    x_96 = 'b111011001;
    x_97 = 'b111001010;
    x_98 = 'b111000000;
    x_99 = 'b111001011;
    x_100 = 'b111000001;
    x_101 = 'b111110000;
    x_102 = 'b000010010;
    x_103 = 'b111001010;
    x_104 = 'b000011011;
    x_105 = 'b111011100;
    x_106 = 'b000101100;
    x_107 = 'b111101011;
    x_108 = 'b000110110;
    x_109 = 'b000000101;
    x_110 = 'b000110000;
    x_111 = 'b000100001;
    x_112 = 'b000001101;
    x_113 = 'b000001001;
    x_114 = 'b111111011;
    x_115 = 'b000000111;
    x_116 = 'b000001011;
    x_117 = 'b000010111;
    x_118 = 'b000011100;
    x_119 = 'b000110111;
    x_120 = 'b000100000;
    x_121 = 'b000010001;
    x_122 = 'b000011110;
    x_123 = 'b000100011;
    x_124 = 'b000110110;
    x_125 = 'b000100011;
    x_126 = 'b000110100;
    x_127 = 'b000110100;
    x_128 = 'b000000001;
    x_129 = 'b111110111;
    x_130 = 'b111100001;
    x_131 = 'b111001011;
    x_132 = 'b111000001;
    x_133 = 'b110111010;
    x_134 = 'b111001010;
    x_135 = 'b000010100;
    x_136 = 'b111110101;
    x_137 = 'b111110010;
    x_138 = 'b111101011;
    x_139 = 'b111001100;
    x_140 = 'b111001011;
    x_141 = 'b111010000;
    x_142 = 'b000011100;
    x_143 = 'b000000101;
    x_144 = 'b111111100;
    x_145 = 'b111101111;
    x_146 = 'b111110101;
    x_147 = 'b111110001;
    x_148 = 'b111101101;
    x_149 = 'b111101111;
    x_150 = 'b111011100;
    x_151 = 'b111011011;
    x_152 = 'b000000100;
    x_153 = 'b000000010;
    x_154 = 'b111001010;
    x_155 = 'b110111110;
    x_156 = 'b111001111;
    x_157 = 'b000001111;
    x_158 = 'b111111010;
    x_159 = 'b111001010;
    x_160 = 'b111011001;
    x_161 = 'b111001010;
    x_162 = 'b111000000;
    x_163 = 'b111001011;
    x_164 = 'b111000001;
    x_165 = 'b111110000;
    x_166 = 'b000010010;
    x_167 = 'b111001010;
    x_168 = 'b000011011;
    x_169 = 'b111011100;
    x_170 = 'b000101100;
    x_171 = 'b111101011;
    x_172 = 'b000110110;
    x_173 = 'b000000101;
    x_174 = 'b000110000;
    x_175 = 'b000100001;
    x_176 = 'b000001101;
    x_177 = 'b000001001;
    x_178 = 'b111111011;
    x_179 = 'b000000111;
    x_180 = 'b000001011;
    x_181 = 'b000010111;
    x_182 = 'b000011100;
    x_183 = 'b000110111;
    x_184 = 'b000100000;
    x_185 = 'b000010001;
    x_186 = 'b000011110;
    x_187 = 'b000100011;
    x_188 = 'b000110110;
    x_189 = 'b000100011;
    x_190 = 'b000110100;
    x_191 = 'b000110100;
    x_192 = 'b000000001;
    x_193 = 'b111110111;
    x_194 = 'b111100001;
    x_195 = 'b111001011;
    x_196 = 'b111000001;
    x_197 = 'b110111010;
    x_198 = 'b111001010;
    x_199 = 'b000010100;
    x_200 = 'b111110101;
    x_201 = 'b111110010;
    x_202 = 'b111101011;
    x_203 = 'b111001100;
    x_204 = 'b111001011;
    x_205 = 'b111010000;
    x_206 = 'b000011100;
    x_207 = 'b000000101;
    x_208 = 'b111111100;
    x_209 = 'b111101111;
    x_210 = 'b111110101;
    x_211 = 'b111110001;
    x_212 = 'b111101101;
    x_213 = 'b111101111;
    x_214 = 'b111011100;
    x_215 = 'b111011011;
    x_216 = 'b000000100;
    x_217 = 'b000000010;
    x_218 = 'b111001010;
    x_219 = 'b110111110;
    x_220 = 'b111001111;
    x_221 = 'b000001111;
    x_222 = 'b111111010;
    x_223 = 'b111001010;
    x_224 = 'b111011001;
    x_225 = 'b111001010;
    x_226 = 'b111000000;
    x_227 = 'b111001011;
    x_228 = 'b111000001;
    x_229 = 'b111110000;
    x_230 = 'b000010010;
    x_231 = 'b111001010;
    x_232 = 'b000011011;
    x_233 = 'b111011100;
    x_234 = 'b000101100;
    x_235 = 'b111101011;
    x_236 = 'b000110110;
    x_237 = 'b000000101;
    x_238 = 'b000110000;
    x_239 = 'b000100001;
    x_240 = 'b000001101;
    x_241 = 'b000001001;
    x_242 = 'b111111011;
    x_243 = 'b000000111;
    x_244 = 'b000001011;
    x_245 = 'b000010111;
    x_246 = 'b000011100;
    x_247 = 'b000110111;
    x_248 = 'b000100000;
    x_249 = 'b000010001;
    x_250 = 'b000011110;
    x_251 = 'b000100011;
    x_252 = 'b000110110;
    x_253 = 'b000100011;
    x_254 = 'b000110100;
    x_255 = 'b000110100;

    h_0 = 'b000000001;
    h_1 = 'b111110111;
    h_2 = 'b111100001;
    h_3 = 'b111001011;
    h_4 = 'b111000001;
    h_5 = 'b110111010;
    h_6 = 'b111001010;
    h_7 = 'b000010100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000000111;
    x_1 = 'b111111011;
    x_2 = 'b111100100;
    x_3 = 'b111001111;
    x_4 = 'b111000111;
    x_5 = 'b110111101;
    x_6 = 'b111001011;
    x_7 = 'b000010111;
    x_8 = 'b111110110;
    x_9 = 'b111110001;
    x_10 = 'b111100101;
    x_11 = 'b111001100;
    x_12 = 'b111000111;
    x_13 = 'b111010000;
    x_14 = 'b000010111;
    x_15 = 'b000000011;
    x_16 = 'b111111001;
    x_17 = 'b111101101;
    x_18 = 'b111110001;
    x_19 = 'b111101001;
    x_20 = 'b111100101;
    x_21 = 'b111110101;
    x_22 = 'b111100011;
    x_23 = 'b111100011;
    x_24 = 'b000001000;
    x_25 = 'b000000111;
    x_26 = 'b111010001;
    x_27 = 'b111000111;
    x_28 = 'b111011101;
    x_29 = 'b000010100;
    x_30 = 'b111111011;
    x_31 = 'b111010100;
    x_32 = 'b111011010;
    x_33 = 'b111001101;
    x_34 = 'b111000111;
    x_35 = 'b111010000;
    x_36 = 'b111000111;
    x_37 = 'b111110100;
    x_38 = 'b000011000;
    x_39 = 'b111010101;
    x_40 = 'b000101010;
    x_41 = 'b111101011;
    x_42 = 'b000101110;
    x_43 = 'b111100100;
    x_44 = 'b000110110;
    x_45 = 'b111111110;
    x_46 = 'b000101010;
    x_47 = 'b000011011;
    x_48 = 'b000001010;
    x_49 = 'b000001000;
    x_50 = 'b111111101;
    x_51 = 'b000000101;
    x_52 = 'b000000110;
    x_53 = 'b000001100;
    x_54 = 'b000001101;
    x_55 = 'b000110000;
    x_56 = 'b000011011;
    x_57 = 'b000010000;
    x_58 = 'b000010110;
    x_59 = 'b000010001;
    x_60 = 'b000101111;
    x_61 = 'b000010110;
    x_62 = 'b000100010;
    x_63 = 'b000101011;
    x_64 = 'b000000111;
    x_65 = 'b111111011;
    x_66 = 'b111100100;
    x_67 = 'b111001111;
    x_68 = 'b111000111;
    x_69 = 'b110111101;
    x_70 = 'b111001011;
    x_71 = 'b000010111;
    x_72 = 'b111110110;
    x_73 = 'b111110001;
    x_74 = 'b111100101;
    x_75 = 'b111001100;
    x_76 = 'b111000111;
    x_77 = 'b111010000;
    x_78 = 'b000010111;
    x_79 = 'b000000011;
    x_80 = 'b111111001;
    x_81 = 'b111101101;
    x_82 = 'b111110001;
    x_83 = 'b111101001;
    x_84 = 'b111100101;
    x_85 = 'b111110101;
    x_86 = 'b111100011;
    x_87 = 'b111100011;
    x_88 = 'b000001000;
    x_89 = 'b000000111;
    x_90 = 'b111010001;
    x_91 = 'b111000111;
    x_92 = 'b111011101;
    x_93 = 'b000010100;
    x_94 = 'b111111011;
    x_95 = 'b111010100;
    x_96 = 'b111011010;
    x_97 = 'b111001101;
    x_98 = 'b111000111;
    x_99 = 'b111010000;
    x_100 = 'b111000111;
    x_101 = 'b111110100;
    x_102 = 'b000011000;
    x_103 = 'b111010101;
    x_104 = 'b000101010;
    x_105 = 'b111101011;
    x_106 = 'b000101110;
    x_107 = 'b111100100;
    x_108 = 'b000110110;
    x_109 = 'b111111110;
    x_110 = 'b000101010;
    x_111 = 'b000011011;
    x_112 = 'b000001010;
    x_113 = 'b000001000;
    x_114 = 'b111111101;
    x_115 = 'b000000101;
    x_116 = 'b000000110;
    x_117 = 'b000001100;
    x_118 = 'b000001101;
    x_119 = 'b000110000;
    x_120 = 'b000011011;
    x_121 = 'b000010000;
    x_122 = 'b000010110;
    x_123 = 'b000010001;
    x_124 = 'b000101111;
    x_125 = 'b000010110;
    x_126 = 'b000100010;
    x_127 = 'b000101011;
    x_128 = 'b000000111;
    x_129 = 'b111111011;
    x_130 = 'b111100100;
    x_131 = 'b111001111;
    x_132 = 'b111000111;
    x_133 = 'b110111101;
    x_134 = 'b111001011;
    x_135 = 'b000010111;
    x_136 = 'b111110110;
    x_137 = 'b111110001;
    x_138 = 'b111100101;
    x_139 = 'b111001100;
    x_140 = 'b111000111;
    x_141 = 'b111010000;
    x_142 = 'b000010111;
    x_143 = 'b000000011;
    x_144 = 'b111111001;
    x_145 = 'b111101101;
    x_146 = 'b111110001;
    x_147 = 'b111101001;
    x_148 = 'b111100101;
    x_149 = 'b111110101;
    x_150 = 'b111100011;
    x_151 = 'b111100011;
    x_152 = 'b000001000;
    x_153 = 'b000000111;
    x_154 = 'b111010001;
    x_155 = 'b111000111;
    x_156 = 'b111011101;
    x_157 = 'b000010100;
    x_158 = 'b111111011;
    x_159 = 'b111010100;
    x_160 = 'b111011010;
    x_161 = 'b111001101;
    x_162 = 'b111000111;
    x_163 = 'b111010000;
    x_164 = 'b111000111;
    x_165 = 'b111110100;
    x_166 = 'b000011000;
    x_167 = 'b111010101;
    x_168 = 'b000101010;
    x_169 = 'b111101011;
    x_170 = 'b000101110;
    x_171 = 'b111100100;
    x_172 = 'b000110110;
    x_173 = 'b111111110;
    x_174 = 'b000101010;
    x_175 = 'b000011011;
    x_176 = 'b000001010;
    x_177 = 'b000001000;
    x_178 = 'b111111101;
    x_179 = 'b000000101;
    x_180 = 'b000000110;
    x_181 = 'b000001100;
    x_182 = 'b000001101;
    x_183 = 'b000110000;
    x_184 = 'b000011011;
    x_185 = 'b000010000;
    x_186 = 'b000010110;
    x_187 = 'b000010001;
    x_188 = 'b000101111;
    x_189 = 'b000010110;
    x_190 = 'b000100010;
    x_191 = 'b000101011;
    x_192 = 'b000000111;
    x_193 = 'b111111011;
    x_194 = 'b111100100;
    x_195 = 'b111001111;
    x_196 = 'b111000111;
    x_197 = 'b110111101;
    x_198 = 'b111001011;
    x_199 = 'b000010111;
    x_200 = 'b111110110;
    x_201 = 'b111110001;
    x_202 = 'b111100101;
    x_203 = 'b111001100;
    x_204 = 'b111000111;
    x_205 = 'b111010000;
    x_206 = 'b000010111;
    x_207 = 'b000000011;
    x_208 = 'b111111001;
    x_209 = 'b111101101;
    x_210 = 'b111110001;
    x_211 = 'b111101001;
    x_212 = 'b111100101;
    x_213 = 'b111110101;
    x_214 = 'b111100011;
    x_215 = 'b111100011;
    x_216 = 'b000001000;
    x_217 = 'b000000111;
    x_218 = 'b111010001;
    x_219 = 'b111000111;
    x_220 = 'b111011101;
    x_221 = 'b000010100;
    x_222 = 'b111111011;
    x_223 = 'b111010100;
    x_224 = 'b111011010;
    x_225 = 'b111001101;
    x_226 = 'b111000111;
    x_227 = 'b111010000;
    x_228 = 'b111000111;
    x_229 = 'b111110100;
    x_230 = 'b000011000;
    x_231 = 'b111010101;
    x_232 = 'b000101010;
    x_233 = 'b111101011;
    x_234 = 'b000101110;
    x_235 = 'b111100100;
    x_236 = 'b000110110;
    x_237 = 'b111111110;
    x_238 = 'b000101010;
    x_239 = 'b000011011;
    x_240 = 'b000001010;
    x_241 = 'b000001000;
    x_242 = 'b111111101;
    x_243 = 'b000000101;
    x_244 = 'b000000110;
    x_245 = 'b000001100;
    x_246 = 'b000001101;
    x_247 = 'b000110000;
    x_248 = 'b000011011;
    x_249 = 'b000010000;
    x_250 = 'b000010110;
    x_251 = 'b000010001;
    x_252 = 'b000101111;
    x_253 = 'b000010110;
    x_254 = 'b000100010;
    x_255 = 'b000101011;

    h_0 = 'b000000111;
    h_1 = 'b111111011;
    h_2 = 'b111100100;
    h_3 = 'b111001111;
    h_4 = 'b111000111;
    h_5 = 'b110111101;
    h_6 = 'b111001011;
    h_7 = 'b000010111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111001010;
    x_1 = 'b111011110;
    x_2 = 'b111100001;
    x_3 = 'b111110101;
    x_4 = 'b111111001;
    x_5 = 'b111111000;
    x_6 = 'b111101000;
    x_7 = 'b111011011;
    x_8 = 'b111101100;
    x_9 = 'b111110011;
    x_10 = 'b111111011;
    x_11 = 'b000000000;
    x_12 = 'b000000011;
    x_13 = 'b111111001;
    x_14 = 'b111101100;
    x_15 = 'b111110100;
    x_16 = 'b111111000;
    x_17 = 'b000000100;
    x_18 = 'b000000101;
    x_19 = 'b000001001;
    x_20 = 'b000001100;
    x_21 = 'b111001100;
    x_22 = 'b111001001;
    x_23 = 'b111010010;
    x_24 = 'b111001000;
    x_25 = 'b111001001;
    x_26 = 'b111010110;
    x_27 = 'b111011001;
    x_28 = 'b111010110;
    x_29 = 'b111000101;
    x_30 = 'b111010011;
    x_31 = 'b111011011;
    x_32 = 'b111011101;
    x_33 = 'b111100011;
    x_34 = 'b111101010;
    x_35 = 'b111101001;
    x_36 = 'b111101000;
    x_37 = 'b111101010;
    x_38 = 'b111001010;
    x_39 = 'b111101011;
    x_40 = 'b111001110;
    x_41 = 'b000000000;
    x_42 = 'b110111110;
    x_43 = 'b000000110;
    x_44 = 'b111100001;
    x_45 = 'b111111100;
    x_46 = 'b111111101;
    x_47 = 'b111111100;
    x_48 = 'b000000011;
    x_49 = 'b000000101;
    x_50 = 'b000000110;
    x_51 = 'b000010010;
    x_52 = 'b000001011;
    x_53 = 'b000010001;
    x_54 = 'b000001011;
    x_55 = 'b000001101;
    x_56 = 'b000001101;
    x_57 = 'b000011100;
    x_58 = 'b000011100;
    x_59 = 'b000010110;
    x_60 = 'b000011101;
    x_61 = 'b000100111;
    x_62 = 'b000001011;
    x_63 = 'b000011010;
    x_64 = 'b111001010;
    x_65 = 'b111011110;
    x_66 = 'b111100001;
    x_67 = 'b111110101;
    x_68 = 'b111111001;
    x_69 = 'b111111000;
    x_70 = 'b111101000;
    x_71 = 'b111011011;
    x_72 = 'b111101100;
    x_73 = 'b111110011;
    x_74 = 'b111111011;
    x_75 = 'b000000000;
    x_76 = 'b000000011;
    x_77 = 'b111111001;
    x_78 = 'b111101100;
    x_79 = 'b111110100;
    x_80 = 'b111111000;
    x_81 = 'b000000100;
    x_82 = 'b000000101;
    x_83 = 'b000001001;
    x_84 = 'b000001100;
    x_85 = 'b111001100;
    x_86 = 'b111001001;
    x_87 = 'b111010010;
    x_88 = 'b111001000;
    x_89 = 'b111001001;
    x_90 = 'b111010110;
    x_91 = 'b111011001;
    x_92 = 'b111010110;
    x_93 = 'b111000101;
    x_94 = 'b111010011;
    x_95 = 'b111011011;
    x_96 = 'b111011101;
    x_97 = 'b111100011;
    x_98 = 'b111101010;
    x_99 = 'b111101001;
    x_100 = 'b111101000;
    x_101 = 'b111101010;
    x_102 = 'b111001010;
    x_103 = 'b111101011;
    x_104 = 'b111001110;
    x_105 = 'b000000000;
    x_106 = 'b110111110;
    x_107 = 'b000000110;
    x_108 = 'b111100001;
    x_109 = 'b111111100;
    x_110 = 'b111111101;
    x_111 = 'b111111100;
    x_112 = 'b000000011;
    x_113 = 'b000000101;
    x_114 = 'b000000110;
    x_115 = 'b000010010;
    x_116 = 'b000001011;
    x_117 = 'b000010001;
    x_118 = 'b000001011;
    x_119 = 'b000001101;
    x_120 = 'b000001101;
    x_121 = 'b000011100;
    x_122 = 'b000011100;
    x_123 = 'b000010110;
    x_124 = 'b000011101;
    x_125 = 'b000100111;
    x_126 = 'b000001011;
    x_127 = 'b000011010;
    x_128 = 'b111001010;
    x_129 = 'b111011110;
    x_130 = 'b111100001;
    x_131 = 'b111110101;
    x_132 = 'b111111001;
    x_133 = 'b111111000;
    x_134 = 'b111101000;
    x_135 = 'b111011011;
    x_136 = 'b111101100;
    x_137 = 'b111110011;
    x_138 = 'b111111011;
    x_139 = 'b000000000;
    x_140 = 'b000000011;
    x_141 = 'b111111001;
    x_142 = 'b111101100;
    x_143 = 'b111110100;
    x_144 = 'b111111000;
    x_145 = 'b000000100;
    x_146 = 'b000000101;
    x_147 = 'b000001001;
    x_148 = 'b000001100;
    x_149 = 'b111001100;
    x_150 = 'b111001001;
    x_151 = 'b111010010;
    x_152 = 'b111001000;
    x_153 = 'b111001001;
    x_154 = 'b111010110;
    x_155 = 'b111011001;
    x_156 = 'b111010110;
    x_157 = 'b111000101;
    x_158 = 'b111010011;
    x_159 = 'b111011011;
    x_160 = 'b111011101;
    x_161 = 'b111100011;
    x_162 = 'b111101010;
    x_163 = 'b111101001;
    x_164 = 'b111101000;
    x_165 = 'b111101010;
    x_166 = 'b111001010;
    x_167 = 'b111101011;
    x_168 = 'b111001110;
    x_169 = 'b000000000;
    x_170 = 'b110111110;
    x_171 = 'b000000110;
    x_172 = 'b111100001;
    x_173 = 'b111111100;
    x_174 = 'b111111101;
    x_175 = 'b111111100;
    x_176 = 'b000000011;
    x_177 = 'b000000101;
    x_178 = 'b000000110;
    x_179 = 'b000010010;
    x_180 = 'b000001011;
    x_181 = 'b000010001;
    x_182 = 'b000001011;
    x_183 = 'b000001101;
    x_184 = 'b000001101;
    x_185 = 'b000011100;
    x_186 = 'b000011100;
    x_187 = 'b000010110;
    x_188 = 'b000011101;
    x_189 = 'b000100111;
    x_190 = 'b000001011;
    x_191 = 'b000011010;
    x_192 = 'b111001010;
    x_193 = 'b111011110;
    x_194 = 'b111100001;
    x_195 = 'b111110101;
    x_196 = 'b111111001;
    x_197 = 'b111111000;
    x_198 = 'b111101000;
    x_199 = 'b111011011;
    x_200 = 'b111101100;
    x_201 = 'b111110011;
    x_202 = 'b111111011;
    x_203 = 'b000000000;
    x_204 = 'b000000011;
    x_205 = 'b111111001;
    x_206 = 'b111101100;
    x_207 = 'b111110100;
    x_208 = 'b111111000;
    x_209 = 'b000000100;
    x_210 = 'b000000101;
    x_211 = 'b000001001;
    x_212 = 'b000001100;
    x_213 = 'b111001100;
    x_214 = 'b111001001;
    x_215 = 'b111010010;
    x_216 = 'b111001000;
    x_217 = 'b111001001;
    x_218 = 'b111010110;
    x_219 = 'b111011001;
    x_220 = 'b111010110;
    x_221 = 'b111000101;
    x_222 = 'b111010011;
    x_223 = 'b111011011;
    x_224 = 'b111011101;
    x_225 = 'b111100011;
    x_226 = 'b111101010;
    x_227 = 'b111101001;
    x_228 = 'b111101000;
    x_229 = 'b111101010;
    x_230 = 'b111001010;
    x_231 = 'b111101011;
    x_232 = 'b111001110;
    x_233 = 'b000000000;
    x_234 = 'b110111110;
    x_235 = 'b000000110;
    x_236 = 'b111100001;
    x_237 = 'b111111100;
    x_238 = 'b111111101;
    x_239 = 'b111111100;
    x_240 = 'b000000011;
    x_241 = 'b000000101;
    x_242 = 'b000000110;
    x_243 = 'b000010010;
    x_244 = 'b000001011;
    x_245 = 'b000010001;
    x_246 = 'b000001011;
    x_247 = 'b000001101;
    x_248 = 'b000001101;
    x_249 = 'b000011100;
    x_250 = 'b000011100;
    x_251 = 'b000010110;
    x_252 = 'b000011101;
    x_253 = 'b000100111;
    x_254 = 'b000001011;
    x_255 = 'b000011010;

    h_0 = 'b111001010;
    h_1 = 'b111011110;
    h_2 = 'b111100001;
    h_3 = 'b111110101;
    h_4 = 'b111111001;
    h_5 = 'b111111000;
    h_6 = 'b111101000;
    h_7 = 'b111011011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111001110;
    x_1 = 'b111100100;
    x_2 = 'b111100111;
    x_3 = 'b111110101;
    x_4 = 'b111111011;
    x_5 = 'b111111110;
    x_6 = 'b111111000;
    x_7 = 'b111100010;
    x_8 = 'b111110001;
    x_9 = 'b111110100;
    x_10 = 'b111110110;
    x_11 = 'b111111111;
    x_12 = 'b000000101;
    x_13 = 'b000000101;
    x_14 = 'b111101011;
    x_15 = 'b111110011;
    x_16 = 'b111110110;
    x_17 = 'b111111100;
    x_18 = 'b111111000;
    x_19 = 'b111111111;
    x_20 = 'b000000101;
    x_21 = 'b111001001;
    x_22 = 'b111001100;
    x_23 = 'b111010111;
    x_24 = 'b111000111;
    x_25 = 'b111001000;
    x_26 = 'b111010111;
    x_27 = 'b111011111;
    x_28 = 'b111011101;
    x_29 = 'b111000111;
    x_30 = 'b111011001;
    x_31 = 'b111011111;
    x_32 = 'b111011101;
    x_33 = 'b111100100;
    x_34 = 'b111101100;
    x_35 = 'b111101011;
    x_36 = 'b111110010;
    x_37 = 'b111110000;
    x_38 = 'b111001100;
    x_39 = 'b111111100;
    x_40 = 'b111010000;
    x_41 = 'b000101001;
    x_42 = 'b110111111;
    x_43 = 'b111011111;
    x_44 = 'b111011000;
    x_45 = 'b111101011;
    x_46 = 'b111110011;
    x_47 = 'b111111001;
    x_48 = 'b000000011;
    x_49 = 'b000000001;
    x_50 = 'b111111110;
    x_51 = 'b000001000;
    x_52 = 'b000000010;
    x_53 = 'b000001011;
    x_54 = 'b000000110;
    x_55 = 'b000001100;
    x_56 = 'b000001011;
    x_57 = 'b000011001;
    x_58 = 'b000011000;
    x_59 = 'b000010101;
    x_60 = 'b000011001;
    x_61 = 'b000100011;
    x_62 = 'b000000101;
    x_63 = 'b000010111;
    x_64 = 'b111001110;
    x_65 = 'b111100100;
    x_66 = 'b111100111;
    x_67 = 'b111110101;
    x_68 = 'b111111011;
    x_69 = 'b111111110;
    x_70 = 'b111111000;
    x_71 = 'b111100010;
    x_72 = 'b111110001;
    x_73 = 'b111110100;
    x_74 = 'b111110110;
    x_75 = 'b111111111;
    x_76 = 'b000000101;
    x_77 = 'b000000101;
    x_78 = 'b111101011;
    x_79 = 'b111110011;
    x_80 = 'b111110110;
    x_81 = 'b111111100;
    x_82 = 'b111111000;
    x_83 = 'b111111111;
    x_84 = 'b000000101;
    x_85 = 'b111001001;
    x_86 = 'b111001100;
    x_87 = 'b111010111;
    x_88 = 'b111000111;
    x_89 = 'b111001000;
    x_90 = 'b111010111;
    x_91 = 'b111011111;
    x_92 = 'b111011101;
    x_93 = 'b111000111;
    x_94 = 'b111011001;
    x_95 = 'b111011111;
    x_96 = 'b111011101;
    x_97 = 'b111100100;
    x_98 = 'b111101100;
    x_99 = 'b111101011;
    x_100 = 'b111110010;
    x_101 = 'b111110000;
    x_102 = 'b111001100;
    x_103 = 'b111111100;
    x_104 = 'b111010000;
    x_105 = 'b000101001;
    x_106 = 'b110111111;
    x_107 = 'b111011111;
    x_108 = 'b111011000;
    x_109 = 'b111101011;
    x_110 = 'b111110011;
    x_111 = 'b111111001;
    x_112 = 'b000000011;
    x_113 = 'b000000001;
    x_114 = 'b111111110;
    x_115 = 'b000001000;
    x_116 = 'b000000010;
    x_117 = 'b000001011;
    x_118 = 'b000000110;
    x_119 = 'b000001100;
    x_120 = 'b000001011;
    x_121 = 'b000011001;
    x_122 = 'b000011000;
    x_123 = 'b000010101;
    x_124 = 'b000011001;
    x_125 = 'b000100011;
    x_126 = 'b000000101;
    x_127 = 'b000010111;
    x_128 = 'b111001110;
    x_129 = 'b111100100;
    x_130 = 'b111100111;
    x_131 = 'b111110101;
    x_132 = 'b111111011;
    x_133 = 'b111111110;
    x_134 = 'b111111000;
    x_135 = 'b111100010;
    x_136 = 'b111110001;
    x_137 = 'b111110100;
    x_138 = 'b111110110;
    x_139 = 'b111111111;
    x_140 = 'b000000101;
    x_141 = 'b000000101;
    x_142 = 'b111101011;
    x_143 = 'b111110011;
    x_144 = 'b111110110;
    x_145 = 'b111111100;
    x_146 = 'b111111000;
    x_147 = 'b111111111;
    x_148 = 'b000000101;
    x_149 = 'b111001001;
    x_150 = 'b111001100;
    x_151 = 'b111010111;
    x_152 = 'b111000111;
    x_153 = 'b111001000;
    x_154 = 'b111010111;
    x_155 = 'b111011111;
    x_156 = 'b111011101;
    x_157 = 'b111000111;
    x_158 = 'b111011001;
    x_159 = 'b111011111;
    x_160 = 'b111011101;
    x_161 = 'b111100100;
    x_162 = 'b111101100;
    x_163 = 'b111101011;
    x_164 = 'b111110010;
    x_165 = 'b111110000;
    x_166 = 'b111001100;
    x_167 = 'b111111100;
    x_168 = 'b111010000;
    x_169 = 'b000101001;
    x_170 = 'b110111111;
    x_171 = 'b111011111;
    x_172 = 'b111011000;
    x_173 = 'b111101011;
    x_174 = 'b111110011;
    x_175 = 'b111111001;
    x_176 = 'b000000011;
    x_177 = 'b000000001;
    x_178 = 'b111111110;
    x_179 = 'b000001000;
    x_180 = 'b000000010;
    x_181 = 'b000001011;
    x_182 = 'b000000110;
    x_183 = 'b000001100;
    x_184 = 'b000001011;
    x_185 = 'b000011001;
    x_186 = 'b000011000;
    x_187 = 'b000010101;
    x_188 = 'b000011001;
    x_189 = 'b000100011;
    x_190 = 'b000000101;
    x_191 = 'b000010111;
    x_192 = 'b111001110;
    x_193 = 'b111100100;
    x_194 = 'b111100111;
    x_195 = 'b111110101;
    x_196 = 'b111111011;
    x_197 = 'b111111110;
    x_198 = 'b111111000;
    x_199 = 'b111100010;
    x_200 = 'b111110001;
    x_201 = 'b111110100;
    x_202 = 'b111110110;
    x_203 = 'b111111111;
    x_204 = 'b000000101;
    x_205 = 'b000000101;
    x_206 = 'b111101011;
    x_207 = 'b111110011;
    x_208 = 'b111110110;
    x_209 = 'b111111100;
    x_210 = 'b111111000;
    x_211 = 'b111111111;
    x_212 = 'b000000101;
    x_213 = 'b111001001;
    x_214 = 'b111001100;
    x_215 = 'b111010111;
    x_216 = 'b111000111;
    x_217 = 'b111001000;
    x_218 = 'b111010111;
    x_219 = 'b111011111;
    x_220 = 'b111011101;
    x_221 = 'b111000111;
    x_222 = 'b111011001;
    x_223 = 'b111011111;
    x_224 = 'b111011101;
    x_225 = 'b111100100;
    x_226 = 'b111101100;
    x_227 = 'b111101011;
    x_228 = 'b111110010;
    x_229 = 'b111110000;
    x_230 = 'b111001100;
    x_231 = 'b111111100;
    x_232 = 'b111010000;
    x_233 = 'b000101001;
    x_234 = 'b110111111;
    x_235 = 'b111011111;
    x_236 = 'b111011000;
    x_237 = 'b111101011;
    x_238 = 'b111110011;
    x_239 = 'b111111001;
    x_240 = 'b000000011;
    x_241 = 'b000000001;
    x_242 = 'b111111110;
    x_243 = 'b000001000;
    x_244 = 'b000000010;
    x_245 = 'b000001011;
    x_246 = 'b000000110;
    x_247 = 'b000001100;
    x_248 = 'b000001011;
    x_249 = 'b000011001;
    x_250 = 'b000011000;
    x_251 = 'b000010101;
    x_252 = 'b000011001;
    x_253 = 'b000100011;
    x_254 = 'b000000101;
    x_255 = 'b000010111;

    h_0 = 'b111001110;
    h_1 = 'b111100100;
    h_2 = 'b111100111;
    h_3 = 'b111110101;
    h_4 = 'b111111011;
    h_5 = 'b111111110;
    h_6 = 'b111111000;
    h_7 = 'b111100010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111010101;
    x_1 = 'b111101011;
    x_2 = 'b111101011;
    x_3 = 'b111110100;
    x_4 = 'b111111001;
    x_5 = 'b111111110;
    x_6 = 'b000000000;
    x_7 = 'b111101011;
    x_8 = 'b111110111;
    x_9 = 'b111110010;
    x_10 = 'b111101111;
    x_11 = 'b111111000;
    x_12 = 'b000000010;
    x_13 = 'b000001010;
    x_14 = 'b111110000;
    x_15 = 'b111110111;
    x_16 = 'b111110100;
    x_17 = 'b111111000;
    x_18 = 'b111110000;
    x_19 = 'b111111000;
    x_20 = 'b000000110;
    x_21 = 'b111010001;
    x_22 = 'b111010001;
    x_23 = 'b111011010;
    x_24 = 'b111001111;
    x_25 = 'b111001111;
    x_26 = 'b111011011;
    x_27 = 'b111100001;
    x_28 = 'b111011101;
    x_29 = 'b111010001;
    x_30 = 'b111011010;
    x_31 = 'b111100011;
    x_32 = 'b111100011;
    x_33 = 'b111100111;
    x_34 = 'b111101110;
    x_35 = 'b111101110;
    x_36 = 'b111110010;
    x_37 = 'b111101110;
    x_38 = 'b111011011;
    x_39 = 'b111111000;
    x_40 = 'b111100000;
    x_41 = 'b000010011;
    x_42 = 'b110111100;
    x_43 = 'b000000110;
    x_44 = 'b111100100;
    x_45 = 'b111111000;
    x_46 = 'b111111111;
    x_47 = 'b000000001;
    x_48 = 'b000001001;
    x_49 = 'b000000100;
    x_50 = 'b111111111;
    x_51 = 'b000000101;
    x_52 = 'b000000000;
    x_53 = 'b000001110;
    x_54 = 'b000010000;
    x_55 = 'b000001110;
    x_56 = 'b000001101;
    x_57 = 'b000011001;
    x_58 = 'b000011011;
    x_59 = 'b000011001;
    x_60 = 'b000010111;
    x_61 = 'b000100001;
    x_62 = 'b000000101;
    x_63 = 'b000011000;
    x_64 = 'b111010101;
    x_65 = 'b111101011;
    x_66 = 'b111101011;
    x_67 = 'b111110100;
    x_68 = 'b111111001;
    x_69 = 'b111111110;
    x_70 = 'b000000000;
    x_71 = 'b111101011;
    x_72 = 'b111110111;
    x_73 = 'b111110010;
    x_74 = 'b111101111;
    x_75 = 'b111111000;
    x_76 = 'b000000010;
    x_77 = 'b000001010;
    x_78 = 'b111110000;
    x_79 = 'b111110111;
    x_80 = 'b111110100;
    x_81 = 'b111111000;
    x_82 = 'b111110000;
    x_83 = 'b111111000;
    x_84 = 'b000000110;
    x_85 = 'b111010001;
    x_86 = 'b111010001;
    x_87 = 'b111011010;
    x_88 = 'b111001111;
    x_89 = 'b111001111;
    x_90 = 'b111011011;
    x_91 = 'b111100001;
    x_92 = 'b111011101;
    x_93 = 'b111010001;
    x_94 = 'b111011010;
    x_95 = 'b111100011;
    x_96 = 'b111100011;
    x_97 = 'b111100111;
    x_98 = 'b111101110;
    x_99 = 'b111101110;
    x_100 = 'b111110010;
    x_101 = 'b111101110;
    x_102 = 'b111011011;
    x_103 = 'b111111000;
    x_104 = 'b111100000;
    x_105 = 'b000010011;
    x_106 = 'b110111100;
    x_107 = 'b000000110;
    x_108 = 'b111100100;
    x_109 = 'b111111000;
    x_110 = 'b111111111;
    x_111 = 'b000000001;
    x_112 = 'b000001001;
    x_113 = 'b000000100;
    x_114 = 'b111111111;
    x_115 = 'b000000101;
    x_116 = 'b000000000;
    x_117 = 'b000001110;
    x_118 = 'b000010000;
    x_119 = 'b000001110;
    x_120 = 'b000001101;
    x_121 = 'b000011001;
    x_122 = 'b000011011;
    x_123 = 'b000011001;
    x_124 = 'b000010111;
    x_125 = 'b000100001;
    x_126 = 'b000000101;
    x_127 = 'b000011000;
    x_128 = 'b111010101;
    x_129 = 'b111101011;
    x_130 = 'b111101011;
    x_131 = 'b111110100;
    x_132 = 'b111111001;
    x_133 = 'b111111110;
    x_134 = 'b000000000;
    x_135 = 'b111101011;
    x_136 = 'b111110111;
    x_137 = 'b111110010;
    x_138 = 'b111101111;
    x_139 = 'b111111000;
    x_140 = 'b000000010;
    x_141 = 'b000001010;
    x_142 = 'b111110000;
    x_143 = 'b111110111;
    x_144 = 'b111110100;
    x_145 = 'b111111000;
    x_146 = 'b111110000;
    x_147 = 'b111111000;
    x_148 = 'b000000110;
    x_149 = 'b111010001;
    x_150 = 'b111010001;
    x_151 = 'b111011010;
    x_152 = 'b111001111;
    x_153 = 'b111001111;
    x_154 = 'b111011011;
    x_155 = 'b111100001;
    x_156 = 'b111011101;
    x_157 = 'b111010001;
    x_158 = 'b111011010;
    x_159 = 'b111100011;
    x_160 = 'b111100011;
    x_161 = 'b111100111;
    x_162 = 'b111101110;
    x_163 = 'b111101110;
    x_164 = 'b111110010;
    x_165 = 'b111101110;
    x_166 = 'b111011011;
    x_167 = 'b111111000;
    x_168 = 'b111100000;
    x_169 = 'b000010011;
    x_170 = 'b110111100;
    x_171 = 'b000000110;
    x_172 = 'b111100100;
    x_173 = 'b111111000;
    x_174 = 'b111111111;
    x_175 = 'b000000001;
    x_176 = 'b000001001;
    x_177 = 'b000000100;
    x_178 = 'b111111111;
    x_179 = 'b000000101;
    x_180 = 'b000000000;
    x_181 = 'b000001110;
    x_182 = 'b000010000;
    x_183 = 'b000001110;
    x_184 = 'b000001101;
    x_185 = 'b000011001;
    x_186 = 'b000011011;
    x_187 = 'b000011001;
    x_188 = 'b000010111;
    x_189 = 'b000100001;
    x_190 = 'b000000101;
    x_191 = 'b000011000;
    x_192 = 'b111010101;
    x_193 = 'b111101011;
    x_194 = 'b111101011;
    x_195 = 'b111110100;
    x_196 = 'b111111001;
    x_197 = 'b111111110;
    x_198 = 'b000000000;
    x_199 = 'b111101011;
    x_200 = 'b111110111;
    x_201 = 'b111110010;
    x_202 = 'b111101111;
    x_203 = 'b111111000;
    x_204 = 'b000000010;
    x_205 = 'b000001010;
    x_206 = 'b111110000;
    x_207 = 'b111110111;
    x_208 = 'b111110100;
    x_209 = 'b111111000;
    x_210 = 'b111110000;
    x_211 = 'b111111000;
    x_212 = 'b000000110;
    x_213 = 'b111010001;
    x_214 = 'b111010001;
    x_215 = 'b111011010;
    x_216 = 'b111001111;
    x_217 = 'b111001111;
    x_218 = 'b111011011;
    x_219 = 'b111100001;
    x_220 = 'b111011101;
    x_221 = 'b111010001;
    x_222 = 'b111011010;
    x_223 = 'b111100011;
    x_224 = 'b111100011;
    x_225 = 'b111100111;
    x_226 = 'b111101110;
    x_227 = 'b111101110;
    x_228 = 'b111110010;
    x_229 = 'b111101110;
    x_230 = 'b111011011;
    x_231 = 'b111111000;
    x_232 = 'b111100000;
    x_233 = 'b000010011;
    x_234 = 'b110111100;
    x_235 = 'b000000110;
    x_236 = 'b111100100;
    x_237 = 'b111111000;
    x_238 = 'b111111111;
    x_239 = 'b000000001;
    x_240 = 'b000001001;
    x_241 = 'b000000100;
    x_242 = 'b111111111;
    x_243 = 'b000000101;
    x_244 = 'b000000000;
    x_245 = 'b000001110;
    x_246 = 'b000010000;
    x_247 = 'b000001110;
    x_248 = 'b000001101;
    x_249 = 'b000011001;
    x_250 = 'b000011011;
    x_251 = 'b000011001;
    x_252 = 'b000010111;
    x_253 = 'b000100001;
    x_254 = 'b000000101;
    x_255 = 'b000011000;

    h_0 = 'b111010101;
    h_1 = 'b111101011;
    h_2 = 'b111101011;
    h_3 = 'b111110100;
    h_4 = 'b111111001;
    h_5 = 'b111111110;
    h_6 = 'b000000000;
    h_7 = 'b111101011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111100010;
    x_1 = 'b111110010;
    x_2 = 'b111101111;
    x_3 = 'b111110101;
    x_4 = 'b111111000;
    x_5 = 'b111111010;
    x_6 = 'b111111000;
    x_7 = 'b111110101;
    x_8 = 'b111111011;
    x_9 = 'b111110101;
    x_10 = 'b111110100;
    x_11 = 'b111110100;
    x_12 = 'b111111000;
    x_13 = 'b111110011;
    x_14 = 'b111111001;
    x_15 = 'b111111010;
    x_16 = 'b111111000;
    x_17 = 'b111111000;
    x_18 = 'b111101011;
    x_19 = 'b111101111;
    x_20 = 'b111111000;
    x_21 = 'b111010001;
    x_22 = 'b111010000;
    x_23 = 'b111011001;
    x_24 = 'b111010000;
    x_25 = 'b111010001;
    x_26 = 'b111011100;
    x_27 = 'b111100001;
    x_28 = 'b111011101;
    x_29 = 'b111010100;
    x_30 = 'b111011111;
    x_31 = 'b111100010;
    x_32 = 'b111100100;
    x_33 = 'b111100111;
    x_34 = 'b111101111;
    x_35 = 'b111110000;
    x_36 = 'b111101100;
    x_37 = 'b111101101;
    x_38 = 'b111011000;
    x_39 = 'b111100101;
    x_40 = 'b111010111;
    x_41 = 'b111010000;
    x_42 = 'b111000100;
    x_43 = 'b111100111;
    x_44 = 'b111100001;
    x_45 = 'b111101100;
    x_46 = 'b111110110;
    x_47 = 'b111110110;
    x_48 = 'b111111101;
    x_49 = 'b111111011;
    x_50 = 'b111111100;
    x_51 = 'b111111110;
    x_52 = 'b111111001;
    x_53 = 'b000000010;
    x_54 = 'b000000011;
    x_55 = 'b111111001;
    x_56 = 'b111111011;
    x_57 = 'b000001110;
    x_58 = 'b000001110;
    x_59 = 'b000001101;
    x_60 = 'b000001100;
    x_61 = 'b000010111;
    x_62 = 'b111111110;
    x_63 = 'b000001100;
    x_64 = 'b111100010;
    x_65 = 'b111110010;
    x_66 = 'b111101111;
    x_67 = 'b111110101;
    x_68 = 'b111111000;
    x_69 = 'b111111010;
    x_70 = 'b111111000;
    x_71 = 'b111110101;
    x_72 = 'b111111011;
    x_73 = 'b111110101;
    x_74 = 'b111110100;
    x_75 = 'b111110100;
    x_76 = 'b111111000;
    x_77 = 'b111110011;
    x_78 = 'b111111001;
    x_79 = 'b111111010;
    x_80 = 'b111111000;
    x_81 = 'b111111000;
    x_82 = 'b111101011;
    x_83 = 'b111101111;
    x_84 = 'b111111000;
    x_85 = 'b111010001;
    x_86 = 'b111010000;
    x_87 = 'b111011001;
    x_88 = 'b111010000;
    x_89 = 'b111010001;
    x_90 = 'b111011100;
    x_91 = 'b111100001;
    x_92 = 'b111011101;
    x_93 = 'b111010100;
    x_94 = 'b111011111;
    x_95 = 'b111100010;
    x_96 = 'b111100100;
    x_97 = 'b111100111;
    x_98 = 'b111101111;
    x_99 = 'b111110000;
    x_100 = 'b111101100;
    x_101 = 'b111101101;
    x_102 = 'b111011000;
    x_103 = 'b111100101;
    x_104 = 'b111010111;
    x_105 = 'b111010000;
    x_106 = 'b111000100;
    x_107 = 'b111100111;
    x_108 = 'b111100001;
    x_109 = 'b111101100;
    x_110 = 'b111110110;
    x_111 = 'b111110110;
    x_112 = 'b111111101;
    x_113 = 'b111111011;
    x_114 = 'b111111100;
    x_115 = 'b111111110;
    x_116 = 'b111111001;
    x_117 = 'b000000010;
    x_118 = 'b000000011;
    x_119 = 'b111111001;
    x_120 = 'b111111011;
    x_121 = 'b000001110;
    x_122 = 'b000001110;
    x_123 = 'b000001101;
    x_124 = 'b000001100;
    x_125 = 'b000010111;
    x_126 = 'b111111110;
    x_127 = 'b000001100;
    x_128 = 'b111100010;
    x_129 = 'b111110010;
    x_130 = 'b111101111;
    x_131 = 'b111110101;
    x_132 = 'b111111000;
    x_133 = 'b111111010;
    x_134 = 'b111111000;
    x_135 = 'b111110101;
    x_136 = 'b111111011;
    x_137 = 'b111110101;
    x_138 = 'b111110100;
    x_139 = 'b111110100;
    x_140 = 'b111111000;
    x_141 = 'b111110011;
    x_142 = 'b111111001;
    x_143 = 'b111111010;
    x_144 = 'b111111000;
    x_145 = 'b111111000;
    x_146 = 'b111101011;
    x_147 = 'b111101111;
    x_148 = 'b111111000;
    x_149 = 'b111010001;
    x_150 = 'b111010000;
    x_151 = 'b111011001;
    x_152 = 'b111010000;
    x_153 = 'b111010001;
    x_154 = 'b111011100;
    x_155 = 'b111100001;
    x_156 = 'b111011101;
    x_157 = 'b111010100;
    x_158 = 'b111011111;
    x_159 = 'b111100010;
    x_160 = 'b111100100;
    x_161 = 'b111100111;
    x_162 = 'b111101111;
    x_163 = 'b111110000;
    x_164 = 'b111101100;
    x_165 = 'b111101101;
    x_166 = 'b111011000;
    x_167 = 'b111100101;
    x_168 = 'b111010111;
    x_169 = 'b111010000;
    x_170 = 'b111000100;
    x_171 = 'b111100111;
    x_172 = 'b111100001;
    x_173 = 'b111101100;
    x_174 = 'b111110110;
    x_175 = 'b111110110;
    x_176 = 'b111111101;
    x_177 = 'b111111011;
    x_178 = 'b111111100;
    x_179 = 'b111111110;
    x_180 = 'b111111001;
    x_181 = 'b000000010;
    x_182 = 'b000000011;
    x_183 = 'b111111001;
    x_184 = 'b111111011;
    x_185 = 'b000001110;
    x_186 = 'b000001110;
    x_187 = 'b000001101;
    x_188 = 'b000001100;
    x_189 = 'b000010111;
    x_190 = 'b111111110;
    x_191 = 'b000001100;
    x_192 = 'b111100010;
    x_193 = 'b111110010;
    x_194 = 'b111101111;
    x_195 = 'b111110101;
    x_196 = 'b111111000;
    x_197 = 'b111111010;
    x_198 = 'b111111000;
    x_199 = 'b111110101;
    x_200 = 'b111111011;
    x_201 = 'b111110101;
    x_202 = 'b111110100;
    x_203 = 'b111110100;
    x_204 = 'b111111000;
    x_205 = 'b111110011;
    x_206 = 'b111111001;
    x_207 = 'b111111010;
    x_208 = 'b111111000;
    x_209 = 'b111111000;
    x_210 = 'b111101011;
    x_211 = 'b111101111;
    x_212 = 'b111111000;
    x_213 = 'b111010001;
    x_214 = 'b111010000;
    x_215 = 'b111011001;
    x_216 = 'b111010000;
    x_217 = 'b111010001;
    x_218 = 'b111011100;
    x_219 = 'b111100001;
    x_220 = 'b111011101;
    x_221 = 'b111010100;
    x_222 = 'b111011111;
    x_223 = 'b111100010;
    x_224 = 'b111100100;
    x_225 = 'b111100111;
    x_226 = 'b111101111;
    x_227 = 'b111110000;
    x_228 = 'b111101100;
    x_229 = 'b111101101;
    x_230 = 'b111011000;
    x_231 = 'b111100101;
    x_232 = 'b111010111;
    x_233 = 'b111010000;
    x_234 = 'b111000100;
    x_235 = 'b111100111;
    x_236 = 'b111100001;
    x_237 = 'b111101100;
    x_238 = 'b111110110;
    x_239 = 'b111110110;
    x_240 = 'b111111101;
    x_241 = 'b111111011;
    x_242 = 'b111111100;
    x_243 = 'b111111110;
    x_244 = 'b111111001;
    x_245 = 'b000000010;
    x_246 = 'b000000011;
    x_247 = 'b111111001;
    x_248 = 'b111111011;
    x_249 = 'b000001110;
    x_250 = 'b000001110;
    x_251 = 'b000001101;
    x_252 = 'b000001100;
    x_253 = 'b000010111;
    x_254 = 'b111111110;
    x_255 = 'b000001100;

    h_0 = 'b111100010;
    h_1 = 'b111110010;
    h_2 = 'b111101111;
    h_3 = 'b111110101;
    h_4 = 'b111111000;
    h_5 = 'b111111010;
    h_6 = 'b111111000;
    h_7 = 'b111110101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111011111;
    x_1 = 'b111101111;
    x_2 = 'b111101110;
    x_3 = 'b111110101;
    x_4 = 'b111110111;
    x_5 = 'b111110111;
    x_6 = 'b111101110;
    x_7 = 'b111101100;
    x_8 = 'b111110111;
    x_9 = 'b111110111;
    x_10 = 'b111111001;
    x_11 = 'b111111100;
    x_12 = 'b111110110;
    x_13 = 'b111101111;
    x_14 = 'b111101010;
    x_15 = 'b111110011;
    x_16 = 'b111111001;
    x_17 = 'b111111100;
    x_18 = 'b111110101;
    x_19 = 'b111110110;
    x_20 = 'b111111100;
    x_21 = 'b111001011;
    x_22 = 'b111001001;
    x_23 = 'b111010001;
    x_24 = 'b111001001;
    x_25 = 'b111001011;
    x_26 = 'b111011001;
    x_27 = 'b111011011;
    x_28 = 'b111010111;
    x_29 = 'b111001110;
    x_30 = 'b111100110;
    x_31 = 'b111100100;
    x_32 = 'b111100011;
    x_33 = 'b111101000;
    x_34 = 'b111101111;
    x_35 = 'b111101110;
    x_36 = 'b111101000;
    x_37 = 'b111110000;
    x_38 = 'b111011010;
    x_39 = 'b111101110;
    x_40 = 'b111100101;
    x_41 = 'b000010001;
    x_42 = 'b111000011;
    x_43 = 'b111101000;
    x_44 = 'b111100010;
    x_45 = 'b111110011;
    x_46 = 'b111101101;
    x_47 = 'b111110001;
    x_48 = 'b000000000;
    x_49 = 'b000000001;
    x_50 = 'b000000110;
    x_51 = 'b000001101;
    x_52 = 'b000001010;
    x_53 = 'b000001110;
    x_54 = 'b000001110;
    x_55 = 'b111110100;
    x_56 = 'b111111010;
    x_57 = 'b000010001;
    x_58 = 'b000010111;
    x_59 = 'b000010101;
    x_60 = 'b000000000;
    x_61 = 'b000001100;
    x_62 = 'b111111001;
    x_63 = 'b111111110;
    x_64 = 'b111011111;
    x_65 = 'b111101111;
    x_66 = 'b111101110;
    x_67 = 'b111110101;
    x_68 = 'b111110111;
    x_69 = 'b111110111;
    x_70 = 'b111101110;
    x_71 = 'b111101100;
    x_72 = 'b111110111;
    x_73 = 'b111110111;
    x_74 = 'b111111001;
    x_75 = 'b111111100;
    x_76 = 'b111110110;
    x_77 = 'b111101111;
    x_78 = 'b111101010;
    x_79 = 'b111110011;
    x_80 = 'b111111001;
    x_81 = 'b111111100;
    x_82 = 'b111110101;
    x_83 = 'b111110110;
    x_84 = 'b111111100;
    x_85 = 'b111001011;
    x_86 = 'b111001001;
    x_87 = 'b111010001;
    x_88 = 'b111001001;
    x_89 = 'b111001011;
    x_90 = 'b111011001;
    x_91 = 'b111011011;
    x_92 = 'b111010111;
    x_93 = 'b111001110;
    x_94 = 'b111100110;
    x_95 = 'b111100100;
    x_96 = 'b111100011;
    x_97 = 'b111101000;
    x_98 = 'b111101111;
    x_99 = 'b111101110;
    x_100 = 'b111101000;
    x_101 = 'b111110000;
    x_102 = 'b111011010;
    x_103 = 'b111101110;
    x_104 = 'b111100101;
    x_105 = 'b000010001;
    x_106 = 'b111000011;
    x_107 = 'b111101000;
    x_108 = 'b111100010;
    x_109 = 'b111110011;
    x_110 = 'b111101101;
    x_111 = 'b111110001;
    x_112 = 'b000000000;
    x_113 = 'b000000001;
    x_114 = 'b000000110;
    x_115 = 'b000001101;
    x_116 = 'b000001010;
    x_117 = 'b000001110;
    x_118 = 'b000001110;
    x_119 = 'b111110100;
    x_120 = 'b111111010;
    x_121 = 'b000010001;
    x_122 = 'b000010111;
    x_123 = 'b000010101;
    x_124 = 'b000000000;
    x_125 = 'b000001100;
    x_126 = 'b111111001;
    x_127 = 'b111111110;
    x_128 = 'b111011111;
    x_129 = 'b111101111;
    x_130 = 'b111101110;
    x_131 = 'b111110101;
    x_132 = 'b111110111;
    x_133 = 'b111110111;
    x_134 = 'b111101110;
    x_135 = 'b111101100;
    x_136 = 'b111110111;
    x_137 = 'b111110111;
    x_138 = 'b111111001;
    x_139 = 'b111111100;
    x_140 = 'b111110110;
    x_141 = 'b111101111;
    x_142 = 'b111101010;
    x_143 = 'b111110011;
    x_144 = 'b111111001;
    x_145 = 'b111111100;
    x_146 = 'b111110101;
    x_147 = 'b111110110;
    x_148 = 'b111111100;
    x_149 = 'b111001011;
    x_150 = 'b111001001;
    x_151 = 'b111010001;
    x_152 = 'b111001001;
    x_153 = 'b111001011;
    x_154 = 'b111011001;
    x_155 = 'b111011011;
    x_156 = 'b111010111;
    x_157 = 'b111001110;
    x_158 = 'b111100110;
    x_159 = 'b111100100;
    x_160 = 'b111100011;
    x_161 = 'b111101000;
    x_162 = 'b111101111;
    x_163 = 'b111101110;
    x_164 = 'b111101000;
    x_165 = 'b111110000;
    x_166 = 'b111011010;
    x_167 = 'b111101110;
    x_168 = 'b111100101;
    x_169 = 'b000010001;
    x_170 = 'b111000011;
    x_171 = 'b111101000;
    x_172 = 'b111100010;
    x_173 = 'b111110011;
    x_174 = 'b111101101;
    x_175 = 'b111110001;
    x_176 = 'b000000000;
    x_177 = 'b000000001;
    x_178 = 'b000000110;
    x_179 = 'b000001101;
    x_180 = 'b000001010;
    x_181 = 'b000001110;
    x_182 = 'b000001110;
    x_183 = 'b111110100;
    x_184 = 'b111111010;
    x_185 = 'b000010001;
    x_186 = 'b000010111;
    x_187 = 'b000010101;
    x_188 = 'b000000000;
    x_189 = 'b000001100;
    x_190 = 'b111111001;
    x_191 = 'b111111110;
    x_192 = 'b111011111;
    x_193 = 'b111101111;
    x_194 = 'b111101110;
    x_195 = 'b111110101;
    x_196 = 'b111110111;
    x_197 = 'b111110111;
    x_198 = 'b111101110;
    x_199 = 'b111101100;
    x_200 = 'b111110111;
    x_201 = 'b111110111;
    x_202 = 'b111111001;
    x_203 = 'b111111100;
    x_204 = 'b111110110;
    x_205 = 'b111101111;
    x_206 = 'b111101010;
    x_207 = 'b111110011;
    x_208 = 'b111111001;
    x_209 = 'b111111100;
    x_210 = 'b111110101;
    x_211 = 'b111110110;
    x_212 = 'b111111100;
    x_213 = 'b111001011;
    x_214 = 'b111001001;
    x_215 = 'b111010001;
    x_216 = 'b111001001;
    x_217 = 'b111001011;
    x_218 = 'b111011001;
    x_219 = 'b111011011;
    x_220 = 'b111010111;
    x_221 = 'b111001110;
    x_222 = 'b111100110;
    x_223 = 'b111100100;
    x_224 = 'b111100011;
    x_225 = 'b111101000;
    x_226 = 'b111101111;
    x_227 = 'b111101110;
    x_228 = 'b111101000;
    x_229 = 'b111110000;
    x_230 = 'b111011010;
    x_231 = 'b111101110;
    x_232 = 'b111100101;
    x_233 = 'b000010001;
    x_234 = 'b111000011;
    x_235 = 'b111101000;
    x_236 = 'b111100010;
    x_237 = 'b111110011;
    x_238 = 'b111101101;
    x_239 = 'b111110001;
    x_240 = 'b000000000;
    x_241 = 'b000000001;
    x_242 = 'b000000110;
    x_243 = 'b000001101;
    x_244 = 'b000001010;
    x_245 = 'b000001110;
    x_246 = 'b000001110;
    x_247 = 'b111110100;
    x_248 = 'b111111010;
    x_249 = 'b000010001;
    x_250 = 'b000010111;
    x_251 = 'b000010101;
    x_252 = 'b000000000;
    x_253 = 'b000001100;
    x_254 = 'b111111001;
    x_255 = 'b111111110;

    h_0 = 'b111011111;
    h_1 = 'b111101111;
    h_2 = 'b111101110;
    h_3 = 'b111110101;
    h_4 = 'b111110111;
    h_5 = 'b111110111;
    h_6 = 'b111101110;
    h_7 = 'b111101100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111100000;
    x_1 = 'b111110000;
    x_2 = 'b111110100;
    x_3 = 'b111111110;
    x_4 = 'b000000010;
    x_5 = 'b000000100;
    x_6 = 'b111111101;
    x_7 = 'b111110010;
    x_8 = 'b111111100;
    x_9 = 'b111111110;
    x_10 = 'b000000000;
    x_11 = 'b000000100;
    x_12 = 'b000001000;
    x_13 = 'b000000101;
    x_14 = 'b111101000;
    x_15 = 'b111110110;
    x_16 = 'b111111101;
    x_17 = 'b000000100;
    x_18 = 'b000000101;
    x_19 = 'b000000110;
    x_20 = 'b000000110;
    x_21 = 'b111001110;
    x_22 = 'b111001111;
    x_23 = 'b111010110;
    x_24 = 'b111001011;
    x_25 = 'b111001100;
    x_26 = 'b111011100;
    x_27 = 'b111011111;
    x_28 = 'b111011010;
    x_29 = 'b111010101;
    x_30 = 'b111011111;
    x_31 = 'b111100011;
    x_32 = 'b111100100;
    x_33 = 'b111101000;
    x_34 = 'b111110010;
    x_35 = 'b111101110;
    x_36 = 'b111101011;
    x_37 = 'b111110011;
    x_38 = 'b111011000;
    x_39 = 'b111101101;
    x_40 = 'b111010000;
    x_41 = 'b111100110;
    x_42 = 'b110111101;
    x_43 = 'b000000100;
    x_44 = 'b111011011;
    x_45 = 'b111100111;
    x_46 = 'b111100110;
    x_47 = 'b111101000;
    x_48 = 'b111110111;
    x_49 = 'b111111000;
    x_50 = 'b000000000;
    x_51 = 'b000001100;
    x_52 = 'b000001000;
    x_53 = 'b000001001;
    x_54 = 'b000000110;
    x_55 = 'b111101110;
    x_56 = 'b111110011;
    x_57 = 'b000001011;
    x_58 = 'b000010000;
    x_59 = 'b000001101;
    x_60 = 'b111110111;
    x_61 = 'b000000101;
    x_62 = 'b111110101;
    x_63 = 'b111110010;
    x_64 = 'b111100000;
    x_65 = 'b111110000;
    x_66 = 'b111110100;
    x_67 = 'b111111110;
    x_68 = 'b000000010;
    x_69 = 'b000000100;
    x_70 = 'b111111101;
    x_71 = 'b111110010;
    x_72 = 'b111111100;
    x_73 = 'b111111110;
    x_74 = 'b000000000;
    x_75 = 'b000000100;
    x_76 = 'b000001000;
    x_77 = 'b000000101;
    x_78 = 'b111101000;
    x_79 = 'b111110110;
    x_80 = 'b111111101;
    x_81 = 'b000000100;
    x_82 = 'b000000101;
    x_83 = 'b000000110;
    x_84 = 'b000000110;
    x_85 = 'b111001110;
    x_86 = 'b111001111;
    x_87 = 'b111010110;
    x_88 = 'b111001011;
    x_89 = 'b111001100;
    x_90 = 'b111011100;
    x_91 = 'b111011111;
    x_92 = 'b111011010;
    x_93 = 'b111010101;
    x_94 = 'b111011111;
    x_95 = 'b111100011;
    x_96 = 'b111100100;
    x_97 = 'b111101000;
    x_98 = 'b111110010;
    x_99 = 'b111101110;
    x_100 = 'b111101011;
    x_101 = 'b111110011;
    x_102 = 'b111011000;
    x_103 = 'b111101101;
    x_104 = 'b111010000;
    x_105 = 'b111100110;
    x_106 = 'b110111101;
    x_107 = 'b000000100;
    x_108 = 'b111011011;
    x_109 = 'b111100111;
    x_110 = 'b111100110;
    x_111 = 'b111101000;
    x_112 = 'b111110111;
    x_113 = 'b111111000;
    x_114 = 'b000000000;
    x_115 = 'b000001100;
    x_116 = 'b000001000;
    x_117 = 'b000001001;
    x_118 = 'b000000110;
    x_119 = 'b111101110;
    x_120 = 'b111110011;
    x_121 = 'b000001011;
    x_122 = 'b000010000;
    x_123 = 'b000001101;
    x_124 = 'b111110111;
    x_125 = 'b000000101;
    x_126 = 'b111110101;
    x_127 = 'b111110010;
    x_128 = 'b111100000;
    x_129 = 'b111110000;
    x_130 = 'b111110100;
    x_131 = 'b111111110;
    x_132 = 'b000000010;
    x_133 = 'b000000100;
    x_134 = 'b111111101;
    x_135 = 'b111110010;
    x_136 = 'b111111100;
    x_137 = 'b111111110;
    x_138 = 'b000000000;
    x_139 = 'b000000100;
    x_140 = 'b000001000;
    x_141 = 'b000000101;
    x_142 = 'b111101000;
    x_143 = 'b111110110;
    x_144 = 'b111111101;
    x_145 = 'b000000100;
    x_146 = 'b000000101;
    x_147 = 'b000000110;
    x_148 = 'b000000110;
    x_149 = 'b111001110;
    x_150 = 'b111001111;
    x_151 = 'b111010110;
    x_152 = 'b111001011;
    x_153 = 'b111001100;
    x_154 = 'b111011100;
    x_155 = 'b111011111;
    x_156 = 'b111011010;
    x_157 = 'b111010101;
    x_158 = 'b111011111;
    x_159 = 'b111100011;
    x_160 = 'b111100100;
    x_161 = 'b111101000;
    x_162 = 'b111110010;
    x_163 = 'b111101110;
    x_164 = 'b111101011;
    x_165 = 'b111110011;
    x_166 = 'b111011000;
    x_167 = 'b111101101;
    x_168 = 'b111010000;
    x_169 = 'b111100110;
    x_170 = 'b110111101;
    x_171 = 'b000000100;
    x_172 = 'b111011011;
    x_173 = 'b111100111;
    x_174 = 'b111100110;
    x_175 = 'b111101000;
    x_176 = 'b111110111;
    x_177 = 'b111111000;
    x_178 = 'b000000000;
    x_179 = 'b000001100;
    x_180 = 'b000001000;
    x_181 = 'b000001001;
    x_182 = 'b000000110;
    x_183 = 'b111101110;
    x_184 = 'b111110011;
    x_185 = 'b000001011;
    x_186 = 'b000010000;
    x_187 = 'b000001101;
    x_188 = 'b111110111;
    x_189 = 'b000000101;
    x_190 = 'b111110101;
    x_191 = 'b111110010;
    x_192 = 'b111100000;
    x_193 = 'b111110000;
    x_194 = 'b111110100;
    x_195 = 'b111111110;
    x_196 = 'b000000010;
    x_197 = 'b000000100;
    x_198 = 'b111111101;
    x_199 = 'b111110010;
    x_200 = 'b111111100;
    x_201 = 'b111111110;
    x_202 = 'b000000000;
    x_203 = 'b000000100;
    x_204 = 'b000001000;
    x_205 = 'b000000101;
    x_206 = 'b111101000;
    x_207 = 'b111110110;
    x_208 = 'b111111101;
    x_209 = 'b000000100;
    x_210 = 'b000000101;
    x_211 = 'b000000110;
    x_212 = 'b000000110;
    x_213 = 'b111001110;
    x_214 = 'b111001111;
    x_215 = 'b111010110;
    x_216 = 'b111001011;
    x_217 = 'b111001100;
    x_218 = 'b111011100;
    x_219 = 'b111011111;
    x_220 = 'b111011010;
    x_221 = 'b111010101;
    x_222 = 'b111011111;
    x_223 = 'b111100011;
    x_224 = 'b111100100;
    x_225 = 'b111101000;
    x_226 = 'b111110010;
    x_227 = 'b111101110;
    x_228 = 'b111101011;
    x_229 = 'b111110011;
    x_230 = 'b111011000;
    x_231 = 'b111101101;
    x_232 = 'b111010000;
    x_233 = 'b111100110;
    x_234 = 'b110111101;
    x_235 = 'b000000100;
    x_236 = 'b111011011;
    x_237 = 'b111100111;
    x_238 = 'b111100110;
    x_239 = 'b111101000;
    x_240 = 'b111110111;
    x_241 = 'b111111000;
    x_242 = 'b000000000;
    x_243 = 'b000001100;
    x_244 = 'b000001000;
    x_245 = 'b000001001;
    x_246 = 'b000000110;
    x_247 = 'b111101110;
    x_248 = 'b111110011;
    x_249 = 'b000001011;
    x_250 = 'b000010000;
    x_251 = 'b000001101;
    x_252 = 'b111110111;
    x_253 = 'b000000101;
    x_254 = 'b111110101;
    x_255 = 'b111110010;

    h_0 = 'b111100000;
    h_1 = 'b111110000;
    h_2 = 'b111110100;
    h_3 = 'b111111110;
    h_4 = 'b000000010;
    h_5 = 'b000000100;
    h_6 = 'b111111101;
    h_7 = 'b111110010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111010001;
    x_1 = 'b111100100;
    x_2 = 'b111100111;
    x_3 = 'b111110111;
    x_4 = 'b111111011;
    x_5 = 'b111111100;
    x_6 = 'b111110010;
    x_7 = 'b111011111;
    x_8 = 'b111101110;
    x_9 = 'b111101111;
    x_10 = 'b111110100;
    x_11 = 'b111111111;
    x_12 = 'b000000101;
    x_13 = 'b111111001;
    x_14 = 'b111011111;
    x_15 = 'b111101000;
    x_16 = 'b111110001;
    x_17 = 'b111111100;
    x_18 = 'b000000010;
    x_19 = 'b000000110;
    x_20 = 'b000000010;
    x_21 = 'b111001010;
    x_22 = 'b111001100;
    x_23 = 'b111010110;
    x_24 = 'b111001000;
    x_25 = 'b111001001;
    x_26 = 'b111010111;
    x_27 = 'b111011111;
    x_28 = 'b111011011;
    x_29 = 'b111001110;
    x_30 = 'b111011110;
    x_31 = 'b111100000;
    x_32 = 'b111011110;
    x_33 = 'b111100011;
    x_34 = 'b111101111;
    x_35 = 'b111101110;
    x_36 = 'b111101110;
    x_37 = 'b111110010;
    x_38 = 'b111001100;
    x_39 = 'b111110011;
    x_40 = 'b111000101;
    x_41 = 'b111100111;
    x_42 = 'b111000010;
    x_43 = 'b111111011;
    x_44 = 'b111011100;
    x_45 = 'b111110001;
    x_46 = 'b111101101;
    x_47 = 'b111101101;
    x_48 = 'b111111000;
    x_49 = 'b111111010;
    x_50 = 'b000000110;
    x_51 = 'b000010101;
    x_52 = 'b000010001;
    x_53 = 'b000010011;
    x_54 = 'b000001111;
    x_55 = 'b111111001;
    x_56 = 'b111111100;
    x_57 = 'b000010110;
    x_58 = 'b000011000;
    x_59 = 'b000010100;
    x_60 = 'b111111000;
    x_61 = 'b000000101;
    x_62 = 'b111110111;
    x_63 = 'b111110001;
    x_64 = 'b111010001;
    x_65 = 'b111100100;
    x_66 = 'b111100111;
    x_67 = 'b111110111;
    x_68 = 'b111111011;
    x_69 = 'b111111100;
    x_70 = 'b111110010;
    x_71 = 'b111011111;
    x_72 = 'b111101110;
    x_73 = 'b111101111;
    x_74 = 'b111110100;
    x_75 = 'b111111111;
    x_76 = 'b000000101;
    x_77 = 'b111111001;
    x_78 = 'b111011111;
    x_79 = 'b111101000;
    x_80 = 'b111110001;
    x_81 = 'b111111100;
    x_82 = 'b000000010;
    x_83 = 'b000000110;
    x_84 = 'b000000010;
    x_85 = 'b111001010;
    x_86 = 'b111001100;
    x_87 = 'b111010110;
    x_88 = 'b111001000;
    x_89 = 'b111001001;
    x_90 = 'b111010111;
    x_91 = 'b111011111;
    x_92 = 'b111011011;
    x_93 = 'b111001110;
    x_94 = 'b111011110;
    x_95 = 'b111100000;
    x_96 = 'b111011110;
    x_97 = 'b111100011;
    x_98 = 'b111101111;
    x_99 = 'b111101110;
    x_100 = 'b111101110;
    x_101 = 'b111110010;
    x_102 = 'b111001100;
    x_103 = 'b111110011;
    x_104 = 'b111000101;
    x_105 = 'b111100111;
    x_106 = 'b111000010;
    x_107 = 'b111111011;
    x_108 = 'b111011100;
    x_109 = 'b111110001;
    x_110 = 'b111101101;
    x_111 = 'b111101101;
    x_112 = 'b111111000;
    x_113 = 'b111111010;
    x_114 = 'b000000110;
    x_115 = 'b000010101;
    x_116 = 'b000010001;
    x_117 = 'b000010011;
    x_118 = 'b000001111;
    x_119 = 'b111111001;
    x_120 = 'b111111100;
    x_121 = 'b000010110;
    x_122 = 'b000011000;
    x_123 = 'b000010100;
    x_124 = 'b111111000;
    x_125 = 'b000000101;
    x_126 = 'b111110111;
    x_127 = 'b111110001;
    x_128 = 'b111010001;
    x_129 = 'b111100100;
    x_130 = 'b111100111;
    x_131 = 'b111110111;
    x_132 = 'b111111011;
    x_133 = 'b111111100;
    x_134 = 'b111110010;
    x_135 = 'b111011111;
    x_136 = 'b111101110;
    x_137 = 'b111101111;
    x_138 = 'b111110100;
    x_139 = 'b111111111;
    x_140 = 'b000000101;
    x_141 = 'b111111001;
    x_142 = 'b111011111;
    x_143 = 'b111101000;
    x_144 = 'b111110001;
    x_145 = 'b111111100;
    x_146 = 'b000000010;
    x_147 = 'b000000110;
    x_148 = 'b000000010;
    x_149 = 'b111001010;
    x_150 = 'b111001100;
    x_151 = 'b111010110;
    x_152 = 'b111001000;
    x_153 = 'b111001001;
    x_154 = 'b111010111;
    x_155 = 'b111011111;
    x_156 = 'b111011011;
    x_157 = 'b111001110;
    x_158 = 'b111011110;
    x_159 = 'b111100000;
    x_160 = 'b111011110;
    x_161 = 'b111100011;
    x_162 = 'b111101111;
    x_163 = 'b111101110;
    x_164 = 'b111101110;
    x_165 = 'b111110010;
    x_166 = 'b111001100;
    x_167 = 'b111110011;
    x_168 = 'b111000101;
    x_169 = 'b111100111;
    x_170 = 'b111000010;
    x_171 = 'b111111011;
    x_172 = 'b111011100;
    x_173 = 'b111110001;
    x_174 = 'b111101101;
    x_175 = 'b111101101;
    x_176 = 'b111111000;
    x_177 = 'b111111010;
    x_178 = 'b000000110;
    x_179 = 'b000010101;
    x_180 = 'b000010001;
    x_181 = 'b000010011;
    x_182 = 'b000001111;
    x_183 = 'b111111001;
    x_184 = 'b111111100;
    x_185 = 'b000010110;
    x_186 = 'b000011000;
    x_187 = 'b000010100;
    x_188 = 'b111111000;
    x_189 = 'b000000101;
    x_190 = 'b111110111;
    x_191 = 'b111110001;
    x_192 = 'b111010001;
    x_193 = 'b111100100;
    x_194 = 'b111100111;
    x_195 = 'b111110111;
    x_196 = 'b111111011;
    x_197 = 'b111111100;
    x_198 = 'b111110010;
    x_199 = 'b111011111;
    x_200 = 'b111101110;
    x_201 = 'b111101111;
    x_202 = 'b111110100;
    x_203 = 'b111111111;
    x_204 = 'b000000101;
    x_205 = 'b111111001;
    x_206 = 'b111011111;
    x_207 = 'b111101000;
    x_208 = 'b111110001;
    x_209 = 'b111111100;
    x_210 = 'b000000010;
    x_211 = 'b000000110;
    x_212 = 'b000000010;
    x_213 = 'b111001010;
    x_214 = 'b111001100;
    x_215 = 'b111010110;
    x_216 = 'b111001000;
    x_217 = 'b111001001;
    x_218 = 'b111010111;
    x_219 = 'b111011111;
    x_220 = 'b111011011;
    x_221 = 'b111001110;
    x_222 = 'b111011110;
    x_223 = 'b111100000;
    x_224 = 'b111011110;
    x_225 = 'b111100011;
    x_226 = 'b111101111;
    x_227 = 'b111101110;
    x_228 = 'b111101110;
    x_229 = 'b111110010;
    x_230 = 'b111001100;
    x_231 = 'b111110011;
    x_232 = 'b111000101;
    x_233 = 'b111100111;
    x_234 = 'b111000010;
    x_235 = 'b111111011;
    x_236 = 'b111011100;
    x_237 = 'b111110001;
    x_238 = 'b111101101;
    x_239 = 'b111101101;
    x_240 = 'b111111000;
    x_241 = 'b111111010;
    x_242 = 'b000000110;
    x_243 = 'b000010101;
    x_244 = 'b000010001;
    x_245 = 'b000010011;
    x_246 = 'b000001111;
    x_247 = 'b111111001;
    x_248 = 'b111111100;
    x_249 = 'b000010110;
    x_250 = 'b000011000;
    x_251 = 'b000010100;
    x_252 = 'b111111000;
    x_253 = 'b000000101;
    x_254 = 'b111110111;
    x_255 = 'b111110001;

    h_0 = 'b111010001;
    h_1 = 'b111100100;
    h_2 = 'b111100111;
    h_3 = 'b111110111;
    h_4 = 'b111111011;
    h_5 = 'b111111100;
    h_6 = 'b111110010;
    h_7 = 'b111011111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111010101;
    x_1 = 'b111101010;
    x_2 = 'b111101010;
    x_3 = 'b111111011;
    x_4 = 'b000000100;
    x_5 = 'b000001001;
    x_6 = 'b111111010;
    x_7 = 'b111101011;
    x_8 = 'b111110010;
    x_9 = 'b111110100;
    x_10 = 'b111111100;
    x_11 = 'b000001011;
    x_12 = 'b000010011;
    x_13 = 'b000001001;
    x_14 = 'b111101000;
    x_15 = 'b111101011;
    x_16 = 'b111110101;
    x_17 = 'b000000100;
    x_18 = 'b000010001;
    x_19 = 'b000010101;
    x_20 = 'b000010011;
    x_21 = 'b111010001;
    x_22 = 'b111010100;
    x_23 = 'b111011010;
    x_24 = 'b111001110;
    x_25 = 'b111001111;
    x_26 = 'b111100000;
    x_27 = 'b111100111;
    x_28 = 'b111011111;
    x_29 = 'b111010100;
    x_30 = 'b111101010;
    x_31 = 'b111101011;
    x_32 = 'b111100100;
    x_33 = 'b111101010;
    x_34 = 'b111110111;
    x_35 = 'b111110111;
    x_36 = 'b111110111;
    x_37 = 'b111110010;
    x_38 = 'b111011101;
    x_39 = 'b111111011;
    x_40 = 'b111101000;
    x_41 = 'b111110101;
    x_42 = 'b111000111;
    x_43 = 'b000000101;
    x_44 = 'b111100101;
    x_45 = 'b000000001;
    x_46 = 'b111110110;
    x_47 = 'b111110011;
    x_48 = 'b111111010;
    x_49 = 'b000000010;
    x_50 = 'b000001110;
    x_51 = 'b000011110;
    x_52 = 'b000011000;
    x_53 = 'b000011010;
    x_54 = 'b000010110;
    x_55 = 'b000000001;
    x_56 = 'b000000011;
    x_57 = 'b000011011;
    x_58 = 'b000011110;
    x_59 = 'b000011001;
    x_60 = 'b000000010;
    x_61 = 'b000010001;
    x_62 = 'b000000010;
    x_63 = 'b111111110;
    x_64 = 'b111010101;
    x_65 = 'b111101010;
    x_66 = 'b111101010;
    x_67 = 'b111111011;
    x_68 = 'b000000100;
    x_69 = 'b000001001;
    x_70 = 'b111111010;
    x_71 = 'b111101011;
    x_72 = 'b111110010;
    x_73 = 'b111110100;
    x_74 = 'b111111100;
    x_75 = 'b000001011;
    x_76 = 'b000010011;
    x_77 = 'b000001001;
    x_78 = 'b111101000;
    x_79 = 'b111101011;
    x_80 = 'b111110101;
    x_81 = 'b000000100;
    x_82 = 'b000010001;
    x_83 = 'b000010101;
    x_84 = 'b000010011;
    x_85 = 'b111010001;
    x_86 = 'b111010100;
    x_87 = 'b111011010;
    x_88 = 'b111001110;
    x_89 = 'b111001111;
    x_90 = 'b111100000;
    x_91 = 'b111100111;
    x_92 = 'b111011111;
    x_93 = 'b111010100;
    x_94 = 'b111101010;
    x_95 = 'b111101011;
    x_96 = 'b111100100;
    x_97 = 'b111101010;
    x_98 = 'b111110111;
    x_99 = 'b111110111;
    x_100 = 'b111110111;
    x_101 = 'b111110010;
    x_102 = 'b111011101;
    x_103 = 'b111111011;
    x_104 = 'b111101000;
    x_105 = 'b111110101;
    x_106 = 'b111000111;
    x_107 = 'b000000101;
    x_108 = 'b111100101;
    x_109 = 'b000000001;
    x_110 = 'b111110110;
    x_111 = 'b111110011;
    x_112 = 'b111111010;
    x_113 = 'b000000010;
    x_114 = 'b000001110;
    x_115 = 'b000011110;
    x_116 = 'b000011000;
    x_117 = 'b000011010;
    x_118 = 'b000010110;
    x_119 = 'b000000001;
    x_120 = 'b000000011;
    x_121 = 'b000011011;
    x_122 = 'b000011110;
    x_123 = 'b000011001;
    x_124 = 'b000000010;
    x_125 = 'b000010001;
    x_126 = 'b000000010;
    x_127 = 'b111111110;
    x_128 = 'b111010101;
    x_129 = 'b111101010;
    x_130 = 'b111101010;
    x_131 = 'b111111011;
    x_132 = 'b000000100;
    x_133 = 'b000001001;
    x_134 = 'b111111010;
    x_135 = 'b111101011;
    x_136 = 'b111110010;
    x_137 = 'b111110100;
    x_138 = 'b111111100;
    x_139 = 'b000001011;
    x_140 = 'b000010011;
    x_141 = 'b000001001;
    x_142 = 'b111101000;
    x_143 = 'b111101011;
    x_144 = 'b111110101;
    x_145 = 'b000000100;
    x_146 = 'b000010001;
    x_147 = 'b000010101;
    x_148 = 'b000010011;
    x_149 = 'b111010001;
    x_150 = 'b111010100;
    x_151 = 'b111011010;
    x_152 = 'b111001110;
    x_153 = 'b111001111;
    x_154 = 'b111100000;
    x_155 = 'b111100111;
    x_156 = 'b111011111;
    x_157 = 'b111010100;
    x_158 = 'b111101010;
    x_159 = 'b111101011;
    x_160 = 'b111100100;
    x_161 = 'b111101010;
    x_162 = 'b111110111;
    x_163 = 'b111110111;
    x_164 = 'b111110111;
    x_165 = 'b111110010;
    x_166 = 'b111011101;
    x_167 = 'b111111011;
    x_168 = 'b111101000;
    x_169 = 'b111110101;
    x_170 = 'b111000111;
    x_171 = 'b000000101;
    x_172 = 'b111100101;
    x_173 = 'b000000001;
    x_174 = 'b111110110;
    x_175 = 'b111110011;
    x_176 = 'b111111010;
    x_177 = 'b000000010;
    x_178 = 'b000001110;
    x_179 = 'b000011110;
    x_180 = 'b000011000;
    x_181 = 'b000011010;
    x_182 = 'b000010110;
    x_183 = 'b000000001;
    x_184 = 'b000000011;
    x_185 = 'b000011011;
    x_186 = 'b000011110;
    x_187 = 'b000011001;
    x_188 = 'b000000010;
    x_189 = 'b000010001;
    x_190 = 'b000000010;
    x_191 = 'b111111110;
    x_192 = 'b111010101;
    x_193 = 'b111101010;
    x_194 = 'b111101010;
    x_195 = 'b111111011;
    x_196 = 'b000000100;
    x_197 = 'b000001001;
    x_198 = 'b111111010;
    x_199 = 'b111101011;
    x_200 = 'b111110010;
    x_201 = 'b111110100;
    x_202 = 'b111111100;
    x_203 = 'b000001011;
    x_204 = 'b000010011;
    x_205 = 'b000001001;
    x_206 = 'b111101000;
    x_207 = 'b111101011;
    x_208 = 'b111110101;
    x_209 = 'b000000100;
    x_210 = 'b000010001;
    x_211 = 'b000010101;
    x_212 = 'b000010011;
    x_213 = 'b111010001;
    x_214 = 'b111010100;
    x_215 = 'b111011010;
    x_216 = 'b111001110;
    x_217 = 'b111001111;
    x_218 = 'b111100000;
    x_219 = 'b111100111;
    x_220 = 'b111011111;
    x_221 = 'b111010100;
    x_222 = 'b111101010;
    x_223 = 'b111101011;
    x_224 = 'b111100100;
    x_225 = 'b111101010;
    x_226 = 'b111110111;
    x_227 = 'b111110111;
    x_228 = 'b111110111;
    x_229 = 'b111110010;
    x_230 = 'b111011101;
    x_231 = 'b111111011;
    x_232 = 'b111101000;
    x_233 = 'b111110101;
    x_234 = 'b111000111;
    x_235 = 'b000000101;
    x_236 = 'b111100101;
    x_237 = 'b000000001;
    x_238 = 'b111110110;
    x_239 = 'b111110011;
    x_240 = 'b111111010;
    x_241 = 'b000000010;
    x_242 = 'b000001110;
    x_243 = 'b000011110;
    x_244 = 'b000011000;
    x_245 = 'b000011010;
    x_246 = 'b000010110;
    x_247 = 'b000000001;
    x_248 = 'b000000011;
    x_249 = 'b000011011;
    x_250 = 'b000011110;
    x_251 = 'b000011001;
    x_252 = 'b000000010;
    x_253 = 'b000010001;
    x_254 = 'b000000010;
    x_255 = 'b111111110;

    h_0 = 'b111010101;
    h_1 = 'b111101010;
    h_2 = 'b111101010;
    h_3 = 'b111111011;
    h_4 = 'b000000100;
    h_5 = 'b000001001;
    h_6 = 'b111111010;
    h_7 = 'b111101011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111100100;
    x_1 = 'b111110010;
    x_2 = 'b111110000;
    x_3 = 'b000000000;
    x_4 = 'b000000110;
    x_5 = 'b000000111;
    x_6 = 'b111111100;
    x_7 = 'b111101110;
    x_8 = 'b111110010;
    x_9 = 'b111110111;
    x_10 = 'b111111111;
    x_11 = 'b000001001;
    x_12 = 'b000001110;
    x_13 = 'b000000001;
    x_14 = 'b111100001;
    x_15 = 'b111101010;
    x_16 = 'b111111000;
    x_17 = 'b000000101;
    x_18 = 'b000001101;
    x_19 = 'b000001110;
    x_20 = 'b000001010;
    x_21 = 'b111011000;
    x_22 = 'b111011001;
    x_23 = 'b111011101;
    x_24 = 'b111010101;
    x_25 = 'b111010110;
    x_26 = 'b111100110;
    x_27 = 'b111100111;
    x_28 = 'b111011101;
    x_29 = 'b111011011;
    x_30 = 'b111110011;
    x_31 = 'b111101011;
    x_32 = 'b111101011;
    x_33 = 'b111101110;
    x_34 = 'b111110111;
    x_35 = 'b111111000;
    x_36 = 'b111110001;
    x_37 = 'b111110010;
    x_38 = 'b111100101;
    x_39 = 'b111110011;
    x_40 = 'b111011110;
    x_41 = 'b000001011;
    x_42 = 'b111000110;
    x_43 = 'b111101110;
    x_44 = 'b111100111;
    x_45 = 'b111101001;
    x_46 = 'b111111000;
    x_47 = 'b111110001;
    x_48 = 'b111111010;
    x_49 = 'b111111101;
    x_50 = 'b000000111;
    x_51 = 'b000001100;
    x_52 = 'b000000101;
    x_53 = 'b000000101;
    x_54 = 'b111111100;
    x_55 = 'b111111101;
    x_56 = 'b111111110;
    x_57 = 'b000001110;
    x_58 = 'b000001001;
    x_59 = 'b000000010;
    x_60 = 'b000000111;
    x_61 = 'b000010000;
    x_62 = 'b111111111;
    x_63 = 'b111111011;
    x_64 = 'b111100100;
    x_65 = 'b111110010;
    x_66 = 'b111110000;
    x_67 = 'b000000000;
    x_68 = 'b000000110;
    x_69 = 'b000000111;
    x_70 = 'b111111100;
    x_71 = 'b111101110;
    x_72 = 'b111110010;
    x_73 = 'b111110111;
    x_74 = 'b111111111;
    x_75 = 'b000001001;
    x_76 = 'b000001110;
    x_77 = 'b000000001;
    x_78 = 'b111100001;
    x_79 = 'b111101010;
    x_80 = 'b111111000;
    x_81 = 'b000000101;
    x_82 = 'b000001101;
    x_83 = 'b000001110;
    x_84 = 'b000001010;
    x_85 = 'b111011000;
    x_86 = 'b111011001;
    x_87 = 'b111011101;
    x_88 = 'b111010101;
    x_89 = 'b111010110;
    x_90 = 'b111100110;
    x_91 = 'b111100111;
    x_92 = 'b111011101;
    x_93 = 'b111011011;
    x_94 = 'b111110011;
    x_95 = 'b111101011;
    x_96 = 'b111101011;
    x_97 = 'b111101110;
    x_98 = 'b111110111;
    x_99 = 'b111111000;
    x_100 = 'b111110001;
    x_101 = 'b111110010;
    x_102 = 'b111100101;
    x_103 = 'b111110011;
    x_104 = 'b111011110;
    x_105 = 'b000001011;
    x_106 = 'b111000110;
    x_107 = 'b111101110;
    x_108 = 'b111100111;
    x_109 = 'b111101001;
    x_110 = 'b111111000;
    x_111 = 'b111110001;
    x_112 = 'b111111010;
    x_113 = 'b111111101;
    x_114 = 'b000000111;
    x_115 = 'b000001100;
    x_116 = 'b000000101;
    x_117 = 'b000000101;
    x_118 = 'b111111100;
    x_119 = 'b111111101;
    x_120 = 'b111111110;
    x_121 = 'b000001110;
    x_122 = 'b000001001;
    x_123 = 'b000000010;
    x_124 = 'b000000111;
    x_125 = 'b000010000;
    x_126 = 'b111111111;
    x_127 = 'b111111011;
    x_128 = 'b111100100;
    x_129 = 'b111110010;
    x_130 = 'b111110000;
    x_131 = 'b000000000;
    x_132 = 'b000000110;
    x_133 = 'b000000111;
    x_134 = 'b111111100;
    x_135 = 'b111101110;
    x_136 = 'b111110010;
    x_137 = 'b111110111;
    x_138 = 'b111111111;
    x_139 = 'b000001001;
    x_140 = 'b000001110;
    x_141 = 'b000000001;
    x_142 = 'b111100001;
    x_143 = 'b111101010;
    x_144 = 'b111111000;
    x_145 = 'b000000101;
    x_146 = 'b000001101;
    x_147 = 'b000001110;
    x_148 = 'b000001010;
    x_149 = 'b111011000;
    x_150 = 'b111011001;
    x_151 = 'b111011101;
    x_152 = 'b111010101;
    x_153 = 'b111010110;
    x_154 = 'b111100110;
    x_155 = 'b111100111;
    x_156 = 'b111011101;
    x_157 = 'b111011011;
    x_158 = 'b111110011;
    x_159 = 'b111101011;
    x_160 = 'b111101011;
    x_161 = 'b111101110;
    x_162 = 'b111110111;
    x_163 = 'b111111000;
    x_164 = 'b111110001;
    x_165 = 'b111110010;
    x_166 = 'b111100101;
    x_167 = 'b111110011;
    x_168 = 'b111011110;
    x_169 = 'b000001011;
    x_170 = 'b111000110;
    x_171 = 'b111101110;
    x_172 = 'b111100111;
    x_173 = 'b111101001;
    x_174 = 'b111111000;
    x_175 = 'b111110001;
    x_176 = 'b111111010;
    x_177 = 'b111111101;
    x_178 = 'b000000111;
    x_179 = 'b000001100;
    x_180 = 'b000000101;
    x_181 = 'b000000101;
    x_182 = 'b111111100;
    x_183 = 'b111111101;
    x_184 = 'b111111110;
    x_185 = 'b000001110;
    x_186 = 'b000001001;
    x_187 = 'b000000010;
    x_188 = 'b000000111;
    x_189 = 'b000010000;
    x_190 = 'b111111111;
    x_191 = 'b111111011;
    x_192 = 'b111100100;
    x_193 = 'b111110010;
    x_194 = 'b111110000;
    x_195 = 'b000000000;
    x_196 = 'b000000110;
    x_197 = 'b000000111;
    x_198 = 'b111111100;
    x_199 = 'b111101110;
    x_200 = 'b111110010;
    x_201 = 'b111110111;
    x_202 = 'b111111111;
    x_203 = 'b000001001;
    x_204 = 'b000001110;
    x_205 = 'b000000001;
    x_206 = 'b111100001;
    x_207 = 'b111101010;
    x_208 = 'b111111000;
    x_209 = 'b000000101;
    x_210 = 'b000001101;
    x_211 = 'b000001110;
    x_212 = 'b000001010;
    x_213 = 'b111011000;
    x_214 = 'b111011001;
    x_215 = 'b111011101;
    x_216 = 'b111010101;
    x_217 = 'b111010110;
    x_218 = 'b111100110;
    x_219 = 'b111100111;
    x_220 = 'b111011101;
    x_221 = 'b111011011;
    x_222 = 'b111110011;
    x_223 = 'b111101011;
    x_224 = 'b111101011;
    x_225 = 'b111101110;
    x_226 = 'b111110111;
    x_227 = 'b111111000;
    x_228 = 'b111110001;
    x_229 = 'b111110010;
    x_230 = 'b111100101;
    x_231 = 'b111110011;
    x_232 = 'b111011110;
    x_233 = 'b000001011;
    x_234 = 'b111000110;
    x_235 = 'b111101110;
    x_236 = 'b111100111;
    x_237 = 'b111101001;
    x_238 = 'b111111000;
    x_239 = 'b111110001;
    x_240 = 'b111111010;
    x_241 = 'b111111101;
    x_242 = 'b000000111;
    x_243 = 'b000001100;
    x_244 = 'b000000101;
    x_245 = 'b000000101;
    x_246 = 'b111111100;
    x_247 = 'b111111101;
    x_248 = 'b111111110;
    x_249 = 'b000001110;
    x_250 = 'b000001001;
    x_251 = 'b000000010;
    x_252 = 'b000000111;
    x_253 = 'b000010000;
    x_254 = 'b111111111;
    x_255 = 'b111111011;

    h_0 = 'b111100100;
    h_1 = 'b111110010;
    h_2 = 'b111110000;
    h_3 = 'b000000000;
    h_4 = 'b000000110;
    h_5 = 'b000000111;
    h_6 = 'b111111100;
    h_7 = 'b111101110;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111100111;
    x_1 = 'b111111000;
    x_2 = 'b111110011;
    x_3 = 'b000000010;
    x_4 = 'b000000010;
    x_5 = 'b000000001;
    x_6 = 'b111111000;
    x_7 = 'b111110011;
    x_8 = 'b111110111;
    x_9 = 'b111111100;
    x_10 = 'b000000010;
    x_11 = 'b000001001;
    x_12 = 'b000001001;
    x_13 = 'b111111111;
    x_14 = 'b111101100;
    x_15 = 'b111110100;
    x_16 = 'b111111110;
    x_17 = 'b000001001;
    x_18 = 'b000000110;
    x_19 = 'b000000110;
    x_20 = 'b000000101;
    x_21 = 'b111011010;
    x_22 = 'b111011010;
    x_23 = 'b111100000;
    x_24 = 'b111011000;
    x_25 = 'b111011000;
    x_26 = 'b111101010;
    x_27 = 'b111101010;
    x_28 = 'b111100010;
    x_29 = 'b111011010;
    x_30 = 'b111110100;
    x_31 = 'b111101111;
    x_32 = 'b111101111;
    x_33 = 'b111110010;
    x_34 = 'b111111010;
    x_35 = 'b111111010;
    x_36 = 'b111110100;
    x_37 = 'b111111100;
    x_38 = 'b111011011;
    x_39 = 'b111111011;
    x_40 = 'b111011001;
    x_41 = 'b000011000;
    x_42 = 'b111001111;
    x_43 = 'b111100111;
    x_44 = 'b111101100;
    x_45 = 'b111110010;
    x_46 = 'b111111110;
    x_47 = 'b111111111;
    x_48 = 'b000001001;
    x_49 = 'b000001000;
    x_50 = 'b000001100;
    x_51 = 'b000001101;
    x_52 = 'b000000111;
    x_53 = 'b000000111;
    x_54 = 'b000000101;
    x_55 = 'b000001101;
    x_56 = 'b000001011;
    x_57 = 'b000010101;
    x_58 = 'b000001001;
    x_59 = 'b000000101;
    x_60 = 'b000001100;
    x_61 = 'b000001100;
    x_62 = 'b111111001;
    x_63 = 'b111111010;
    x_64 = 'b111100111;
    x_65 = 'b111111000;
    x_66 = 'b111110011;
    x_67 = 'b000000010;
    x_68 = 'b000000010;
    x_69 = 'b000000001;
    x_70 = 'b111111000;
    x_71 = 'b111110011;
    x_72 = 'b111110111;
    x_73 = 'b111111100;
    x_74 = 'b000000010;
    x_75 = 'b000001001;
    x_76 = 'b000001001;
    x_77 = 'b111111111;
    x_78 = 'b111101100;
    x_79 = 'b111110100;
    x_80 = 'b111111110;
    x_81 = 'b000001001;
    x_82 = 'b000000110;
    x_83 = 'b000000110;
    x_84 = 'b000000101;
    x_85 = 'b111011010;
    x_86 = 'b111011010;
    x_87 = 'b111100000;
    x_88 = 'b111011000;
    x_89 = 'b111011000;
    x_90 = 'b111101010;
    x_91 = 'b111101010;
    x_92 = 'b111100010;
    x_93 = 'b111011010;
    x_94 = 'b111110100;
    x_95 = 'b111101111;
    x_96 = 'b111101111;
    x_97 = 'b111110010;
    x_98 = 'b111111010;
    x_99 = 'b111111010;
    x_100 = 'b111110100;
    x_101 = 'b111111100;
    x_102 = 'b111011011;
    x_103 = 'b111111011;
    x_104 = 'b111011001;
    x_105 = 'b000011000;
    x_106 = 'b111001111;
    x_107 = 'b111100111;
    x_108 = 'b111101100;
    x_109 = 'b111110010;
    x_110 = 'b111111110;
    x_111 = 'b111111111;
    x_112 = 'b000001001;
    x_113 = 'b000001000;
    x_114 = 'b000001100;
    x_115 = 'b000001101;
    x_116 = 'b000000111;
    x_117 = 'b000000111;
    x_118 = 'b000000101;
    x_119 = 'b000001101;
    x_120 = 'b000001011;
    x_121 = 'b000010101;
    x_122 = 'b000001001;
    x_123 = 'b000000101;
    x_124 = 'b000001100;
    x_125 = 'b000001100;
    x_126 = 'b111111001;
    x_127 = 'b111111010;
    x_128 = 'b111100111;
    x_129 = 'b111111000;
    x_130 = 'b111110011;
    x_131 = 'b000000010;
    x_132 = 'b000000010;
    x_133 = 'b000000001;
    x_134 = 'b111111000;
    x_135 = 'b111110011;
    x_136 = 'b111110111;
    x_137 = 'b111111100;
    x_138 = 'b000000010;
    x_139 = 'b000001001;
    x_140 = 'b000001001;
    x_141 = 'b111111111;
    x_142 = 'b111101100;
    x_143 = 'b111110100;
    x_144 = 'b111111110;
    x_145 = 'b000001001;
    x_146 = 'b000000110;
    x_147 = 'b000000110;
    x_148 = 'b000000101;
    x_149 = 'b111011010;
    x_150 = 'b111011010;
    x_151 = 'b111100000;
    x_152 = 'b111011000;
    x_153 = 'b111011000;
    x_154 = 'b111101010;
    x_155 = 'b111101010;
    x_156 = 'b111100010;
    x_157 = 'b111011010;
    x_158 = 'b111110100;
    x_159 = 'b111101111;
    x_160 = 'b111101111;
    x_161 = 'b111110010;
    x_162 = 'b111111010;
    x_163 = 'b111111010;
    x_164 = 'b111110100;
    x_165 = 'b111111100;
    x_166 = 'b111011011;
    x_167 = 'b111111011;
    x_168 = 'b111011001;
    x_169 = 'b000011000;
    x_170 = 'b111001111;
    x_171 = 'b111100111;
    x_172 = 'b111101100;
    x_173 = 'b111110010;
    x_174 = 'b111111110;
    x_175 = 'b111111111;
    x_176 = 'b000001001;
    x_177 = 'b000001000;
    x_178 = 'b000001100;
    x_179 = 'b000001101;
    x_180 = 'b000000111;
    x_181 = 'b000000111;
    x_182 = 'b000000101;
    x_183 = 'b000001101;
    x_184 = 'b000001011;
    x_185 = 'b000010101;
    x_186 = 'b000001001;
    x_187 = 'b000000101;
    x_188 = 'b000001100;
    x_189 = 'b000001100;
    x_190 = 'b111111001;
    x_191 = 'b111111010;
    x_192 = 'b111100111;
    x_193 = 'b111111000;
    x_194 = 'b111110011;
    x_195 = 'b000000010;
    x_196 = 'b000000010;
    x_197 = 'b000000001;
    x_198 = 'b111111000;
    x_199 = 'b111110011;
    x_200 = 'b111110111;
    x_201 = 'b111111100;
    x_202 = 'b000000010;
    x_203 = 'b000001001;
    x_204 = 'b000001001;
    x_205 = 'b111111111;
    x_206 = 'b111101100;
    x_207 = 'b111110100;
    x_208 = 'b111111110;
    x_209 = 'b000001001;
    x_210 = 'b000000110;
    x_211 = 'b000000110;
    x_212 = 'b000000101;
    x_213 = 'b111011010;
    x_214 = 'b111011010;
    x_215 = 'b111100000;
    x_216 = 'b111011000;
    x_217 = 'b111011000;
    x_218 = 'b111101010;
    x_219 = 'b111101010;
    x_220 = 'b111100010;
    x_221 = 'b111011010;
    x_222 = 'b111110100;
    x_223 = 'b111101111;
    x_224 = 'b111101111;
    x_225 = 'b111110010;
    x_226 = 'b111111010;
    x_227 = 'b111111010;
    x_228 = 'b111110100;
    x_229 = 'b111111100;
    x_230 = 'b111011011;
    x_231 = 'b111111011;
    x_232 = 'b111011001;
    x_233 = 'b000011000;
    x_234 = 'b111001111;
    x_235 = 'b111100111;
    x_236 = 'b111101100;
    x_237 = 'b111110010;
    x_238 = 'b111111110;
    x_239 = 'b111111111;
    x_240 = 'b000001001;
    x_241 = 'b000001000;
    x_242 = 'b000001100;
    x_243 = 'b000001101;
    x_244 = 'b000000111;
    x_245 = 'b000000111;
    x_246 = 'b000000101;
    x_247 = 'b000001101;
    x_248 = 'b000001011;
    x_249 = 'b000010101;
    x_250 = 'b000001001;
    x_251 = 'b000000101;
    x_252 = 'b000001100;
    x_253 = 'b000001100;
    x_254 = 'b111111001;
    x_255 = 'b111111010;

    h_0 = 'b111100111;
    h_1 = 'b111111000;
    h_2 = 'b111110011;
    h_3 = 'b000000010;
    h_4 = 'b000000010;
    h_5 = 'b000000001;
    h_6 = 'b111111000;
    h_7 = 'b111110011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111100100;
    x_1 = 'b111111010;
    x_2 = 'b111110100;
    x_3 = 'b000000010;
    x_4 = 'b000000001;
    x_5 = 'b000000100;
    x_6 = 'b111111010;
    x_7 = 'b111111100;
    x_8 = 'b000000000;
    x_9 = 'b111111110;
    x_10 = 'b111111111;
    x_11 = 'b000001001;
    x_12 = 'b000000110;
    x_13 = 'b000000001;
    x_14 = 'b111110111;
    x_15 = 'b111111101;
    x_16 = 'b000000000;
    x_17 = 'b000000100;
    x_18 = 'b000000000;
    x_19 = 'b111111111;
    x_20 = 'b000000010;
    x_21 = 'b111011011;
    x_22 = 'b111011101;
    x_23 = 'b111100010;
    x_24 = 'b111010101;
    x_25 = 'b111010110;
    x_26 = 'b111101010;
    x_27 = 'b111101011;
    x_28 = 'b111100101;
    x_29 = 'b111010110;
    x_30 = 'b111101100;
    x_31 = 'b111101010;
    x_32 = 'b111101001;
    x_33 = 'b111101100;
    x_34 = 'b111110101;
    x_35 = 'b111110011;
    x_36 = 'b111110001;
    x_37 = 'b111110101;
    x_38 = 'b111011111;
    x_39 = 'b111101111;
    x_40 = 'b111100111;
    x_41 = 'b111101100;
    x_42 = 'b111010111;
    x_43 = 'b111011011;
    x_44 = 'b111101110;
    x_45 = 'b111100100;
    x_46 = 'b111111110;
    x_47 = 'b111111100;
    x_48 = 'b000000011;
    x_49 = 'b111111101;
    x_50 = 'b111111010;
    x_51 = 'b111111010;
    x_52 = 'b111110001;
    x_53 = 'b111110111;
    x_54 = 'b111110110;
    x_55 = 'b000000111;
    x_56 = 'b000000011;
    x_57 = 'b000000101;
    x_58 = 'b111110111;
    x_59 = 'b111111100;
    x_60 = 'b000001101;
    x_61 = 'b000000111;
    x_62 = 'b111110101;
    x_63 = 'b111111101;
    x_64 = 'b111100100;
    x_65 = 'b111111010;
    x_66 = 'b111110100;
    x_67 = 'b000000010;
    x_68 = 'b000000001;
    x_69 = 'b000000100;
    x_70 = 'b111111010;
    x_71 = 'b111111100;
    x_72 = 'b000000000;
    x_73 = 'b111111110;
    x_74 = 'b111111111;
    x_75 = 'b000001001;
    x_76 = 'b000000110;
    x_77 = 'b000000001;
    x_78 = 'b111110111;
    x_79 = 'b111111101;
    x_80 = 'b000000000;
    x_81 = 'b000000100;
    x_82 = 'b000000000;
    x_83 = 'b111111111;
    x_84 = 'b000000010;
    x_85 = 'b111011011;
    x_86 = 'b111011101;
    x_87 = 'b111100010;
    x_88 = 'b111010101;
    x_89 = 'b111010110;
    x_90 = 'b111101010;
    x_91 = 'b111101011;
    x_92 = 'b111100101;
    x_93 = 'b111010110;
    x_94 = 'b111101100;
    x_95 = 'b111101010;
    x_96 = 'b111101001;
    x_97 = 'b111101100;
    x_98 = 'b111110101;
    x_99 = 'b111110011;
    x_100 = 'b111110001;
    x_101 = 'b111110101;
    x_102 = 'b111011111;
    x_103 = 'b111101111;
    x_104 = 'b111100111;
    x_105 = 'b111101100;
    x_106 = 'b111010111;
    x_107 = 'b111011011;
    x_108 = 'b111101110;
    x_109 = 'b111100100;
    x_110 = 'b111111110;
    x_111 = 'b111111100;
    x_112 = 'b000000011;
    x_113 = 'b111111101;
    x_114 = 'b111111010;
    x_115 = 'b111111010;
    x_116 = 'b111110001;
    x_117 = 'b111110111;
    x_118 = 'b111110110;
    x_119 = 'b000000111;
    x_120 = 'b000000011;
    x_121 = 'b000000101;
    x_122 = 'b111110111;
    x_123 = 'b111111100;
    x_124 = 'b000001101;
    x_125 = 'b000000111;
    x_126 = 'b111110101;
    x_127 = 'b111111101;
    x_128 = 'b111100100;
    x_129 = 'b111111010;
    x_130 = 'b111110100;
    x_131 = 'b000000010;
    x_132 = 'b000000001;
    x_133 = 'b000000100;
    x_134 = 'b111111010;
    x_135 = 'b111111100;
    x_136 = 'b000000000;
    x_137 = 'b111111110;
    x_138 = 'b111111111;
    x_139 = 'b000001001;
    x_140 = 'b000000110;
    x_141 = 'b000000001;
    x_142 = 'b111110111;
    x_143 = 'b111111101;
    x_144 = 'b000000000;
    x_145 = 'b000000100;
    x_146 = 'b000000000;
    x_147 = 'b111111111;
    x_148 = 'b000000010;
    x_149 = 'b111011011;
    x_150 = 'b111011101;
    x_151 = 'b111100010;
    x_152 = 'b111010101;
    x_153 = 'b111010110;
    x_154 = 'b111101010;
    x_155 = 'b111101011;
    x_156 = 'b111100101;
    x_157 = 'b111010110;
    x_158 = 'b111101100;
    x_159 = 'b111101010;
    x_160 = 'b111101001;
    x_161 = 'b111101100;
    x_162 = 'b111110101;
    x_163 = 'b111110011;
    x_164 = 'b111110001;
    x_165 = 'b111110101;
    x_166 = 'b111011111;
    x_167 = 'b111101111;
    x_168 = 'b111100111;
    x_169 = 'b111101100;
    x_170 = 'b111010111;
    x_171 = 'b111011011;
    x_172 = 'b111101110;
    x_173 = 'b111100100;
    x_174 = 'b111111110;
    x_175 = 'b111111100;
    x_176 = 'b000000011;
    x_177 = 'b111111101;
    x_178 = 'b111111010;
    x_179 = 'b111111010;
    x_180 = 'b111110001;
    x_181 = 'b111110111;
    x_182 = 'b111110110;
    x_183 = 'b000000111;
    x_184 = 'b000000011;
    x_185 = 'b000000101;
    x_186 = 'b111110111;
    x_187 = 'b111111100;
    x_188 = 'b000001101;
    x_189 = 'b000000111;
    x_190 = 'b111110101;
    x_191 = 'b111111101;
    x_192 = 'b111100100;
    x_193 = 'b111111010;
    x_194 = 'b111110100;
    x_195 = 'b000000010;
    x_196 = 'b000000001;
    x_197 = 'b000000100;
    x_198 = 'b111111010;
    x_199 = 'b111111100;
    x_200 = 'b000000000;
    x_201 = 'b111111110;
    x_202 = 'b111111111;
    x_203 = 'b000001001;
    x_204 = 'b000000110;
    x_205 = 'b000000001;
    x_206 = 'b111110111;
    x_207 = 'b111111101;
    x_208 = 'b000000000;
    x_209 = 'b000000100;
    x_210 = 'b000000000;
    x_211 = 'b111111111;
    x_212 = 'b000000010;
    x_213 = 'b111011011;
    x_214 = 'b111011101;
    x_215 = 'b111100010;
    x_216 = 'b111010101;
    x_217 = 'b111010110;
    x_218 = 'b111101010;
    x_219 = 'b111101011;
    x_220 = 'b111100101;
    x_221 = 'b111010110;
    x_222 = 'b111101100;
    x_223 = 'b111101010;
    x_224 = 'b111101001;
    x_225 = 'b111101100;
    x_226 = 'b111110101;
    x_227 = 'b111110011;
    x_228 = 'b111110001;
    x_229 = 'b111110101;
    x_230 = 'b111011111;
    x_231 = 'b111101111;
    x_232 = 'b111100111;
    x_233 = 'b111101100;
    x_234 = 'b111010111;
    x_235 = 'b111011011;
    x_236 = 'b111101110;
    x_237 = 'b111100100;
    x_238 = 'b111111110;
    x_239 = 'b111111100;
    x_240 = 'b000000011;
    x_241 = 'b111111101;
    x_242 = 'b111111010;
    x_243 = 'b111111010;
    x_244 = 'b111110001;
    x_245 = 'b111110111;
    x_246 = 'b111110110;
    x_247 = 'b000000111;
    x_248 = 'b000000011;
    x_249 = 'b000000101;
    x_250 = 'b111110111;
    x_251 = 'b111111100;
    x_252 = 'b000001101;
    x_253 = 'b000000111;
    x_254 = 'b111110101;
    x_255 = 'b111111101;

    h_0 = 'b111100100;
    h_1 = 'b111111010;
    h_2 = 'b111110100;
    h_3 = 'b000000010;
    h_4 = 'b000000001;
    h_5 = 'b000000100;
    h_6 = 'b111111010;
    h_7 = 'b111111100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111011101;
    x_1 = 'b111101000;
    x_2 = 'b111100111;
    x_3 = 'b111110111;
    x_4 = 'b111110110;
    x_5 = 'b111110011;
    x_6 = 'b111101011;
    x_7 = 'b111101100;
    x_8 = 'b111110001;
    x_9 = 'b111101110;
    x_10 = 'b111101111;
    x_11 = 'b111111010;
    x_12 = 'b111110011;
    x_13 = 'b111101001;
    x_14 = 'b111101110;
    x_15 = 'b111110000;
    x_16 = 'b111110001;
    x_17 = 'b111110001;
    x_18 = 'b111101101;
    x_19 = 'b111101110;
    x_20 = 'b111110000;
    x_21 = 'b111011011;
    x_22 = 'b111011100;
    x_23 = 'b111100001;
    x_24 = 'b111010110;
    x_25 = 'b111010110;
    x_26 = 'b111101010;
    x_27 = 'b111101000;
    x_28 = 'b111100010;
    x_29 = 'b111011001;
    x_30 = 'b111101100;
    x_31 = 'b111100110;
    x_32 = 'b111101010;
    x_33 = 'b111101111;
    x_34 = 'b111110110;
    x_35 = 'b111110011;
    x_36 = 'b111101100;
    x_37 = 'b111110001;
    x_38 = 'b111101101;
    x_39 = 'b111101010;
    x_40 = 'b111110100;
    x_41 = 'b111100010;
    x_42 = 'b111101010;
    x_43 = 'b111100111;
    x_44 = 'b111110000;
    x_45 = 'b111101100;
    x_46 = 'b000000001;
    x_47 = 'b111111110;
    x_48 = 'b000000010;
    x_49 = 'b111111010;
    x_50 = 'b111110110;
    x_51 = 'b111110110;
    x_52 = 'b111110010;
    x_53 = 'b111111101;
    x_54 = 'b000000000;
    x_55 = 'b000001100;
    x_56 = 'b000001000;
    x_57 = 'b000000100;
    x_58 = 'b111111010;
    x_59 = 'b000000110;
    x_60 = 'b000001100;
    x_61 = 'b000000110;
    x_62 = 'b111110111;
    x_63 = 'b000000111;
    x_64 = 'b111011101;
    x_65 = 'b111101000;
    x_66 = 'b111100111;
    x_67 = 'b111110111;
    x_68 = 'b111110110;
    x_69 = 'b111110011;
    x_70 = 'b111101011;
    x_71 = 'b111101100;
    x_72 = 'b111110001;
    x_73 = 'b111101110;
    x_74 = 'b111101111;
    x_75 = 'b111111010;
    x_76 = 'b111110011;
    x_77 = 'b111101001;
    x_78 = 'b111101110;
    x_79 = 'b111110000;
    x_80 = 'b111110001;
    x_81 = 'b111110001;
    x_82 = 'b111101101;
    x_83 = 'b111101110;
    x_84 = 'b111110000;
    x_85 = 'b111011011;
    x_86 = 'b111011100;
    x_87 = 'b111100001;
    x_88 = 'b111010110;
    x_89 = 'b111010110;
    x_90 = 'b111101010;
    x_91 = 'b111101000;
    x_92 = 'b111100010;
    x_93 = 'b111011001;
    x_94 = 'b111101100;
    x_95 = 'b111100110;
    x_96 = 'b111101010;
    x_97 = 'b111101111;
    x_98 = 'b111110110;
    x_99 = 'b111110011;
    x_100 = 'b111101100;
    x_101 = 'b111110001;
    x_102 = 'b111101101;
    x_103 = 'b111101010;
    x_104 = 'b111110100;
    x_105 = 'b111100010;
    x_106 = 'b111101010;
    x_107 = 'b111100111;
    x_108 = 'b111110000;
    x_109 = 'b111101100;
    x_110 = 'b000000001;
    x_111 = 'b111111110;
    x_112 = 'b000000010;
    x_113 = 'b111111010;
    x_114 = 'b111110110;
    x_115 = 'b111110110;
    x_116 = 'b111110010;
    x_117 = 'b111111101;
    x_118 = 'b000000000;
    x_119 = 'b000001100;
    x_120 = 'b000001000;
    x_121 = 'b000000100;
    x_122 = 'b111111010;
    x_123 = 'b000000110;
    x_124 = 'b000001100;
    x_125 = 'b000000110;
    x_126 = 'b111110111;
    x_127 = 'b000000111;
    x_128 = 'b111011101;
    x_129 = 'b111101000;
    x_130 = 'b111100111;
    x_131 = 'b111110111;
    x_132 = 'b111110110;
    x_133 = 'b111110011;
    x_134 = 'b111101011;
    x_135 = 'b111101100;
    x_136 = 'b111110001;
    x_137 = 'b111101110;
    x_138 = 'b111101111;
    x_139 = 'b111111010;
    x_140 = 'b111110011;
    x_141 = 'b111101001;
    x_142 = 'b111101110;
    x_143 = 'b111110000;
    x_144 = 'b111110001;
    x_145 = 'b111110001;
    x_146 = 'b111101101;
    x_147 = 'b111101110;
    x_148 = 'b111110000;
    x_149 = 'b111011011;
    x_150 = 'b111011100;
    x_151 = 'b111100001;
    x_152 = 'b111010110;
    x_153 = 'b111010110;
    x_154 = 'b111101010;
    x_155 = 'b111101000;
    x_156 = 'b111100010;
    x_157 = 'b111011001;
    x_158 = 'b111101100;
    x_159 = 'b111100110;
    x_160 = 'b111101010;
    x_161 = 'b111101111;
    x_162 = 'b111110110;
    x_163 = 'b111110011;
    x_164 = 'b111101100;
    x_165 = 'b111110001;
    x_166 = 'b111101101;
    x_167 = 'b111101010;
    x_168 = 'b111110100;
    x_169 = 'b111100010;
    x_170 = 'b111101010;
    x_171 = 'b111100111;
    x_172 = 'b111110000;
    x_173 = 'b111101100;
    x_174 = 'b000000001;
    x_175 = 'b111111110;
    x_176 = 'b000000010;
    x_177 = 'b111111010;
    x_178 = 'b111110110;
    x_179 = 'b111110110;
    x_180 = 'b111110010;
    x_181 = 'b111111101;
    x_182 = 'b000000000;
    x_183 = 'b000001100;
    x_184 = 'b000001000;
    x_185 = 'b000000100;
    x_186 = 'b111111010;
    x_187 = 'b000000110;
    x_188 = 'b000001100;
    x_189 = 'b000000110;
    x_190 = 'b111110111;
    x_191 = 'b000000111;
    x_192 = 'b111011101;
    x_193 = 'b111101000;
    x_194 = 'b111100111;
    x_195 = 'b111110111;
    x_196 = 'b111110110;
    x_197 = 'b111110011;
    x_198 = 'b111101011;
    x_199 = 'b111101100;
    x_200 = 'b111110001;
    x_201 = 'b111101110;
    x_202 = 'b111101111;
    x_203 = 'b111111010;
    x_204 = 'b111110011;
    x_205 = 'b111101001;
    x_206 = 'b111101110;
    x_207 = 'b111110000;
    x_208 = 'b111110001;
    x_209 = 'b111110001;
    x_210 = 'b111101101;
    x_211 = 'b111101110;
    x_212 = 'b111110000;
    x_213 = 'b111011011;
    x_214 = 'b111011100;
    x_215 = 'b111100001;
    x_216 = 'b111010110;
    x_217 = 'b111010110;
    x_218 = 'b111101010;
    x_219 = 'b111101000;
    x_220 = 'b111100010;
    x_221 = 'b111011001;
    x_222 = 'b111101100;
    x_223 = 'b111100110;
    x_224 = 'b111101010;
    x_225 = 'b111101111;
    x_226 = 'b111110110;
    x_227 = 'b111110011;
    x_228 = 'b111101100;
    x_229 = 'b111110001;
    x_230 = 'b111101101;
    x_231 = 'b111101010;
    x_232 = 'b111110100;
    x_233 = 'b111100010;
    x_234 = 'b111101010;
    x_235 = 'b111100111;
    x_236 = 'b111110000;
    x_237 = 'b111101100;
    x_238 = 'b000000001;
    x_239 = 'b111111110;
    x_240 = 'b000000010;
    x_241 = 'b111111010;
    x_242 = 'b111110110;
    x_243 = 'b111110110;
    x_244 = 'b111110010;
    x_245 = 'b111111101;
    x_246 = 'b000000000;
    x_247 = 'b000001100;
    x_248 = 'b000001000;
    x_249 = 'b000000100;
    x_250 = 'b111111010;
    x_251 = 'b000000110;
    x_252 = 'b000001100;
    x_253 = 'b000000110;
    x_254 = 'b111110111;
    x_255 = 'b000000111;

    h_0 = 'b111011101;
    h_1 = 'b111101000;
    h_2 = 'b111100111;
    h_3 = 'b111110111;
    h_4 = 'b111110110;
    h_5 = 'b111110011;
    h_6 = 'b111101011;
    h_7 = 'b111101100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111110001;
    x_1 = 'b111111011;
    x_2 = 'b111111000;
    x_3 = 'b000000111;
    x_4 = 'b000000110;
    x_5 = 'b000000001;
    x_6 = 'b111110101;
    x_7 = 'b000001011;
    x_8 = 'b000000110;
    x_9 = 'b000000000;
    x_10 = 'b000000001;
    x_11 = 'b000001101;
    x_12 = 'b000000100;
    x_13 = 'b111111001;
    x_14 = 'b000000011;
    x_15 = 'b000000101;
    x_16 = 'b000000010;
    x_17 = 'b000000010;
    x_18 = 'b111111100;
    x_19 = 'b111111111;
    x_20 = 'b000000100;
    x_21 = 'b111100011;
    x_22 = 'b111100101;
    x_23 = 'b111100111;
    x_24 = 'b111100010;
    x_25 = 'b111100010;
    x_26 = 'b111110101;
    x_27 = 'b111110010;
    x_28 = 'b111100111;
    x_29 = 'b111101001;
    x_30 = 'b000000000;
    x_31 = 'b111110110;
    x_32 = 'b111110111;
    x_33 = 'b111111010;
    x_34 = 'b000000011;
    x_35 = 'b111111111;
    x_36 = 'b111110111;
    x_37 = 'b111111001;
    x_38 = 'b111111100;
    x_39 = 'b111101101;
    x_40 = 'b000000010;
    x_41 = 'b111110000;
    x_42 = 'b111101000;
    x_43 = 'b111111101;
    x_44 = 'b000000000;
    x_45 = 'b111110010;
    x_46 = 'b000001011;
    x_47 = 'b000001000;
    x_48 = 'b000001100;
    x_49 = 'b000000001;
    x_50 = 'b111111010;
    x_51 = 'b111111000;
    x_52 = 'b111110010;
    x_53 = 'b111111011;
    x_54 = 'b111111101;
    x_55 = 'b000001110;
    x_56 = 'b000001010;
    x_57 = 'b000000010;
    x_58 = 'b111110110;
    x_59 = 'b111111010;
    x_60 = 'b000001110;
    x_61 = 'b000001010;
    x_62 = 'b111110111;
    x_63 = 'b000010010;
    x_64 = 'b111110001;
    x_65 = 'b111111011;
    x_66 = 'b111111000;
    x_67 = 'b000000111;
    x_68 = 'b000000110;
    x_69 = 'b000000001;
    x_70 = 'b111110101;
    x_71 = 'b000001011;
    x_72 = 'b000000110;
    x_73 = 'b000000000;
    x_74 = 'b000000001;
    x_75 = 'b000001101;
    x_76 = 'b000000100;
    x_77 = 'b111111001;
    x_78 = 'b000000011;
    x_79 = 'b000000101;
    x_80 = 'b000000010;
    x_81 = 'b000000010;
    x_82 = 'b111111100;
    x_83 = 'b111111111;
    x_84 = 'b000000100;
    x_85 = 'b111100011;
    x_86 = 'b111100101;
    x_87 = 'b111100111;
    x_88 = 'b111100010;
    x_89 = 'b111100010;
    x_90 = 'b111110101;
    x_91 = 'b111110010;
    x_92 = 'b111100111;
    x_93 = 'b111101001;
    x_94 = 'b000000000;
    x_95 = 'b111110110;
    x_96 = 'b111110111;
    x_97 = 'b111111010;
    x_98 = 'b000000011;
    x_99 = 'b111111111;
    x_100 = 'b111110111;
    x_101 = 'b111111001;
    x_102 = 'b111111100;
    x_103 = 'b111101101;
    x_104 = 'b000000010;
    x_105 = 'b111110000;
    x_106 = 'b111101000;
    x_107 = 'b111111101;
    x_108 = 'b000000000;
    x_109 = 'b111110010;
    x_110 = 'b000001011;
    x_111 = 'b000001000;
    x_112 = 'b000001100;
    x_113 = 'b000000001;
    x_114 = 'b111111010;
    x_115 = 'b111111000;
    x_116 = 'b111110010;
    x_117 = 'b111111011;
    x_118 = 'b111111101;
    x_119 = 'b000001110;
    x_120 = 'b000001010;
    x_121 = 'b000000010;
    x_122 = 'b111110110;
    x_123 = 'b111111010;
    x_124 = 'b000001110;
    x_125 = 'b000001010;
    x_126 = 'b111110111;
    x_127 = 'b000010010;
    x_128 = 'b111110001;
    x_129 = 'b111111011;
    x_130 = 'b111111000;
    x_131 = 'b000000111;
    x_132 = 'b000000110;
    x_133 = 'b000000001;
    x_134 = 'b111110101;
    x_135 = 'b000001011;
    x_136 = 'b000000110;
    x_137 = 'b000000000;
    x_138 = 'b000000001;
    x_139 = 'b000001101;
    x_140 = 'b000000100;
    x_141 = 'b111111001;
    x_142 = 'b000000011;
    x_143 = 'b000000101;
    x_144 = 'b000000010;
    x_145 = 'b000000010;
    x_146 = 'b111111100;
    x_147 = 'b111111111;
    x_148 = 'b000000100;
    x_149 = 'b111100011;
    x_150 = 'b111100101;
    x_151 = 'b111100111;
    x_152 = 'b111100010;
    x_153 = 'b111100010;
    x_154 = 'b111110101;
    x_155 = 'b111110010;
    x_156 = 'b111100111;
    x_157 = 'b111101001;
    x_158 = 'b000000000;
    x_159 = 'b111110110;
    x_160 = 'b111110111;
    x_161 = 'b111111010;
    x_162 = 'b000000011;
    x_163 = 'b111111111;
    x_164 = 'b111110111;
    x_165 = 'b111111001;
    x_166 = 'b111111100;
    x_167 = 'b111101101;
    x_168 = 'b000000010;
    x_169 = 'b111110000;
    x_170 = 'b111101000;
    x_171 = 'b111111101;
    x_172 = 'b000000000;
    x_173 = 'b111110010;
    x_174 = 'b000001011;
    x_175 = 'b000001000;
    x_176 = 'b000001100;
    x_177 = 'b000000001;
    x_178 = 'b111111010;
    x_179 = 'b111111000;
    x_180 = 'b111110010;
    x_181 = 'b111111011;
    x_182 = 'b111111101;
    x_183 = 'b000001110;
    x_184 = 'b000001010;
    x_185 = 'b000000010;
    x_186 = 'b111110110;
    x_187 = 'b111111010;
    x_188 = 'b000001110;
    x_189 = 'b000001010;
    x_190 = 'b111110111;
    x_191 = 'b000010010;
    x_192 = 'b111110001;
    x_193 = 'b111111011;
    x_194 = 'b111111000;
    x_195 = 'b000000111;
    x_196 = 'b000000110;
    x_197 = 'b000000001;
    x_198 = 'b111110101;
    x_199 = 'b000001011;
    x_200 = 'b000000110;
    x_201 = 'b000000000;
    x_202 = 'b000000001;
    x_203 = 'b000001101;
    x_204 = 'b000000100;
    x_205 = 'b111111001;
    x_206 = 'b000000011;
    x_207 = 'b000000101;
    x_208 = 'b000000010;
    x_209 = 'b000000010;
    x_210 = 'b111111100;
    x_211 = 'b111111111;
    x_212 = 'b000000100;
    x_213 = 'b111100011;
    x_214 = 'b111100101;
    x_215 = 'b111100111;
    x_216 = 'b111100010;
    x_217 = 'b111100010;
    x_218 = 'b111110101;
    x_219 = 'b111110010;
    x_220 = 'b111100111;
    x_221 = 'b111101001;
    x_222 = 'b000000000;
    x_223 = 'b111110110;
    x_224 = 'b111110111;
    x_225 = 'b111111010;
    x_226 = 'b000000011;
    x_227 = 'b111111111;
    x_228 = 'b111110111;
    x_229 = 'b111111001;
    x_230 = 'b111111100;
    x_231 = 'b111101101;
    x_232 = 'b000000010;
    x_233 = 'b111110000;
    x_234 = 'b111101000;
    x_235 = 'b111111101;
    x_236 = 'b000000000;
    x_237 = 'b111110010;
    x_238 = 'b000001011;
    x_239 = 'b000001000;
    x_240 = 'b000001100;
    x_241 = 'b000000001;
    x_242 = 'b111111010;
    x_243 = 'b111111000;
    x_244 = 'b111110010;
    x_245 = 'b111111011;
    x_246 = 'b111111101;
    x_247 = 'b000001110;
    x_248 = 'b000001010;
    x_249 = 'b000000010;
    x_250 = 'b111110110;
    x_251 = 'b111111010;
    x_252 = 'b000001110;
    x_253 = 'b000001010;
    x_254 = 'b111110111;
    x_255 = 'b000010010;

    h_0 = 'b111110001;
    h_1 = 'b111111011;
    h_2 = 'b111111000;
    h_3 = 'b000000111;
    h_4 = 'b000000110;
    h_5 = 'b000000001;
    h_6 = 'b111110101;
    h_7 = 'b000001011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111110101;
    x_1 = 'b111111011;
    x_2 = 'b111110100;
    x_3 = 'b111111111;
    x_4 = 'b111111101;
    x_5 = 'b111111001;
    x_6 = 'b111101110;
    x_7 = 'b000000100;
    x_8 = 'b111111111;
    x_9 = 'b111111001;
    x_10 = 'b111110111;
    x_11 = 'b111111101;
    x_12 = 'b111110001;
    x_13 = 'b111101001;
    x_14 = 'b111110100;
    x_15 = 'b111111000;
    x_16 = 'b111110101;
    x_17 = 'b111110101;
    x_18 = 'b111101011;
    x_19 = 'b111101001;
    x_20 = 'b111101010;
    x_21 = 'b111011110;
    x_22 = 'b111011111;
    x_23 = 'b111100000;
    x_24 = 'b111011011;
    x_25 = 'b111011100;
    x_26 = 'b111101010;
    x_27 = 'b111101001;
    x_28 = 'b111100000;
    x_29 = 'b111011001;
    x_30 = 'b111111101;
    x_31 = 'b111101000;
    x_32 = 'b111101000;
    x_33 = 'b111101001;
    x_34 = 'b111110011;
    x_35 = 'b111110000;
    x_36 = 'b111101001;
    x_37 = 'b111101011;
    x_38 = 'b111100100;
    x_39 = 'b111011110;
    x_40 = 'b111100100;
    x_41 = 'b111101100;
    x_42 = 'b111001011;
    x_43 = 'b111011101;
    x_44 = 'b111101001;
    x_45 = 'b111001100;
    x_46 = 'b111110010;
    x_47 = 'b111101110;
    x_48 = 'b111110000;
    x_49 = 'b111100111;
    x_50 = 'b111100011;
    x_51 = 'b111100000;
    x_52 = 'b111011001;
    x_53 = 'b111011111;
    x_54 = 'b111011100;
    x_55 = 'b111111001;
    x_56 = 'b111110110;
    x_57 = 'b111101110;
    x_58 = 'b111100011;
    x_59 = 'b111100101;
    x_60 = 'b000000111;
    x_61 = 'b111111111;
    x_62 = 'b111100110;
    x_63 = 'b000000110;
    x_64 = 'b111110101;
    x_65 = 'b111111011;
    x_66 = 'b111110100;
    x_67 = 'b111111111;
    x_68 = 'b111111101;
    x_69 = 'b111111001;
    x_70 = 'b111101110;
    x_71 = 'b000000100;
    x_72 = 'b111111111;
    x_73 = 'b111111001;
    x_74 = 'b111110111;
    x_75 = 'b111111101;
    x_76 = 'b111110001;
    x_77 = 'b111101001;
    x_78 = 'b111110100;
    x_79 = 'b111111000;
    x_80 = 'b111110101;
    x_81 = 'b111110101;
    x_82 = 'b111101011;
    x_83 = 'b111101001;
    x_84 = 'b111101010;
    x_85 = 'b111011110;
    x_86 = 'b111011111;
    x_87 = 'b111100000;
    x_88 = 'b111011011;
    x_89 = 'b111011100;
    x_90 = 'b111101010;
    x_91 = 'b111101001;
    x_92 = 'b111100000;
    x_93 = 'b111011001;
    x_94 = 'b111111101;
    x_95 = 'b111101000;
    x_96 = 'b111101000;
    x_97 = 'b111101001;
    x_98 = 'b111110011;
    x_99 = 'b111110000;
    x_100 = 'b111101001;
    x_101 = 'b111101011;
    x_102 = 'b111100100;
    x_103 = 'b111011110;
    x_104 = 'b111100100;
    x_105 = 'b111101100;
    x_106 = 'b111001011;
    x_107 = 'b111011101;
    x_108 = 'b111101001;
    x_109 = 'b111001100;
    x_110 = 'b111110010;
    x_111 = 'b111101110;
    x_112 = 'b111110000;
    x_113 = 'b111100111;
    x_114 = 'b111100011;
    x_115 = 'b111100000;
    x_116 = 'b111011001;
    x_117 = 'b111011111;
    x_118 = 'b111011100;
    x_119 = 'b111111001;
    x_120 = 'b111110110;
    x_121 = 'b111101110;
    x_122 = 'b111100011;
    x_123 = 'b111100101;
    x_124 = 'b000000111;
    x_125 = 'b111111111;
    x_126 = 'b111100110;
    x_127 = 'b000000110;
    x_128 = 'b111110101;
    x_129 = 'b111111011;
    x_130 = 'b111110100;
    x_131 = 'b111111111;
    x_132 = 'b111111101;
    x_133 = 'b111111001;
    x_134 = 'b111101110;
    x_135 = 'b000000100;
    x_136 = 'b111111111;
    x_137 = 'b111111001;
    x_138 = 'b111110111;
    x_139 = 'b111111101;
    x_140 = 'b111110001;
    x_141 = 'b111101001;
    x_142 = 'b111110100;
    x_143 = 'b111111000;
    x_144 = 'b111110101;
    x_145 = 'b111110101;
    x_146 = 'b111101011;
    x_147 = 'b111101001;
    x_148 = 'b111101010;
    x_149 = 'b111011110;
    x_150 = 'b111011111;
    x_151 = 'b111100000;
    x_152 = 'b111011011;
    x_153 = 'b111011100;
    x_154 = 'b111101010;
    x_155 = 'b111101001;
    x_156 = 'b111100000;
    x_157 = 'b111011001;
    x_158 = 'b111111101;
    x_159 = 'b111101000;
    x_160 = 'b111101000;
    x_161 = 'b111101001;
    x_162 = 'b111110011;
    x_163 = 'b111110000;
    x_164 = 'b111101001;
    x_165 = 'b111101011;
    x_166 = 'b111100100;
    x_167 = 'b111011110;
    x_168 = 'b111100100;
    x_169 = 'b111101100;
    x_170 = 'b111001011;
    x_171 = 'b111011101;
    x_172 = 'b111101001;
    x_173 = 'b111001100;
    x_174 = 'b111110010;
    x_175 = 'b111101110;
    x_176 = 'b111110000;
    x_177 = 'b111100111;
    x_178 = 'b111100011;
    x_179 = 'b111100000;
    x_180 = 'b111011001;
    x_181 = 'b111011111;
    x_182 = 'b111011100;
    x_183 = 'b111111001;
    x_184 = 'b111110110;
    x_185 = 'b111101110;
    x_186 = 'b111100011;
    x_187 = 'b111100101;
    x_188 = 'b000000111;
    x_189 = 'b111111111;
    x_190 = 'b111100110;
    x_191 = 'b000000110;
    x_192 = 'b111110101;
    x_193 = 'b111111011;
    x_194 = 'b111110100;
    x_195 = 'b111111111;
    x_196 = 'b111111101;
    x_197 = 'b111111001;
    x_198 = 'b111101110;
    x_199 = 'b000000100;
    x_200 = 'b111111111;
    x_201 = 'b111111001;
    x_202 = 'b111110111;
    x_203 = 'b111111101;
    x_204 = 'b111110001;
    x_205 = 'b111101001;
    x_206 = 'b111110100;
    x_207 = 'b111111000;
    x_208 = 'b111110101;
    x_209 = 'b111110101;
    x_210 = 'b111101011;
    x_211 = 'b111101001;
    x_212 = 'b111101010;
    x_213 = 'b111011110;
    x_214 = 'b111011111;
    x_215 = 'b111100000;
    x_216 = 'b111011011;
    x_217 = 'b111011100;
    x_218 = 'b111101010;
    x_219 = 'b111101001;
    x_220 = 'b111100000;
    x_221 = 'b111011001;
    x_222 = 'b111111101;
    x_223 = 'b111101000;
    x_224 = 'b111101000;
    x_225 = 'b111101001;
    x_226 = 'b111110011;
    x_227 = 'b111110000;
    x_228 = 'b111101001;
    x_229 = 'b111101011;
    x_230 = 'b111100100;
    x_231 = 'b111011110;
    x_232 = 'b111100100;
    x_233 = 'b111101100;
    x_234 = 'b111001011;
    x_235 = 'b111011101;
    x_236 = 'b111101001;
    x_237 = 'b111001100;
    x_238 = 'b111110010;
    x_239 = 'b111101110;
    x_240 = 'b111110000;
    x_241 = 'b111100111;
    x_242 = 'b111100011;
    x_243 = 'b111100000;
    x_244 = 'b111011001;
    x_245 = 'b111011111;
    x_246 = 'b111011100;
    x_247 = 'b111111001;
    x_248 = 'b111110110;
    x_249 = 'b111101110;
    x_250 = 'b111100011;
    x_251 = 'b111100101;
    x_252 = 'b000000111;
    x_253 = 'b111111111;
    x_254 = 'b111100110;
    x_255 = 'b000000110;

    h_0 = 'b111110101;
    h_1 = 'b111111011;
    h_2 = 'b111110100;
    h_3 = 'b111111111;
    h_4 = 'b111111101;
    h_5 = 'b111111001;
    h_6 = 'b111101110;
    h_7 = 'b000000100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111101001;
    x_1 = 'b111110010;
    x_2 = 'b111101101;
    x_3 = 'b111110100;
    x_4 = 'b111110101;
    x_5 = 'b111110011;
    x_6 = 'b111101110;
    x_7 = 'b111110000;
    x_8 = 'b111110001;
    x_9 = 'b111101111;
    x_10 = 'b111101101;
    x_11 = 'b111110111;
    x_12 = 'b111101100;
    x_13 = 'b111101001;
    x_14 = 'b111100111;
    x_15 = 'b111101001;
    x_16 = 'b111101010;
    x_17 = 'b111101011;
    x_18 = 'b111100111;
    x_19 = 'b111100111;
    x_20 = 'b111101001;
    x_21 = 'b111011111;
    x_22 = 'b111100000;
    x_23 = 'b111100001;
    x_24 = 'b111011110;
    x_25 = 'b111011101;
    x_26 = 'b111101111;
    x_27 = 'b111101100;
    x_28 = 'b111100000;
    x_29 = 'b111100000;
    x_30 = 'b111111010;
    x_31 = 'b111101011;
    x_32 = 'b111110000;
    x_33 = 'b111110010;
    x_34 = 'b111111001;
    x_35 = 'b111110110;
    x_36 = 'b111101111;
    x_37 = 'b111110001;
    x_38 = 'b111101011;
    x_39 = 'b111110100;
    x_40 = 'b111110011;
    x_41 = 'b000001100;
    x_42 = 'b111010010;
    x_43 = 'b111010000;
    x_44 = 'b111101011;
    x_45 = 'b111011001;
    x_46 = 'b111110101;
    x_47 = 'b111101110;
    x_48 = 'b111110001;
    x_49 = 'b111101100;
    x_50 = 'b111101011;
    x_51 = 'b111110000;
    x_52 = 'b111101001;
    x_53 = 'b111101110;
    x_54 = 'b111101011;
    x_55 = 'b111111100;
    x_56 = 'b111111001;
    x_57 = 'b111111001;
    x_58 = 'b111110110;
    x_59 = 'b111110110;
    x_60 = 'b111111111;
    x_61 = 'b111110111;
    x_62 = 'b111011111;
    x_63 = 'b111111011;
    x_64 = 'b111101001;
    x_65 = 'b111110010;
    x_66 = 'b111101101;
    x_67 = 'b111110100;
    x_68 = 'b111110101;
    x_69 = 'b111110011;
    x_70 = 'b111101110;
    x_71 = 'b111110000;
    x_72 = 'b111110001;
    x_73 = 'b111101111;
    x_74 = 'b111101101;
    x_75 = 'b111110111;
    x_76 = 'b111101100;
    x_77 = 'b111101001;
    x_78 = 'b111100111;
    x_79 = 'b111101001;
    x_80 = 'b111101010;
    x_81 = 'b111101011;
    x_82 = 'b111100111;
    x_83 = 'b111100111;
    x_84 = 'b111101001;
    x_85 = 'b111011111;
    x_86 = 'b111100000;
    x_87 = 'b111100001;
    x_88 = 'b111011110;
    x_89 = 'b111011101;
    x_90 = 'b111101111;
    x_91 = 'b111101100;
    x_92 = 'b111100000;
    x_93 = 'b111100000;
    x_94 = 'b111111010;
    x_95 = 'b111101011;
    x_96 = 'b111110000;
    x_97 = 'b111110010;
    x_98 = 'b111111001;
    x_99 = 'b111110110;
    x_100 = 'b111101111;
    x_101 = 'b111110001;
    x_102 = 'b111101011;
    x_103 = 'b111110100;
    x_104 = 'b111110011;
    x_105 = 'b000001100;
    x_106 = 'b111010010;
    x_107 = 'b111010000;
    x_108 = 'b111101011;
    x_109 = 'b111011001;
    x_110 = 'b111110101;
    x_111 = 'b111101110;
    x_112 = 'b111110001;
    x_113 = 'b111101100;
    x_114 = 'b111101011;
    x_115 = 'b111110000;
    x_116 = 'b111101001;
    x_117 = 'b111101110;
    x_118 = 'b111101011;
    x_119 = 'b111111100;
    x_120 = 'b111111001;
    x_121 = 'b111111001;
    x_122 = 'b111110110;
    x_123 = 'b111110110;
    x_124 = 'b111111111;
    x_125 = 'b111110111;
    x_126 = 'b111011111;
    x_127 = 'b111111011;
    x_128 = 'b111101001;
    x_129 = 'b111110010;
    x_130 = 'b111101101;
    x_131 = 'b111110100;
    x_132 = 'b111110101;
    x_133 = 'b111110011;
    x_134 = 'b111101110;
    x_135 = 'b111110000;
    x_136 = 'b111110001;
    x_137 = 'b111101111;
    x_138 = 'b111101101;
    x_139 = 'b111110111;
    x_140 = 'b111101100;
    x_141 = 'b111101001;
    x_142 = 'b111100111;
    x_143 = 'b111101001;
    x_144 = 'b111101010;
    x_145 = 'b111101011;
    x_146 = 'b111100111;
    x_147 = 'b111100111;
    x_148 = 'b111101001;
    x_149 = 'b111011111;
    x_150 = 'b111100000;
    x_151 = 'b111100001;
    x_152 = 'b111011110;
    x_153 = 'b111011101;
    x_154 = 'b111101111;
    x_155 = 'b111101100;
    x_156 = 'b111100000;
    x_157 = 'b111100000;
    x_158 = 'b111111010;
    x_159 = 'b111101011;
    x_160 = 'b111110000;
    x_161 = 'b111110010;
    x_162 = 'b111111001;
    x_163 = 'b111110110;
    x_164 = 'b111101111;
    x_165 = 'b111110001;
    x_166 = 'b111101011;
    x_167 = 'b111110100;
    x_168 = 'b111110011;
    x_169 = 'b000001100;
    x_170 = 'b111010010;
    x_171 = 'b111010000;
    x_172 = 'b111101011;
    x_173 = 'b111011001;
    x_174 = 'b111110101;
    x_175 = 'b111101110;
    x_176 = 'b111110001;
    x_177 = 'b111101100;
    x_178 = 'b111101011;
    x_179 = 'b111110000;
    x_180 = 'b111101001;
    x_181 = 'b111101110;
    x_182 = 'b111101011;
    x_183 = 'b111111100;
    x_184 = 'b111111001;
    x_185 = 'b111111001;
    x_186 = 'b111110110;
    x_187 = 'b111110110;
    x_188 = 'b111111111;
    x_189 = 'b111110111;
    x_190 = 'b111011111;
    x_191 = 'b111111011;
    x_192 = 'b111101001;
    x_193 = 'b111110010;
    x_194 = 'b111101101;
    x_195 = 'b111110100;
    x_196 = 'b111110101;
    x_197 = 'b111110011;
    x_198 = 'b111101110;
    x_199 = 'b111110000;
    x_200 = 'b111110001;
    x_201 = 'b111101111;
    x_202 = 'b111101101;
    x_203 = 'b111110111;
    x_204 = 'b111101100;
    x_205 = 'b111101001;
    x_206 = 'b111100111;
    x_207 = 'b111101001;
    x_208 = 'b111101010;
    x_209 = 'b111101011;
    x_210 = 'b111100111;
    x_211 = 'b111100111;
    x_212 = 'b111101001;
    x_213 = 'b111011111;
    x_214 = 'b111100000;
    x_215 = 'b111100001;
    x_216 = 'b111011110;
    x_217 = 'b111011101;
    x_218 = 'b111101111;
    x_219 = 'b111101100;
    x_220 = 'b111100000;
    x_221 = 'b111100000;
    x_222 = 'b111111010;
    x_223 = 'b111101011;
    x_224 = 'b111110000;
    x_225 = 'b111110010;
    x_226 = 'b111111001;
    x_227 = 'b111110110;
    x_228 = 'b111101111;
    x_229 = 'b111110001;
    x_230 = 'b111101011;
    x_231 = 'b111110100;
    x_232 = 'b111110011;
    x_233 = 'b000001100;
    x_234 = 'b111010010;
    x_235 = 'b111010000;
    x_236 = 'b111101011;
    x_237 = 'b111011001;
    x_238 = 'b111110101;
    x_239 = 'b111101110;
    x_240 = 'b111110001;
    x_241 = 'b111101100;
    x_242 = 'b111101011;
    x_243 = 'b111110000;
    x_244 = 'b111101001;
    x_245 = 'b111101110;
    x_246 = 'b111101011;
    x_247 = 'b111111100;
    x_248 = 'b111111001;
    x_249 = 'b111111001;
    x_250 = 'b111110110;
    x_251 = 'b111110110;
    x_252 = 'b111111111;
    x_253 = 'b111110111;
    x_254 = 'b111011111;
    x_255 = 'b111111011;

    h_0 = 'b111101001;
    h_1 = 'b111110010;
    h_2 = 'b111101101;
    h_3 = 'b111110100;
    h_4 = 'b111110101;
    h_5 = 'b111110011;
    h_6 = 'b111101110;
    h_7 = 'b111110000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111101011;
    x_1 = 'b111110110;
    x_2 = 'b111110100;
    x_3 = 'b111111101;
    x_4 = 'b111111111;
    x_5 = 'b000000000;
    x_6 = 'b111110101;
    x_7 = 'b111111000;
    x_8 = 'b111110101;
    x_9 = 'b111110100;
    x_10 = 'b111110101;
    x_11 = 'b000000001;
    x_12 = 'b111111011;
    x_13 = 'b111111000;
    x_14 = 'b111101011;
    x_15 = 'b111101101;
    x_16 = 'b111110010;
    x_17 = 'b111110010;
    x_18 = 'b111110101;
    x_19 = 'b111111000;
    x_20 = 'b111111000;
    x_21 = 'b111100000;
    x_22 = 'b111011110;
    x_23 = 'b111100000;
    x_24 = 'b111011110;
    x_25 = 'b111011111;
    x_26 = 'b111101101;
    x_27 = 'b111101010;
    x_28 = 'b111011111;
    x_29 = 'b111100011;
    x_30 = 'b111110101;
    x_31 = 'b111101110;
    x_32 = 'b111101111;
    x_33 = 'b111110011;
    x_34 = 'b111111001;
    x_35 = 'b111110100;
    x_36 = 'b111101110;
    x_37 = 'b111110001;
    x_38 = 'b111101100;
    x_39 = 'b111110111;
    x_40 = 'b111011010;
    x_41 = 'b111111010;
    x_42 = 'b111001111;
    x_43 = 'b111110111;
    x_44 = 'b111101001;
    x_45 = 'b111101101;
    x_46 = 'b111110001;
    x_47 = 'b111101110;
    x_48 = 'b111110001;
    x_49 = 'b111110011;
    x_50 = 'b111110101;
    x_51 = 'b111111110;
    x_52 = 'b111111010;
    x_53 = 'b111111110;
    x_54 = 'b111111011;
    x_55 = 'b111111000;
    x_56 = 'b111110101;
    x_57 = 'b000000001;
    x_58 = 'b000000100;
    x_59 = 'b000000100;
    x_60 = 'b111111100;
    x_61 = 'b111111010;
    x_62 = 'b111101011;
    x_63 = 'b111111110;
    x_64 = 'b111101011;
    x_65 = 'b111110110;
    x_66 = 'b111110100;
    x_67 = 'b111111101;
    x_68 = 'b111111111;
    x_69 = 'b000000000;
    x_70 = 'b111110101;
    x_71 = 'b111111000;
    x_72 = 'b111110101;
    x_73 = 'b111110100;
    x_74 = 'b111110101;
    x_75 = 'b000000001;
    x_76 = 'b111111011;
    x_77 = 'b111111000;
    x_78 = 'b111101011;
    x_79 = 'b111101101;
    x_80 = 'b111110010;
    x_81 = 'b111110010;
    x_82 = 'b111110101;
    x_83 = 'b111111000;
    x_84 = 'b111111000;
    x_85 = 'b111100000;
    x_86 = 'b111011110;
    x_87 = 'b111100000;
    x_88 = 'b111011110;
    x_89 = 'b111011111;
    x_90 = 'b111101101;
    x_91 = 'b111101010;
    x_92 = 'b111011111;
    x_93 = 'b111100011;
    x_94 = 'b111110101;
    x_95 = 'b111101110;
    x_96 = 'b111101111;
    x_97 = 'b111110011;
    x_98 = 'b111111001;
    x_99 = 'b111110100;
    x_100 = 'b111101110;
    x_101 = 'b111110001;
    x_102 = 'b111101100;
    x_103 = 'b111110111;
    x_104 = 'b111011010;
    x_105 = 'b111111010;
    x_106 = 'b111001111;
    x_107 = 'b111110111;
    x_108 = 'b111101001;
    x_109 = 'b111101101;
    x_110 = 'b111110001;
    x_111 = 'b111101110;
    x_112 = 'b111110001;
    x_113 = 'b111110011;
    x_114 = 'b111110101;
    x_115 = 'b111111110;
    x_116 = 'b111111010;
    x_117 = 'b111111110;
    x_118 = 'b111111011;
    x_119 = 'b111111000;
    x_120 = 'b111110101;
    x_121 = 'b000000001;
    x_122 = 'b000000100;
    x_123 = 'b000000100;
    x_124 = 'b111111100;
    x_125 = 'b111111010;
    x_126 = 'b111101011;
    x_127 = 'b111111110;
    x_128 = 'b111101011;
    x_129 = 'b111110110;
    x_130 = 'b111110100;
    x_131 = 'b111111101;
    x_132 = 'b111111111;
    x_133 = 'b000000000;
    x_134 = 'b111110101;
    x_135 = 'b111111000;
    x_136 = 'b111110101;
    x_137 = 'b111110100;
    x_138 = 'b111110101;
    x_139 = 'b000000001;
    x_140 = 'b111111011;
    x_141 = 'b111111000;
    x_142 = 'b111101011;
    x_143 = 'b111101101;
    x_144 = 'b111110010;
    x_145 = 'b111110010;
    x_146 = 'b111110101;
    x_147 = 'b111111000;
    x_148 = 'b111111000;
    x_149 = 'b111100000;
    x_150 = 'b111011110;
    x_151 = 'b111100000;
    x_152 = 'b111011110;
    x_153 = 'b111011111;
    x_154 = 'b111101101;
    x_155 = 'b111101010;
    x_156 = 'b111011111;
    x_157 = 'b111100011;
    x_158 = 'b111110101;
    x_159 = 'b111101110;
    x_160 = 'b111101111;
    x_161 = 'b111110011;
    x_162 = 'b111111001;
    x_163 = 'b111110100;
    x_164 = 'b111101110;
    x_165 = 'b111110001;
    x_166 = 'b111101100;
    x_167 = 'b111110111;
    x_168 = 'b111011010;
    x_169 = 'b111111010;
    x_170 = 'b111001111;
    x_171 = 'b111110111;
    x_172 = 'b111101001;
    x_173 = 'b111101101;
    x_174 = 'b111110001;
    x_175 = 'b111101110;
    x_176 = 'b111110001;
    x_177 = 'b111110011;
    x_178 = 'b111110101;
    x_179 = 'b111111110;
    x_180 = 'b111111010;
    x_181 = 'b111111110;
    x_182 = 'b111111011;
    x_183 = 'b111111000;
    x_184 = 'b111110101;
    x_185 = 'b000000001;
    x_186 = 'b000000100;
    x_187 = 'b000000100;
    x_188 = 'b111111100;
    x_189 = 'b111111010;
    x_190 = 'b111101011;
    x_191 = 'b111111110;
    x_192 = 'b111101011;
    x_193 = 'b111110110;
    x_194 = 'b111110100;
    x_195 = 'b111111101;
    x_196 = 'b111111111;
    x_197 = 'b000000000;
    x_198 = 'b111110101;
    x_199 = 'b111111000;
    x_200 = 'b111110101;
    x_201 = 'b111110100;
    x_202 = 'b111110101;
    x_203 = 'b000000001;
    x_204 = 'b111111011;
    x_205 = 'b111111000;
    x_206 = 'b111101011;
    x_207 = 'b111101101;
    x_208 = 'b111110010;
    x_209 = 'b111110010;
    x_210 = 'b111110101;
    x_211 = 'b111111000;
    x_212 = 'b111111000;
    x_213 = 'b111100000;
    x_214 = 'b111011110;
    x_215 = 'b111100000;
    x_216 = 'b111011110;
    x_217 = 'b111011111;
    x_218 = 'b111101101;
    x_219 = 'b111101010;
    x_220 = 'b111011111;
    x_221 = 'b111100011;
    x_222 = 'b111110101;
    x_223 = 'b111101110;
    x_224 = 'b111101111;
    x_225 = 'b111110011;
    x_226 = 'b111111001;
    x_227 = 'b111110100;
    x_228 = 'b111101110;
    x_229 = 'b111110001;
    x_230 = 'b111101100;
    x_231 = 'b111110111;
    x_232 = 'b111011010;
    x_233 = 'b111111010;
    x_234 = 'b111001111;
    x_235 = 'b111110111;
    x_236 = 'b111101001;
    x_237 = 'b111101101;
    x_238 = 'b111110001;
    x_239 = 'b111101110;
    x_240 = 'b111110001;
    x_241 = 'b111110011;
    x_242 = 'b111110101;
    x_243 = 'b111111110;
    x_244 = 'b111111010;
    x_245 = 'b111111110;
    x_246 = 'b111111011;
    x_247 = 'b111111000;
    x_248 = 'b111110101;
    x_249 = 'b000000001;
    x_250 = 'b000000100;
    x_251 = 'b000000100;
    x_252 = 'b111111100;
    x_253 = 'b111111010;
    x_254 = 'b111101011;
    x_255 = 'b111111110;

    h_0 = 'b111101011;
    h_1 = 'b111110110;
    h_2 = 'b111110100;
    h_3 = 'b111111101;
    h_4 = 'b111111111;
    h_5 = 'b000000000;
    h_6 = 'b111110101;
    h_7 = 'b111111000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000001110;
    x_1 = 'b000001110;
    x_2 = 'b000000110;
    x_3 = 'b000001100;
    x_4 = 'b000010000;
    x_5 = 'b000000111;
    x_6 = 'b000000111;
    x_7 = 'b000000011;
    x_8 = 'b000001010;
    x_9 = 'b000001100;
    x_10 = 'b000010001;
    x_11 = 'b000000010;
    x_12 = 'b000001011;
    x_13 = 'b000010000;
    x_14 = 'b000001011;
    x_15 = 'b000001100;
    x_16 = 'b000001101;
    x_17 = 'b000001011;
    x_18 = 'b000001011;
    x_19 = 'b000010000;
    x_20 = 'b000001000;
    x_21 = 'b000000100;
    x_22 = 'b000000110;
    x_23 = 'b111111100;
    x_24 = 'b111111011;
    x_25 = 'b111111100;
    x_26 = 'b111111100;
    x_27 = 'b111111101;
    x_28 = 'b000000100;
    x_29 = 'b000000110;
    x_30 = 'b111111100;
    x_31 = 'b111110110;
    x_32 = 'b111111101;
    x_33 = 'b111111011;
    x_34 = 'b111111000;
    x_35 = 'b111111011;
    x_36 = 'b111111011;
    x_37 = 'b000001000;
    x_38 = 'b111111100;
    x_39 = 'b000001100;
    x_40 = 'b111111111;
    x_41 = 'b111110000;
    x_42 = 'b111111011;
    x_43 = 'b000011110;
    x_44 = 'b111110001;
    x_45 = 'b000010101;
    x_46 = 'b000001000;
    x_47 = 'b000000111;
    x_48 = 'b000001001;
    x_49 = 'b000001000;
    x_50 = 'b000001101;
    x_51 = 'b000001111;
    x_52 = 'b000001101;
    x_53 = 'b000001011;
    x_54 = 'b000000111;
    x_55 = 'b000001010;
    x_56 = 'b000000111;
    x_57 = 'b000010010;
    x_58 = 'b000010101;
    x_59 = 'b000010111;
    x_60 = 'b000010111;
    x_61 = 'b000100101;
    x_62 = 'b000010010;
    x_63 = 'b000001111;
    x_64 = 'b000001110;
    x_65 = 'b000001110;
    x_66 = 'b000000110;
    x_67 = 'b000001100;
    x_68 = 'b000010000;
    x_69 = 'b000000111;
    x_70 = 'b000000111;
    x_71 = 'b000000011;
    x_72 = 'b000001010;
    x_73 = 'b000001100;
    x_74 = 'b000010001;
    x_75 = 'b000000010;
    x_76 = 'b000001011;
    x_77 = 'b000010000;
    x_78 = 'b000001011;
    x_79 = 'b000001100;
    x_80 = 'b000001101;
    x_81 = 'b000001011;
    x_82 = 'b000001011;
    x_83 = 'b000010000;
    x_84 = 'b000001000;
    x_85 = 'b000000100;
    x_86 = 'b000000110;
    x_87 = 'b111111100;
    x_88 = 'b111111011;
    x_89 = 'b111111100;
    x_90 = 'b111111100;
    x_91 = 'b111111101;
    x_92 = 'b000000100;
    x_93 = 'b000000110;
    x_94 = 'b111111100;
    x_95 = 'b111110110;
    x_96 = 'b111111101;
    x_97 = 'b111111011;
    x_98 = 'b111111000;
    x_99 = 'b111111011;
    x_100 = 'b111111011;
    x_101 = 'b000001000;
    x_102 = 'b111111100;
    x_103 = 'b000001100;
    x_104 = 'b111111111;
    x_105 = 'b111110000;
    x_106 = 'b111111011;
    x_107 = 'b000011110;
    x_108 = 'b111110001;
    x_109 = 'b000010101;
    x_110 = 'b000001000;
    x_111 = 'b000000111;
    x_112 = 'b000001001;
    x_113 = 'b000001000;
    x_114 = 'b000001101;
    x_115 = 'b000001111;
    x_116 = 'b000001101;
    x_117 = 'b000001011;
    x_118 = 'b000000111;
    x_119 = 'b000001010;
    x_120 = 'b000000111;
    x_121 = 'b000010010;
    x_122 = 'b000010101;
    x_123 = 'b000010111;
    x_124 = 'b000010111;
    x_125 = 'b000100101;
    x_126 = 'b000010010;
    x_127 = 'b000001111;
    x_128 = 'b000001110;
    x_129 = 'b000001110;
    x_130 = 'b000000110;
    x_131 = 'b000001100;
    x_132 = 'b000010000;
    x_133 = 'b000000111;
    x_134 = 'b000000111;
    x_135 = 'b000000011;
    x_136 = 'b000001010;
    x_137 = 'b000001100;
    x_138 = 'b000010001;
    x_139 = 'b000000010;
    x_140 = 'b000001011;
    x_141 = 'b000010000;
    x_142 = 'b000001011;
    x_143 = 'b000001100;
    x_144 = 'b000001101;
    x_145 = 'b000001011;
    x_146 = 'b000001011;
    x_147 = 'b000010000;
    x_148 = 'b000001000;
    x_149 = 'b000000100;
    x_150 = 'b000000110;
    x_151 = 'b111111100;
    x_152 = 'b111111011;
    x_153 = 'b111111100;
    x_154 = 'b111111100;
    x_155 = 'b111111101;
    x_156 = 'b000000100;
    x_157 = 'b000000110;
    x_158 = 'b111111100;
    x_159 = 'b111110110;
    x_160 = 'b111111101;
    x_161 = 'b111111011;
    x_162 = 'b111111000;
    x_163 = 'b111111011;
    x_164 = 'b111111011;
    x_165 = 'b000001000;
    x_166 = 'b111111100;
    x_167 = 'b000001100;
    x_168 = 'b111111111;
    x_169 = 'b111110000;
    x_170 = 'b111111011;
    x_171 = 'b000011110;
    x_172 = 'b111110001;
    x_173 = 'b000010101;
    x_174 = 'b000001000;
    x_175 = 'b000000111;
    x_176 = 'b000001001;
    x_177 = 'b000001000;
    x_178 = 'b000001101;
    x_179 = 'b000001111;
    x_180 = 'b000001101;
    x_181 = 'b000001011;
    x_182 = 'b000000111;
    x_183 = 'b000001010;
    x_184 = 'b000000111;
    x_185 = 'b000010010;
    x_186 = 'b000010101;
    x_187 = 'b000010111;
    x_188 = 'b000010111;
    x_189 = 'b000100101;
    x_190 = 'b000010010;
    x_191 = 'b000001111;
    x_192 = 'b000001110;
    x_193 = 'b000001110;
    x_194 = 'b000000110;
    x_195 = 'b000001100;
    x_196 = 'b000010000;
    x_197 = 'b000000111;
    x_198 = 'b000000111;
    x_199 = 'b000000011;
    x_200 = 'b000001010;
    x_201 = 'b000001100;
    x_202 = 'b000010001;
    x_203 = 'b000000010;
    x_204 = 'b000001011;
    x_205 = 'b000010000;
    x_206 = 'b000001011;
    x_207 = 'b000001100;
    x_208 = 'b000001101;
    x_209 = 'b000001011;
    x_210 = 'b000001011;
    x_211 = 'b000010000;
    x_212 = 'b000001000;
    x_213 = 'b000000100;
    x_214 = 'b000000110;
    x_215 = 'b111111100;
    x_216 = 'b111111011;
    x_217 = 'b111111100;
    x_218 = 'b111111100;
    x_219 = 'b111111101;
    x_220 = 'b000000100;
    x_221 = 'b000000110;
    x_222 = 'b111111100;
    x_223 = 'b111110110;
    x_224 = 'b111111101;
    x_225 = 'b111111011;
    x_226 = 'b111111000;
    x_227 = 'b111111011;
    x_228 = 'b111111011;
    x_229 = 'b000001000;
    x_230 = 'b111111100;
    x_231 = 'b000001100;
    x_232 = 'b111111111;
    x_233 = 'b111110000;
    x_234 = 'b111111011;
    x_235 = 'b000011110;
    x_236 = 'b111110001;
    x_237 = 'b000010101;
    x_238 = 'b000001000;
    x_239 = 'b000000111;
    x_240 = 'b000001001;
    x_241 = 'b000001000;
    x_242 = 'b000001101;
    x_243 = 'b000001111;
    x_244 = 'b000001101;
    x_245 = 'b000001011;
    x_246 = 'b000000111;
    x_247 = 'b000001010;
    x_248 = 'b000000111;
    x_249 = 'b000010010;
    x_250 = 'b000010101;
    x_251 = 'b000010111;
    x_252 = 'b000010111;
    x_253 = 'b000100101;
    x_254 = 'b000010010;
    x_255 = 'b000001111;

    h_0 = 'b000001110;
    h_1 = 'b000001110;
    h_2 = 'b000000110;
    h_3 = 'b000001100;
    h_4 = 'b000010000;
    h_5 = 'b000000111;
    h_6 = 'b000000111;
    h_7 = 'b000000011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000000101;
    x_1 = 'b000000110;
    x_2 = 'b000000001;
    x_3 = 'b000001010;
    x_4 = 'b000001101;
    x_5 = 'b000000000;
    x_6 = 'b111111110;
    x_7 = 'b111111011;
    x_8 = 'b000000011;
    x_9 = 'b000001001;
    x_10 = 'b000001101;
    x_11 = 'b000000011;
    x_12 = 'b000000110;
    x_13 = 'b000000111;
    x_14 = 'b000000110;
    x_15 = 'b000000100;
    x_16 = 'b000000110;
    x_17 = 'b000000110;
    x_18 = 'b000001000;
    x_19 = 'b000001011;
    x_20 = 'b000000010;
    x_21 = 'b000000111;
    x_22 = 'b000001001;
    x_23 = 'b000000000;
    x_24 = 'b111111100;
    x_25 = 'b111111101;
    x_26 = 'b000000000;
    x_27 = 'b000000001;
    x_28 = 'b000000110;
    x_29 = 'b000000011;
    x_30 = 'b111111100;
    x_31 = 'b111111000;
    x_32 = 'b000000001;
    x_33 = 'b000000001;
    x_34 = 'b111111101;
    x_35 = 'b111111101;
    x_36 = 'b111111000;
    x_37 = 'b000000110;
    x_38 = 'b111111001;
    x_39 = 'b000000000;
    x_40 = 'b000000000;
    x_41 = 'b111011010;
    x_42 = 'b111101101;
    x_43 = 'b000010000;
    x_44 = 'b111101100;
    x_45 = 'b000100001;
    x_46 = 'b000000011;
    x_47 = 'b000000011;
    x_48 = 'b000000111;
    x_49 = 'b000001000;
    x_50 = 'b000001011;
    x_51 = 'b000001111;
    x_52 = 'b000001100;
    x_53 = 'b000001100;
    x_54 = 'b000001101;
    x_55 = 'b000001001;
    x_56 = 'b000000110;
    x_57 = 'b000010001;
    x_58 = 'b000010010;
    x_59 = 'b000011000;
    x_60 = 'b000010111;
    x_61 = 'b000100000;
    x_62 = 'b000001010;
    x_63 = 'b000010010;
    x_64 = 'b000000101;
    x_65 = 'b000000110;
    x_66 = 'b000000001;
    x_67 = 'b000001010;
    x_68 = 'b000001101;
    x_69 = 'b000000000;
    x_70 = 'b111111110;
    x_71 = 'b111111011;
    x_72 = 'b000000011;
    x_73 = 'b000001001;
    x_74 = 'b000001101;
    x_75 = 'b000000011;
    x_76 = 'b000000110;
    x_77 = 'b000000111;
    x_78 = 'b000000110;
    x_79 = 'b000000100;
    x_80 = 'b000000110;
    x_81 = 'b000000110;
    x_82 = 'b000001000;
    x_83 = 'b000001011;
    x_84 = 'b000000010;
    x_85 = 'b000000111;
    x_86 = 'b000001001;
    x_87 = 'b000000000;
    x_88 = 'b111111100;
    x_89 = 'b111111101;
    x_90 = 'b000000000;
    x_91 = 'b000000001;
    x_92 = 'b000000110;
    x_93 = 'b000000011;
    x_94 = 'b111111100;
    x_95 = 'b111111000;
    x_96 = 'b000000001;
    x_97 = 'b000000001;
    x_98 = 'b111111101;
    x_99 = 'b111111101;
    x_100 = 'b111111000;
    x_101 = 'b000000110;
    x_102 = 'b111111001;
    x_103 = 'b000000000;
    x_104 = 'b000000000;
    x_105 = 'b111011010;
    x_106 = 'b111101101;
    x_107 = 'b000010000;
    x_108 = 'b111101100;
    x_109 = 'b000100001;
    x_110 = 'b000000011;
    x_111 = 'b000000011;
    x_112 = 'b000000111;
    x_113 = 'b000001000;
    x_114 = 'b000001011;
    x_115 = 'b000001111;
    x_116 = 'b000001100;
    x_117 = 'b000001100;
    x_118 = 'b000001101;
    x_119 = 'b000001001;
    x_120 = 'b000000110;
    x_121 = 'b000010001;
    x_122 = 'b000010010;
    x_123 = 'b000011000;
    x_124 = 'b000010111;
    x_125 = 'b000100000;
    x_126 = 'b000001010;
    x_127 = 'b000010010;
    x_128 = 'b000000101;
    x_129 = 'b000000110;
    x_130 = 'b000000001;
    x_131 = 'b000001010;
    x_132 = 'b000001101;
    x_133 = 'b000000000;
    x_134 = 'b111111110;
    x_135 = 'b111111011;
    x_136 = 'b000000011;
    x_137 = 'b000001001;
    x_138 = 'b000001101;
    x_139 = 'b000000011;
    x_140 = 'b000000110;
    x_141 = 'b000000111;
    x_142 = 'b000000110;
    x_143 = 'b000000100;
    x_144 = 'b000000110;
    x_145 = 'b000000110;
    x_146 = 'b000001000;
    x_147 = 'b000001011;
    x_148 = 'b000000010;
    x_149 = 'b000000111;
    x_150 = 'b000001001;
    x_151 = 'b000000000;
    x_152 = 'b111111100;
    x_153 = 'b111111101;
    x_154 = 'b000000000;
    x_155 = 'b000000001;
    x_156 = 'b000000110;
    x_157 = 'b000000011;
    x_158 = 'b111111100;
    x_159 = 'b111111000;
    x_160 = 'b000000001;
    x_161 = 'b000000001;
    x_162 = 'b111111101;
    x_163 = 'b111111101;
    x_164 = 'b111111000;
    x_165 = 'b000000110;
    x_166 = 'b111111001;
    x_167 = 'b000000000;
    x_168 = 'b000000000;
    x_169 = 'b111011010;
    x_170 = 'b111101101;
    x_171 = 'b000010000;
    x_172 = 'b111101100;
    x_173 = 'b000100001;
    x_174 = 'b000000011;
    x_175 = 'b000000011;
    x_176 = 'b000000111;
    x_177 = 'b000001000;
    x_178 = 'b000001011;
    x_179 = 'b000001111;
    x_180 = 'b000001100;
    x_181 = 'b000001100;
    x_182 = 'b000001101;
    x_183 = 'b000001001;
    x_184 = 'b000000110;
    x_185 = 'b000010001;
    x_186 = 'b000010010;
    x_187 = 'b000011000;
    x_188 = 'b000010111;
    x_189 = 'b000100000;
    x_190 = 'b000001010;
    x_191 = 'b000010010;
    x_192 = 'b000000101;
    x_193 = 'b000000110;
    x_194 = 'b000000001;
    x_195 = 'b000001010;
    x_196 = 'b000001101;
    x_197 = 'b000000000;
    x_198 = 'b111111110;
    x_199 = 'b111111011;
    x_200 = 'b000000011;
    x_201 = 'b000001001;
    x_202 = 'b000001101;
    x_203 = 'b000000011;
    x_204 = 'b000000110;
    x_205 = 'b000000111;
    x_206 = 'b000000110;
    x_207 = 'b000000100;
    x_208 = 'b000000110;
    x_209 = 'b000000110;
    x_210 = 'b000001000;
    x_211 = 'b000001011;
    x_212 = 'b000000010;
    x_213 = 'b000000111;
    x_214 = 'b000001001;
    x_215 = 'b000000000;
    x_216 = 'b111111100;
    x_217 = 'b111111101;
    x_218 = 'b000000000;
    x_219 = 'b000000001;
    x_220 = 'b000000110;
    x_221 = 'b000000011;
    x_222 = 'b111111100;
    x_223 = 'b111111000;
    x_224 = 'b000000001;
    x_225 = 'b000000001;
    x_226 = 'b111111101;
    x_227 = 'b111111101;
    x_228 = 'b111111000;
    x_229 = 'b000000110;
    x_230 = 'b111111001;
    x_231 = 'b000000000;
    x_232 = 'b000000000;
    x_233 = 'b111011010;
    x_234 = 'b111101101;
    x_235 = 'b000010000;
    x_236 = 'b111101100;
    x_237 = 'b000100001;
    x_238 = 'b000000011;
    x_239 = 'b000000011;
    x_240 = 'b000000111;
    x_241 = 'b000001000;
    x_242 = 'b000001011;
    x_243 = 'b000001111;
    x_244 = 'b000001100;
    x_245 = 'b000001100;
    x_246 = 'b000001101;
    x_247 = 'b000001001;
    x_248 = 'b000000110;
    x_249 = 'b000010001;
    x_250 = 'b000010010;
    x_251 = 'b000011000;
    x_252 = 'b000010111;
    x_253 = 'b000100000;
    x_254 = 'b000001010;
    x_255 = 'b000010010;

    h_0 = 'b000000101;
    h_1 = 'b000000110;
    h_2 = 'b000000001;
    h_3 = 'b000001010;
    h_4 = 'b000001101;
    h_5 = 'b000000000;
    h_6 = 'b111111110;
    h_7 = 'b111111011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111111011;
    x_1 = 'b000000000;
    x_2 = 'b000000000;
    x_3 = 'b000001100;
    x_4 = 'b000001110;
    x_5 = 'b000000000;
    x_6 = 'b111111010;
    x_7 = 'b111101111;
    x_8 = 'b111111010;
    x_9 = 'b000000101;
    x_10 = 'b000001111;
    x_11 = 'b000000000;
    x_12 = 'b000000011;
    x_13 = 'b000000110;
    x_14 = 'b111110111;
    x_15 = 'b111111110;
    x_16 = 'b000000010;
    x_17 = 'b000000100;
    x_18 = 'b000000100;
    x_19 = 'b000000101;
    x_20 = 'b111111111;
    x_21 = 'b111111101;
    x_22 = 'b111111110;
    x_23 = 'b111111000;
    x_24 = 'b111101101;
    x_25 = 'b111101110;
    x_26 = 'b111110100;
    x_27 = 'b111110101;
    x_28 = 'b111111110;
    x_29 = 'b111110010;
    x_30 = 'b111101001;
    x_31 = 'b111101110;
    x_32 = 'b111110011;
    x_33 = 'b111110101;
    x_34 = 'b111110000;
    x_35 = 'b111101110;
    x_36 = 'b111101000;
    x_37 = 'b111111000;
    x_38 = 'b111100111;
    x_39 = 'b111111010;
    x_40 = 'b111100101;
    x_41 = 'b111100100;
    x_42 = 'b111100010;
    x_43 = 'b111111110;
    x_44 = 'b111100000;
    x_45 = 'b000011111;
    x_46 = 'b111111000;
    x_47 = 'b111111100;
    x_48 = 'b000000000;
    x_49 = 'b000000010;
    x_50 = 'b000000011;
    x_51 = 'b000000101;
    x_52 = 'b000000010;
    x_53 = 'b000000101;
    x_54 = 'b000001101;
    x_55 = 'b000001010;
    x_56 = 'b000000011;
    x_57 = 'b000001001;
    x_58 = 'b000001011;
    x_59 = 'b000011000;
    x_60 = 'b000010101;
    x_61 = 'b000011100;
    x_62 = 'b000000010;
    x_63 = 'b000010001;
    x_64 = 'b111111011;
    x_65 = 'b000000000;
    x_66 = 'b000000000;
    x_67 = 'b000001100;
    x_68 = 'b000001110;
    x_69 = 'b000000000;
    x_70 = 'b111111010;
    x_71 = 'b111101111;
    x_72 = 'b111111010;
    x_73 = 'b000000101;
    x_74 = 'b000001111;
    x_75 = 'b000000000;
    x_76 = 'b000000011;
    x_77 = 'b000000110;
    x_78 = 'b111110111;
    x_79 = 'b111111110;
    x_80 = 'b000000010;
    x_81 = 'b000000100;
    x_82 = 'b000000100;
    x_83 = 'b000000101;
    x_84 = 'b111111111;
    x_85 = 'b111111101;
    x_86 = 'b111111110;
    x_87 = 'b111111000;
    x_88 = 'b111101101;
    x_89 = 'b111101110;
    x_90 = 'b111110100;
    x_91 = 'b111110101;
    x_92 = 'b111111110;
    x_93 = 'b111110010;
    x_94 = 'b111101001;
    x_95 = 'b111101110;
    x_96 = 'b111110011;
    x_97 = 'b111110101;
    x_98 = 'b111110000;
    x_99 = 'b111101110;
    x_100 = 'b111101000;
    x_101 = 'b111111000;
    x_102 = 'b111100111;
    x_103 = 'b111111010;
    x_104 = 'b111100101;
    x_105 = 'b111100100;
    x_106 = 'b111100010;
    x_107 = 'b111111110;
    x_108 = 'b111100000;
    x_109 = 'b000011111;
    x_110 = 'b111111000;
    x_111 = 'b111111100;
    x_112 = 'b000000000;
    x_113 = 'b000000010;
    x_114 = 'b000000011;
    x_115 = 'b000000101;
    x_116 = 'b000000010;
    x_117 = 'b000000101;
    x_118 = 'b000001101;
    x_119 = 'b000001010;
    x_120 = 'b000000011;
    x_121 = 'b000001001;
    x_122 = 'b000001011;
    x_123 = 'b000011000;
    x_124 = 'b000010101;
    x_125 = 'b000011100;
    x_126 = 'b000000010;
    x_127 = 'b000010001;
    x_128 = 'b111111011;
    x_129 = 'b000000000;
    x_130 = 'b000000000;
    x_131 = 'b000001100;
    x_132 = 'b000001110;
    x_133 = 'b000000000;
    x_134 = 'b111111010;
    x_135 = 'b111101111;
    x_136 = 'b111111010;
    x_137 = 'b000000101;
    x_138 = 'b000001111;
    x_139 = 'b000000000;
    x_140 = 'b000000011;
    x_141 = 'b000000110;
    x_142 = 'b111110111;
    x_143 = 'b111111110;
    x_144 = 'b000000010;
    x_145 = 'b000000100;
    x_146 = 'b000000100;
    x_147 = 'b000000101;
    x_148 = 'b111111111;
    x_149 = 'b111111101;
    x_150 = 'b111111110;
    x_151 = 'b111111000;
    x_152 = 'b111101101;
    x_153 = 'b111101110;
    x_154 = 'b111110100;
    x_155 = 'b111110101;
    x_156 = 'b111111110;
    x_157 = 'b111110010;
    x_158 = 'b111101001;
    x_159 = 'b111101110;
    x_160 = 'b111110011;
    x_161 = 'b111110101;
    x_162 = 'b111110000;
    x_163 = 'b111101110;
    x_164 = 'b111101000;
    x_165 = 'b111111000;
    x_166 = 'b111100111;
    x_167 = 'b111111010;
    x_168 = 'b111100101;
    x_169 = 'b111100100;
    x_170 = 'b111100010;
    x_171 = 'b111111110;
    x_172 = 'b111100000;
    x_173 = 'b000011111;
    x_174 = 'b111111000;
    x_175 = 'b111111100;
    x_176 = 'b000000000;
    x_177 = 'b000000010;
    x_178 = 'b000000011;
    x_179 = 'b000000101;
    x_180 = 'b000000010;
    x_181 = 'b000000101;
    x_182 = 'b000001101;
    x_183 = 'b000001010;
    x_184 = 'b000000011;
    x_185 = 'b000001001;
    x_186 = 'b000001011;
    x_187 = 'b000011000;
    x_188 = 'b000010101;
    x_189 = 'b000011100;
    x_190 = 'b000000010;
    x_191 = 'b000010001;
    x_192 = 'b111111011;
    x_193 = 'b000000000;
    x_194 = 'b000000000;
    x_195 = 'b000001100;
    x_196 = 'b000001110;
    x_197 = 'b000000000;
    x_198 = 'b111111010;
    x_199 = 'b111101111;
    x_200 = 'b111111010;
    x_201 = 'b000000101;
    x_202 = 'b000001111;
    x_203 = 'b000000000;
    x_204 = 'b000000011;
    x_205 = 'b000000110;
    x_206 = 'b111110111;
    x_207 = 'b111111110;
    x_208 = 'b000000010;
    x_209 = 'b000000100;
    x_210 = 'b000000100;
    x_211 = 'b000000101;
    x_212 = 'b111111111;
    x_213 = 'b111111101;
    x_214 = 'b111111110;
    x_215 = 'b111111000;
    x_216 = 'b111101101;
    x_217 = 'b111101110;
    x_218 = 'b111110100;
    x_219 = 'b111110101;
    x_220 = 'b111111110;
    x_221 = 'b111110010;
    x_222 = 'b111101001;
    x_223 = 'b111101110;
    x_224 = 'b111110011;
    x_225 = 'b111110101;
    x_226 = 'b111110000;
    x_227 = 'b111101110;
    x_228 = 'b111101000;
    x_229 = 'b111111000;
    x_230 = 'b111100111;
    x_231 = 'b111111010;
    x_232 = 'b111100101;
    x_233 = 'b111100100;
    x_234 = 'b111100010;
    x_235 = 'b111111110;
    x_236 = 'b111100000;
    x_237 = 'b000011111;
    x_238 = 'b111111000;
    x_239 = 'b111111100;
    x_240 = 'b000000000;
    x_241 = 'b000000010;
    x_242 = 'b000000011;
    x_243 = 'b000000101;
    x_244 = 'b000000010;
    x_245 = 'b000000101;
    x_246 = 'b000001101;
    x_247 = 'b000001010;
    x_248 = 'b000000011;
    x_249 = 'b000001001;
    x_250 = 'b000001011;
    x_251 = 'b000011000;
    x_252 = 'b000010101;
    x_253 = 'b000011100;
    x_254 = 'b000000010;
    x_255 = 'b000010001;

    h_0 = 'b111111011;
    h_1 = 'b000000000;
    h_2 = 'b000000000;
    h_3 = 'b000001100;
    h_4 = 'b000001110;
    h_5 = 'b000000000;
    h_6 = 'b111111010;
    h_7 = 'b111101111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111101101;
    x_1 = 'b111110011;
    x_2 = 'b111110010;
    x_3 = 'b111111100;
    x_4 = 'b111111110;
    x_5 = 'b111110000;
    x_6 = 'b111101001;
    x_7 = 'b111100001;
    x_8 = 'b111110000;
    x_9 = 'b111111010;
    x_10 = 'b000000100;
    x_11 = 'b111101110;
    x_12 = 'b111110101;
    x_13 = 'b111111110;
    x_14 = 'b111110111;
    x_15 = 'b111111101;
    x_16 = 'b111111011;
    x_17 = 'b111111010;
    x_18 = 'b111110110;
    x_19 = 'b111111000;
    x_20 = 'b111110011;
    x_21 = 'b111111010;
    x_22 = 'b111111000;
    x_23 = 'b111110001;
    x_24 = 'b111101100;
    x_25 = 'b111101100;
    x_26 = 'b111101111;
    x_27 = 'b111101101;
    x_28 = 'b111110101;
    x_29 = 'b111110100;
    x_30 = 'b111101011;
    x_31 = 'b111100101;
    x_32 = 'b111110000;
    x_33 = 'b111101110;
    x_34 = 'b111101001;
    x_35 = 'b111101011;
    x_36 = 'b111100010;
    x_37 = 'b111110010;
    x_38 = 'b111110000;
    x_39 = 'b000000011;
    x_40 = 'b111111011;
    x_41 = 'b111111101;
    x_42 = 'b111110010;
    x_43 = 'b111101100;
    x_44 = 'b111101010;
    x_45 = 'b000001110;
    x_46 = 'b000000010;
    x_47 = 'b000000001;
    x_48 = 'b111111100;
    x_49 = 'b111111111;
    x_50 = 'b111111001;
    x_51 = 'b111111000;
    x_52 = 'b111110100;
    x_53 = 'b111110111;
    x_54 = 'b000000111;
    x_55 = 'b000001110;
    x_56 = 'b000000010;
    x_57 = 'b111111111;
    x_58 = 'b000000011;
    x_59 = 'b000011000;
    x_60 = 'b000010101;
    x_61 = 'b000011010;
    x_62 = 'b000000000;
    x_63 = 'b000010001;
    x_64 = 'b111101101;
    x_65 = 'b111110011;
    x_66 = 'b111110010;
    x_67 = 'b111111100;
    x_68 = 'b111111110;
    x_69 = 'b111110000;
    x_70 = 'b111101001;
    x_71 = 'b111100001;
    x_72 = 'b111110000;
    x_73 = 'b111111010;
    x_74 = 'b000000100;
    x_75 = 'b111101110;
    x_76 = 'b111110101;
    x_77 = 'b111111110;
    x_78 = 'b111110111;
    x_79 = 'b111111101;
    x_80 = 'b111111011;
    x_81 = 'b111111010;
    x_82 = 'b111110110;
    x_83 = 'b111111000;
    x_84 = 'b111110011;
    x_85 = 'b111111010;
    x_86 = 'b111111000;
    x_87 = 'b111110001;
    x_88 = 'b111101100;
    x_89 = 'b111101100;
    x_90 = 'b111101111;
    x_91 = 'b111101101;
    x_92 = 'b111110101;
    x_93 = 'b111110100;
    x_94 = 'b111101011;
    x_95 = 'b111100101;
    x_96 = 'b111110000;
    x_97 = 'b111101110;
    x_98 = 'b111101001;
    x_99 = 'b111101011;
    x_100 = 'b111100010;
    x_101 = 'b111110010;
    x_102 = 'b111110000;
    x_103 = 'b000000011;
    x_104 = 'b111111011;
    x_105 = 'b111111101;
    x_106 = 'b111110010;
    x_107 = 'b111101100;
    x_108 = 'b111101010;
    x_109 = 'b000001110;
    x_110 = 'b000000010;
    x_111 = 'b000000001;
    x_112 = 'b111111100;
    x_113 = 'b111111111;
    x_114 = 'b111111001;
    x_115 = 'b111111000;
    x_116 = 'b111110100;
    x_117 = 'b111110111;
    x_118 = 'b000000111;
    x_119 = 'b000001110;
    x_120 = 'b000000010;
    x_121 = 'b111111111;
    x_122 = 'b000000011;
    x_123 = 'b000011000;
    x_124 = 'b000010101;
    x_125 = 'b000011010;
    x_126 = 'b000000000;
    x_127 = 'b000010001;
    x_128 = 'b111101101;
    x_129 = 'b111110011;
    x_130 = 'b111110010;
    x_131 = 'b111111100;
    x_132 = 'b111111110;
    x_133 = 'b111110000;
    x_134 = 'b111101001;
    x_135 = 'b111100001;
    x_136 = 'b111110000;
    x_137 = 'b111111010;
    x_138 = 'b000000100;
    x_139 = 'b111101110;
    x_140 = 'b111110101;
    x_141 = 'b111111110;
    x_142 = 'b111110111;
    x_143 = 'b111111101;
    x_144 = 'b111111011;
    x_145 = 'b111111010;
    x_146 = 'b111110110;
    x_147 = 'b111111000;
    x_148 = 'b111110011;
    x_149 = 'b111111010;
    x_150 = 'b111111000;
    x_151 = 'b111110001;
    x_152 = 'b111101100;
    x_153 = 'b111101100;
    x_154 = 'b111101111;
    x_155 = 'b111101101;
    x_156 = 'b111110101;
    x_157 = 'b111110100;
    x_158 = 'b111101011;
    x_159 = 'b111100101;
    x_160 = 'b111110000;
    x_161 = 'b111101110;
    x_162 = 'b111101001;
    x_163 = 'b111101011;
    x_164 = 'b111100010;
    x_165 = 'b111110010;
    x_166 = 'b111110000;
    x_167 = 'b000000011;
    x_168 = 'b111111011;
    x_169 = 'b111111101;
    x_170 = 'b111110010;
    x_171 = 'b111101100;
    x_172 = 'b111101010;
    x_173 = 'b000001110;
    x_174 = 'b000000010;
    x_175 = 'b000000001;
    x_176 = 'b111111100;
    x_177 = 'b111111111;
    x_178 = 'b111111001;
    x_179 = 'b111111000;
    x_180 = 'b111110100;
    x_181 = 'b111110111;
    x_182 = 'b000000111;
    x_183 = 'b000001110;
    x_184 = 'b000000010;
    x_185 = 'b111111111;
    x_186 = 'b000000011;
    x_187 = 'b000011000;
    x_188 = 'b000010101;
    x_189 = 'b000011010;
    x_190 = 'b000000000;
    x_191 = 'b000010001;
    x_192 = 'b111101101;
    x_193 = 'b111110011;
    x_194 = 'b111110010;
    x_195 = 'b111111100;
    x_196 = 'b111111110;
    x_197 = 'b111110000;
    x_198 = 'b111101001;
    x_199 = 'b111100001;
    x_200 = 'b111110000;
    x_201 = 'b111111010;
    x_202 = 'b000000100;
    x_203 = 'b111101110;
    x_204 = 'b111110101;
    x_205 = 'b111111110;
    x_206 = 'b111110111;
    x_207 = 'b111111101;
    x_208 = 'b111111011;
    x_209 = 'b111111010;
    x_210 = 'b111110110;
    x_211 = 'b111111000;
    x_212 = 'b111110011;
    x_213 = 'b111111010;
    x_214 = 'b111111000;
    x_215 = 'b111110001;
    x_216 = 'b111101100;
    x_217 = 'b111101100;
    x_218 = 'b111101111;
    x_219 = 'b111101101;
    x_220 = 'b111110101;
    x_221 = 'b111110100;
    x_222 = 'b111101011;
    x_223 = 'b111100101;
    x_224 = 'b111110000;
    x_225 = 'b111101110;
    x_226 = 'b111101001;
    x_227 = 'b111101011;
    x_228 = 'b111100010;
    x_229 = 'b111110010;
    x_230 = 'b111110000;
    x_231 = 'b000000011;
    x_232 = 'b111111011;
    x_233 = 'b111111101;
    x_234 = 'b111110010;
    x_235 = 'b111101100;
    x_236 = 'b111101010;
    x_237 = 'b000001110;
    x_238 = 'b000000010;
    x_239 = 'b000000001;
    x_240 = 'b111111100;
    x_241 = 'b111111111;
    x_242 = 'b111111001;
    x_243 = 'b111111000;
    x_244 = 'b111110100;
    x_245 = 'b111110111;
    x_246 = 'b000000111;
    x_247 = 'b000001110;
    x_248 = 'b000000010;
    x_249 = 'b111111111;
    x_250 = 'b000000011;
    x_251 = 'b000011000;
    x_252 = 'b000010101;
    x_253 = 'b000011010;
    x_254 = 'b000000000;
    x_255 = 'b000010001;

    h_0 = 'b111101101;
    h_1 = 'b111110011;
    h_2 = 'b111110010;
    h_3 = 'b111111100;
    h_4 = 'b111111110;
    h_5 = 'b111110000;
    h_6 = 'b111101001;
    h_7 = 'b111100001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111110101;
    x_1 = 'b111111010;
    x_2 = 'b111110000;
    x_3 = 'b111110110;
    x_4 = 'b111110110;
    x_5 = 'b111101011;
    x_6 = 'b111101011;
    x_7 = 'b111101100;
    x_8 = 'b111110101;
    x_9 = 'b111110111;
    x_10 = 'b111111100;
    x_11 = 'b111101000;
    x_12 = 'b111101011;
    x_13 = 'b111111001;
    x_14 = 'b111111011;
    x_15 = 'b111111101;
    x_16 = 'b111110111;
    x_17 = 'b111110001;
    x_18 = 'b111101001;
    x_19 = 'b111101010;
    x_20 = 'b111100101;
    x_21 = 'b111110110;
    x_22 = 'b111110011;
    x_23 = 'b111101101;
    x_24 = 'b111101000;
    x_25 = 'b111101000;
    x_26 = 'b111101000;
    x_27 = 'b111101001;
    x_28 = 'b111110011;
    x_29 = 'b111101011;
    x_30 = 'b111100110;
    x_31 = 'b111100100;
    x_32 = 'b111101101;
    x_33 = 'b111101000;
    x_34 = 'b111100011;
    x_35 = 'b111100101;
    x_36 = 'b111100000;
    x_37 = 'b111101110;
    x_38 = 'b111101010;
    x_39 = 'b111110111;
    x_40 = 'b111101101;
    x_41 = 'b111100100;
    x_42 = 'b111100111;
    x_43 = 'b000010000;
    x_44 = 'b111101011;
    x_45 = 'b000001001;
    x_46 = 'b000000010;
    x_47 = 'b000000000;
    x_48 = 'b111111000;
    x_49 = 'b111111011;
    x_50 = 'b111110001;
    x_51 = 'b111110000;
    x_52 = 'b111101100;
    x_53 = 'b111110100;
    x_54 = 'b000000101;
    x_55 = 'b000000111;
    x_56 = 'b111111101;
    x_57 = 'b111110110;
    x_58 = 'b111111110;
    x_59 = 'b000011010;
    x_60 = 'b000010011;
    x_61 = 'b000010111;
    x_62 = 'b000000100;
    x_63 = 'b000010001;
    x_64 = 'b111110101;
    x_65 = 'b111111010;
    x_66 = 'b111110000;
    x_67 = 'b111110110;
    x_68 = 'b111110110;
    x_69 = 'b111101011;
    x_70 = 'b111101011;
    x_71 = 'b111101100;
    x_72 = 'b111110101;
    x_73 = 'b111110111;
    x_74 = 'b111111100;
    x_75 = 'b111101000;
    x_76 = 'b111101011;
    x_77 = 'b111111001;
    x_78 = 'b111111011;
    x_79 = 'b111111101;
    x_80 = 'b111110111;
    x_81 = 'b111110001;
    x_82 = 'b111101001;
    x_83 = 'b111101010;
    x_84 = 'b111100101;
    x_85 = 'b111110110;
    x_86 = 'b111110011;
    x_87 = 'b111101101;
    x_88 = 'b111101000;
    x_89 = 'b111101000;
    x_90 = 'b111101000;
    x_91 = 'b111101001;
    x_92 = 'b111110011;
    x_93 = 'b111101011;
    x_94 = 'b111100110;
    x_95 = 'b111100100;
    x_96 = 'b111101101;
    x_97 = 'b111101000;
    x_98 = 'b111100011;
    x_99 = 'b111100101;
    x_100 = 'b111100000;
    x_101 = 'b111101110;
    x_102 = 'b111101010;
    x_103 = 'b111110111;
    x_104 = 'b111101101;
    x_105 = 'b111100100;
    x_106 = 'b111100111;
    x_107 = 'b000010000;
    x_108 = 'b111101011;
    x_109 = 'b000001001;
    x_110 = 'b000000010;
    x_111 = 'b000000000;
    x_112 = 'b111111000;
    x_113 = 'b111111011;
    x_114 = 'b111110001;
    x_115 = 'b111110000;
    x_116 = 'b111101100;
    x_117 = 'b111110100;
    x_118 = 'b000000101;
    x_119 = 'b000000111;
    x_120 = 'b111111101;
    x_121 = 'b111110110;
    x_122 = 'b111111110;
    x_123 = 'b000011010;
    x_124 = 'b000010011;
    x_125 = 'b000010111;
    x_126 = 'b000000100;
    x_127 = 'b000010001;
    x_128 = 'b111110101;
    x_129 = 'b111111010;
    x_130 = 'b111110000;
    x_131 = 'b111110110;
    x_132 = 'b111110110;
    x_133 = 'b111101011;
    x_134 = 'b111101011;
    x_135 = 'b111101100;
    x_136 = 'b111110101;
    x_137 = 'b111110111;
    x_138 = 'b111111100;
    x_139 = 'b111101000;
    x_140 = 'b111101011;
    x_141 = 'b111111001;
    x_142 = 'b111111011;
    x_143 = 'b111111101;
    x_144 = 'b111110111;
    x_145 = 'b111110001;
    x_146 = 'b111101001;
    x_147 = 'b111101010;
    x_148 = 'b111100101;
    x_149 = 'b111110110;
    x_150 = 'b111110011;
    x_151 = 'b111101101;
    x_152 = 'b111101000;
    x_153 = 'b111101000;
    x_154 = 'b111101000;
    x_155 = 'b111101001;
    x_156 = 'b111110011;
    x_157 = 'b111101011;
    x_158 = 'b111100110;
    x_159 = 'b111100100;
    x_160 = 'b111101101;
    x_161 = 'b111101000;
    x_162 = 'b111100011;
    x_163 = 'b111100101;
    x_164 = 'b111100000;
    x_165 = 'b111101110;
    x_166 = 'b111101010;
    x_167 = 'b111110111;
    x_168 = 'b111101101;
    x_169 = 'b111100100;
    x_170 = 'b111100111;
    x_171 = 'b000010000;
    x_172 = 'b111101011;
    x_173 = 'b000001001;
    x_174 = 'b000000010;
    x_175 = 'b000000000;
    x_176 = 'b111111000;
    x_177 = 'b111111011;
    x_178 = 'b111110001;
    x_179 = 'b111110000;
    x_180 = 'b111101100;
    x_181 = 'b111110100;
    x_182 = 'b000000101;
    x_183 = 'b000000111;
    x_184 = 'b111111101;
    x_185 = 'b111110110;
    x_186 = 'b111111110;
    x_187 = 'b000011010;
    x_188 = 'b000010011;
    x_189 = 'b000010111;
    x_190 = 'b000000100;
    x_191 = 'b000010001;
    x_192 = 'b111110101;
    x_193 = 'b111111010;
    x_194 = 'b111110000;
    x_195 = 'b111110110;
    x_196 = 'b111110110;
    x_197 = 'b111101011;
    x_198 = 'b111101011;
    x_199 = 'b111101100;
    x_200 = 'b111110101;
    x_201 = 'b111110111;
    x_202 = 'b111111100;
    x_203 = 'b111101000;
    x_204 = 'b111101011;
    x_205 = 'b111111001;
    x_206 = 'b111111011;
    x_207 = 'b111111101;
    x_208 = 'b111110111;
    x_209 = 'b111110001;
    x_210 = 'b111101001;
    x_211 = 'b111101010;
    x_212 = 'b111100101;
    x_213 = 'b111110110;
    x_214 = 'b111110011;
    x_215 = 'b111101101;
    x_216 = 'b111101000;
    x_217 = 'b111101000;
    x_218 = 'b111101000;
    x_219 = 'b111101001;
    x_220 = 'b111110011;
    x_221 = 'b111101011;
    x_222 = 'b111100110;
    x_223 = 'b111100100;
    x_224 = 'b111101101;
    x_225 = 'b111101000;
    x_226 = 'b111100011;
    x_227 = 'b111100101;
    x_228 = 'b111100000;
    x_229 = 'b111101110;
    x_230 = 'b111101010;
    x_231 = 'b111110111;
    x_232 = 'b111101101;
    x_233 = 'b111100100;
    x_234 = 'b111100111;
    x_235 = 'b000010000;
    x_236 = 'b111101011;
    x_237 = 'b000001001;
    x_238 = 'b000000010;
    x_239 = 'b000000000;
    x_240 = 'b111111000;
    x_241 = 'b111111011;
    x_242 = 'b111110001;
    x_243 = 'b111110000;
    x_244 = 'b111101100;
    x_245 = 'b111110100;
    x_246 = 'b000000101;
    x_247 = 'b000000111;
    x_248 = 'b111111101;
    x_249 = 'b111110110;
    x_250 = 'b111111110;
    x_251 = 'b000011010;
    x_252 = 'b000010011;
    x_253 = 'b000010111;
    x_254 = 'b000000100;
    x_255 = 'b000010001;

    h_0 = 'b111110101;
    h_1 = 'b111111010;
    h_2 = 'b111110000;
    h_3 = 'b111110110;
    h_4 = 'b111110110;
    h_5 = 'b111101011;
    h_6 = 'b111101011;
    h_7 = 'b111101100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111110101;
    x_1 = 'b111111010;
    x_2 = 'b111110011;
    x_3 = 'b111110101;
    x_4 = 'b111111010;
    x_5 = 'b111110000;
    x_6 = 'b111101101;
    x_7 = 'b111110011;
    x_8 = 'b111111010;
    x_9 = 'b111111100;
    x_10 = 'b111111110;
    x_11 = 'b111101101;
    x_12 = 'b111110000;
    x_13 = 'b111111001;
    x_14 = 'b000000010;
    x_15 = 'b000000100;
    x_16 = 'b111111011;
    x_17 = 'b111110100;
    x_18 = 'b111101100;
    x_19 = 'b111101101;
    x_20 = 'b111101000;
    x_21 = 'b111111100;
    x_22 = 'b111110110;
    x_23 = 'b111101110;
    x_24 = 'b111101110;
    x_25 = 'b111101110;
    x_26 = 'b111101111;
    x_27 = 'b111101110;
    x_28 = 'b111110011;
    x_29 = 'b111110110;
    x_30 = 'b111101111;
    x_31 = 'b111101110;
    x_32 = 'b111110110;
    x_33 = 'b111110010;
    x_34 = 'b111101101;
    x_35 = 'b111110000;
    x_36 = 'b111101011;
    x_37 = 'b111110100;
    x_38 = 'b111110101;
    x_39 = 'b000000000;
    x_40 = 'b111111110;
    x_41 = 'b111011111;
    x_42 = 'b111111110;
    x_43 = 'b000010000;
    x_44 = 'b111111010;
    x_45 = 'b000010010;
    x_46 = 'b000001001;
    x_47 = 'b000000101;
    x_48 = 'b111111101;
    x_49 = 'b111111101;
    x_50 = 'b111110010;
    x_51 = 'b111110001;
    x_52 = 'b111101110;
    x_53 = 'b111110111;
    x_54 = 'b000000010;
    x_55 = 'b000000110;
    x_56 = 'b111111100;
    x_57 = 'b111110011;
    x_58 = 'b111111100;
    x_59 = 'b000010011;
    x_60 = 'b000010000;
    x_61 = 'b000010010;
    x_62 = 'b000000101;
    x_63 = 'b000001101;
    x_64 = 'b111110101;
    x_65 = 'b111111010;
    x_66 = 'b111110011;
    x_67 = 'b111110101;
    x_68 = 'b111111010;
    x_69 = 'b111110000;
    x_70 = 'b111101101;
    x_71 = 'b111110011;
    x_72 = 'b111111010;
    x_73 = 'b111111100;
    x_74 = 'b111111110;
    x_75 = 'b111101101;
    x_76 = 'b111110000;
    x_77 = 'b111111001;
    x_78 = 'b000000010;
    x_79 = 'b000000100;
    x_80 = 'b111111011;
    x_81 = 'b111110100;
    x_82 = 'b111101100;
    x_83 = 'b111101101;
    x_84 = 'b111101000;
    x_85 = 'b111111100;
    x_86 = 'b111110110;
    x_87 = 'b111101110;
    x_88 = 'b111101110;
    x_89 = 'b111101110;
    x_90 = 'b111101111;
    x_91 = 'b111101110;
    x_92 = 'b111110011;
    x_93 = 'b111110110;
    x_94 = 'b111101111;
    x_95 = 'b111101110;
    x_96 = 'b111110110;
    x_97 = 'b111110010;
    x_98 = 'b111101101;
    x_99 = 'b111110000;
    x_100 = 'b111101011;
    x_101 = 'b111110100;
    x_102 = 'b111110101;
    x_103 = 'b000000000;
    x_104 = 'b111111110;
    x_105 = 'b111011111;
    x_106 = 'b111111110;
    x_107 = 'b000010000;
    x_108 = 'b111111010;
    x_109 = 'b000010010;
    x_110 = 'b000001001;
    x_111 = 'b000000101;
    x_112 = 'b111111101;
    x_113 = 'b111111101;
    x_114 = 'b111110010;
    x_115 = 'b111110001;
    x_116 = 'b111101110;
    x_117 = 'b111110111;
    x_118 = 'b000000010;
    x_119 = 'b000000110;
    x_120 = 'b111111100;
    x_121 = 'b111110011;
    x_122 = 'b111111100;
    x_123 = 'b000010011;
    x_124 = 'b000010000;
    x_125 = 'b000010010;
    x_126 = 'b000000101;
    x_127 = 'b000001101;
    x_128 = 'b111110101;
    x_129 = 'b111111010;
    x_130 = 'b111110011;
    x_131 = 'b111110101;
    x_132 = 'b111111010;
    x_133 = 'b111110000;
    x_134 = 'b111101101;
    x_135 = 'b111110011;
    x_136 = 'b111111010;
    x_137 = 'b111111100;
    x_138 = 'b111111110;
    x_139 = 'b111101101;
    x_140 = 'b111110000;
    x_141 = 'b111111001;
    x_142 = 'b000000010;
    x_143 = 'b000000100;
    x_144 = 'b111111011;
    x_145 = 'b111110100;
    x_146 = 'b111101100;
    x_147 = 'b111101101;
    x_148 = 'b111101000;
    x_149 = 'b111111100;
    x_150 = 'b111110110;
    x_151 = 'b111101110;
    x_152 = 'b111101110;
    x_153 = 'b111101110;
    x_154 = 'b111101111;
    x_155 = 'b111101110;
    x_156 = 'b111110011;
    x_157 = 'b111110110;
    x_158 = 'b111101111;
    x_159 = 'b111101110;
    x_160 = 'b111110110;
    x_161 = 'b111110010;
    x_162 = 'b111101101;
    x_163 = 'b111110000;
    x_164 = 'b111101011;
    x_165 = 'b111110100;
    x_166 = 'b111110101;
    x_167 = 'b000000000;
    x_168 = 'b111111110;
    x_169 = 'b111011111;
    x_170 = 'b111111110;
    x_171 = 'b000010000;
    x_172 = 'b111111010;
    x_173 = 'b000010010;
    x_174 = 'b000001001;
    x_175 = 'b000000101;
    x_176 = 'b111111101;
    x_177 = 'b111111101;
    x_178 = 'b111110010;
    x_179 = 'b111110001;
    x_180 = 'b111101110;
    x_181 = 'b111110111;
    x_182 = 'b000000010;
    x_183 = 'b000000110;
    x_184 = 'b111111100;
    x_185 = 'b111110011;
    x_186 = 'b111111100;
    x_187 = 'b000010011;
    x_188 = 'b000010000;
    x_189 = 'b000010010;
    x_190 = 'b000000101;
    x_191 = 'b000001101;
    x_192 = 'b111110101;
    x_193 = 'b111111010;
    x_194 = 'b111110011;
    x_195 = 'b111110101;
    x_196 = 'b111111010;
    x_197 = 'b111110000;
    x_198 = 'b111101101;
    x_199 = 'b111110011;
    x_200 = 'b111111010;
    x_201 = 'b111111100;
    x_202 = 'b111111110;
    x_203 = 'b111101101;
    x_204 = 'b111110000;
    x_205 = 'b111111001;
    x_206 = 'b000000010;
    x_207 = 'b000000100;
    x_208 = 'b111111011;
    x_209 = 'b111110100;
    x_210 = 'b111101100;
    x_211 = 'b111101101;
    x_212 = 'b111101000;
    x_213 = 'b111111100;
    x_214 = 'b111110110;
    x_215 = 'b111101110;
    x_216 = 'b111101110;
    x_217 = 'b111101110;
    x_218 = 'b111101111;
    x_219 = 'b111101110;
    x_220 = 'b111110011;
    x_221 = 'b111110110;
    x_222 = 'b111101111;
    x_223 = 'b111101110;
    x_224 = 'b111110110;
    x_225 = 'b111110010;
    x_226 = 'b111101101;
    x_227 = 'b111110000;
    x_228 = 'b111101011;
    x_229 = 'b111110100;
    x_230 = 'b111110101;
    x_231 = 'b000000000;
    x_232 = 'b111111110;
    x_233 = 'b111011111;
    x_234 = 'b111111110;
    x_235 = 'b000010000;
    x_236 = 'b111111010;
    x_237 = 'b000010010;
    x_238 = 'b000001001;
    x_239 = 'b000000101;
    x_240 = 'b111111101;
    x_241 = 'b111111101;
    x_242 = 'b111110010;
    x_243 = 'b111110001;
    x_244 = 'b111101110;
    x_245 = 'b111110111;
    x_246 = 'b000000010;
    x_247 = 'b000000110;
    x_248 = 'b111111100;
    x_249 = 'b111110011;
    x_250 = 'b111111100;
    x_251 = 'b000010011;
    x_252 = 'b000010000;
    x_253 = 'b000010010;
    x_254 = 'b000000101;
    x_255 = 'b000001101;

    h_0 = 'b111110101;
    h_1 = 'b111111010;
    h_2 = 'b111110011;
    h_3 = 'b111110101;
    h_4 = 'b111111010;
    h_5 = 'b111110000;
    h_6 = 'b111101101;
    h_7 = 'b111110011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000000001;
    x_1 = 'b000000011;
    x_2 = 'b111111010;
    x_3 = 'b111111011;
    x_4 = 'b000000010;
    x_5 = 'b111111110;
    x_6 = 'b111111111;
    x_7 = 'b111111011;
    x_8 = 'b000000000;
    x_9 = 'b000000010;
    x_10 = 'b000000100;
    x_11 = 'b111110100;
    x_12 = 'b111111111;
    x_13 = 'b000001001;
    x_14 = 'b000001001;
    x_15 = 'b000000111;
    x_16 = 'b000000000;
    x_17 = 'b111111001;
    x_18 = 'b111110110;
    x_19 = 'b111111001;
    x_20 = 'b111110101;
    x_21 = 'b000000111;
    x_22 = 'b000000011;
    x_23 = 'b111111010;
    x_24 = 'b111111010;
    x_25 = 'b111111001;
    x_26 = 'b111110110;
    x_27 = 'b111111011;
    x_28 = 'b111111111;
    x_29 = 'b000000101;
    x_30 = 'b111111011;
    x_31 = 'b111110011;
    x_32 = 'b111111010;
    x_33 = 'b111110101;
    x_34 = 'b111110011;
    x_35 = 'b111111000;
    x_36 = 'b111111000;
    x_37 = 'b111111111;
    x_38 = 'b000000001;
    x_39 = 'b000010110;
    x_40 = 'b000010000;
    x_41 = 'b000000101;
    x_42 = 'b000000111;
    x_43 = 'b000010001;
    x_44 = 'b111111110;
    x_45 = 'b000011001;
    x_46 = 'b000001101;
    x_47 = 'b000001011;
    x_48 = 'b000000010;
    x_49 = 'b111111111;
    x_50 = 'b111110111;
    x_51 = 'b111110010;
    x_52 = 'b111110010;
    x_53 = 'b111111010;
    x_54 = 'b111111111;
    x_55 = 'b000001001;
    x_56 = 'b000000010;
    x_57 = 'b111110101;
    x_58 = 'b111110110;
    x_59 = 'b000000110;
    x_60 = 'b000001001;
    x_61 = 'b000000101;
    x_62 = 'b111111001;
    x_63 = 'b111111111;
    x_64 = 'b000000001;
    x_65 = 'b000000011;
    x_66 = 'b111111010;
    x_67 = 'b111111011;
    x_68 = 'b000000010;
    x_69 = 'b111111110;
    x_70 = 'b111111111;
    x_71 = 'b111111011;
    x_72 = 'b000000000;
    x_73 = 'b000000010;
    x_74 = 'b000000100;
    x_75 = 'b111110100;
    x_76 = 'b111111111;
    x_77 = 'b000001001;
    x_78 = 'b000001001;
    x_79 = 'b000000111;
    x_80 = 'b000000000;
    x_81 = 'b111111001;
    x_82 = 'b111110110;
    x_83 = 'b111111001;
    x_84 = 'b111110101;
    x_85 = 'b000000111;
    x_86 = 'b000000011;
    x_87 = 'b111111010;
    x_88 = 'b111111010;
    x_89 = 'b111111001;
    x_90 = 'b111110110;
    x_91 = 'b111111011;
    x_92 = 'b111111111;
    x_93 = 'b000000101;
    x_94 = 'b111111011;
    x_95 = 'b111110011;
    x_96 = 'b111111010;
    x_97 = 'b111110101;
    x_98 = 'b111110011;
    x_99 = 'b111111000;
    x_100 = 'b111111000;
    x_101 = 'b111111111;
    x_102 = 'b000000001;
    x_103 = 'b000010110;
    x_104 = 'b000010000;
    x_105 = 'b000000101;
    x_106 = 'b000000111;
    x_107 = 'b000010001;
    x_108 = 'b111111110;
    x_109 = 'b000011001;
    x_110 = 'b000001101;
    x_111 = 'b000001011;
    x_112 = 'b000000010;
    x_113 = 'b111111111;
    x_114 = 'b111110111;
    x_115 = 'b111110010;
    x_116 = 'b111110010;
    x_117 = 'b111111010;
    x_118 = 'b111111111;
    x_119 = 'b000001001;
    x_120 = 'b000000010;
    x_121 = 'b111110101;
    x_122 = 'b111110110;
    x_123 = 'b000000110;
    x_124 = 'b000001001;
    x_125 = 'b000000101;
    x_126 = 'b111111001;
    x_127 = 'b111111111;
    x_128 = 'b000000001;
    x_129 = 'b000000011;
    x_130 = 'b111111010;
    x_131 = 'b111111011;
    x_132 = 'b000000010;
    x_133 = 'b111111110;
    x_134 = 'b111111111;
    x_135 = 'b111111011;
    x_136 = 'b000000000;
    x_137 = 'b000000010;
    x_138 = 'b000000100;
    x_139 = 'b111110100;
    x_140 = 'b111111111;
    x_141 = 'b000001001;
    x_142 = 'b000001001;
    x_143 = 'b000000111;
    x_144 = 'b000000000;
    x_145 = 'b111111001;
    x_146 = 'b111110110;
    x_147 = 'b111111001;
    x_148 = 'b111110101;
    x_149 = 'b000000111;
    x_150 = 'b000000011;
    x_151 = 'b111111010;
    x_152 = 'b111111010;
    x_153 = 'b111111001;
    x_154 = 'b111110110;
    x_155 = 'b111111011;
    x_156 = 'b111111111;
    x_157 = 'b000000101;
    x_158 = 'b111111011;
    x_159 = 'b111110011;
    x_160 = 'b111111010;
    x_161 = 'b111110101;
    x_162 = 'b111110011;
    x_163 = 'b111111000;
    x_164 = 'b111111000;
    x_165 = 'b111111111;
    x_166 = 'b000000001;
    x_167 = 'b000010110;
    x_168 = 'b000010000;
    x_169 = 'b000000101;
    x_170 = 'b000000111;
    x_171 = 'b000010001;
    x_172 = 'b111111110;
    x_173 = 'b000011001;
    x_174 = 'b000001101;
    x_175 = 'b000001011;
    x_176 = 'b000000010;
    x_177 = 'b111111111;
    x_178 = 'b111110111;
    x_179 = 'b111110010;
    x_180 = 'b111110010;
    x_181 = 'b111111010;
    x_182 = 'b111111111;
    x_183 = 'b000001001;
    x_184 = 'b000000010;
    x_185 = 'b111110101;
    x_186 = 'b111110110;
    x_187 = 'b000000110;
    x_188 = 'b000001001;
    x_189 = 'b000000101;
    x_190 = 'b111111001;
    x_191 = 'b111111111;
    x_192 = 'b000000001;
    x_193 = 'b000000011;
    x_194 = 'b111111010;
    x_195 = 'b111111011;
    x_196 = 'b000000010;
    x_197 = 'b111111110;
    x_198 = 'b111111111;
    x_199 = 'b111111011;
    x_200 = 'b000000000;
    x_201 = 'b000000010;
    x_202 = 'b000000100;
    x_203 = 'b111110100;
    x_204 = 'b111111111;
    x_205 = 'b000001001;
    x_206 = 'b000001001;
    x_207 = 'b000000111;
    x_208 = 'b000000000;
    x_209 = 'b111111001;
    x_210 = 'b111110110;
    x_211 = 'b111111001;
    x_212 = 'b111110101;
    x_213 = 'b000000111;
    x_214 = 'b000000011;
    x_215 = 'b111111010;
    x_216 = 'b111111010;
    x_217 = 'b111111001;
    x_218 = 'b111110110;
    x_219 = 'b111111011;
    x_220 = 'b111111111;
    x_221 = 'b000000101;
    x_222 = 'b111111011;
    x_223 = 'b111110011;
    x_224 = 'b111111010;
    x_225 = 'b111110101;
    x_226 = 'b111110011;
    x_227 = 'b111111000;
    x_228 = 'b111111000;
    x_229 = 'b111111111;
    x_230 = 'b000000001;
    x_231 = 'b000010110;
    x_232 = 'b000010000;
    x_233 = 'b000000101;
    x_234 = 'b000000111;
    x_235 = 'b000010001;
    x_236 = 'b111111110;
    x_237 = 'b000011001;
    x_238 = 'b000001101;
    x_239 = 'b000001011;
    x_240 = 'b000000010;
    x_241 = 'b111111111;
    x_242 = 'b111110111;
    x_243 = 'b111110010;
    x_244 = 'b111110010;
    x_245 = 'b111111010;
    x_246 = 'b111111111;
    x_247 = 'b000001001;
    x_248 = 'b000000010;
    x_249 = 'b111110101;
    x_250 = 'b111110110;
    x_251 = 'b000000110;
    x_252 = 'b000001001;
    x_253 = 'b000000101;
    x_254 = 'b111111001;
    x_255 = 'b111111111;

    h_0 = 'b000000001;
    h_1 = 'b000000011;
    h_2 = 'b111111010;
    h_3 = 'b111111011;
    h_4 = 'b000000010;
    h_5 = 'b111111110;
    h_6 = 'b111111111;
    h_7 = 'b111111011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000001000;
    x_1 = 'b000001000;
    x_2 = 'b111111111;
    x_3 = 'b000000000;
    x_4 = 'b000000100;
    x_5 = 'b000000000;
    x_6 = 'b000000000;
    x_7 = 'b000000100;
    x_8 = 'b000000111;
    x_9 = 'b000001010;
    x_10 = 'b000010001;
    x_11 = 'b111111011;
    x_12 = 'b000000111;
    x_13 = 'b000001110;
    x_14 = 'b000010101;
    x_15 = 'b000010000;
    x_16 = 'b000001000;
    x_17 = 'b000000010;
    x_18 = 'b111111110;
    x_19 = 'b000000010;
    x_20 = 'b111111110;
    x_21 = 'b111111111;
    x_22 = 'b000000000;
    x_23 = 'b111111000;
    x_24 = 'b111110110;
    x_25 = 'b111110101;
    x_26 = 'b111110001;
    x_27 = 'b111111000;
    x_28 = 'b000000000;
    x_29 = 'b000000000;
    x_30 = 'b111110101;
    x_31 = 'b111110001;
    x_32 = 'b111111000;
    x_33 = 'b111110010;
    x_34 = 'b111101101;
    x_35 = 'b111110001;
    x_36 = 'b111110000;
    x_37 = 'b111110010;
    x_38 = 'b000000000;
    x_39 = 'b000001011;
    x_40 = 'b000011000;
    x_41 = 'b111101110;
    x_42 = 'b111110001;
    x_43 = 'b000011110;
    x_44 = 'b000000101;
    x_45 = 'b000011011;
    x_46 = 'b000011101;
    x_47 = 'b000011010;
    x_48 = 'b000001101;
    x_49 = 'b000001101;
    x_50 = 'b000000010;
    x_51 = 'b111110101;
    x_52 = 'b111110100;
    x_53 = 'b111111010;
    x_54 = 'b111111011;
    x_55 = 'b000010010;
    x_56 = 'b000010000;
    x_57 = 'b111111010;
    x_58 = 'b111101101;
    x_59 = 'b111111000;
    x_60 = 'b000001001;
    x_61 = 'b111111001;
    x_62 = 'b111100101;
    x_63 = 'b111110110;
    x_64 = 'b000001000;
    x_65 = 'b000001000;
    x_66 = 'b111111111;
    x_67 = 'b000000000;
    x_68 = 'b000000100;
    x_69 = 'b000000000;
    x_70 = 'b000000000;
    x_71 = 'b000000100;
    x_72 = 'b000000111;
    x_73 = 'b000001010;
    x_74 = 'b000010001;
    x_75 = 'b111111011;
    x_76 = 'b000000111;
    x_77 = 'b000001110;
    x_78 = 'b000010101;
    x_79 = 'b000010000;
    x_80 = 'b000001000;
    x_81 = 'b000000010;
    x_82 = 'b111111110;
    x_83 = 'b000000010;
    x_84 = 'b111111110;
    x_85 = 'b111111111;
    x_86 = 'b000000000;
    x_87 = 'b111111000;
    x_88 = 'b111110110;
    x_89 = 'b111110101;
    x_90 = 'b111110001;
    x_91 = 'b111111000;
    x_92 = 'b000000000;
    x_93 = 'b000000000;
    x_94 = 'b111110101;
    x_95 = 'b111110001;
    x_96 = 'b111111000;
    x_97 = 'b111110010;
    x_98 = 'b111101101;
    x_99 = 'b111110001;
    x_100 = 'b111110000;
    x_101 = 'b111110010;
    x_102 = 'b000000000;
    x_103 = 'b000001011;
    x_104 = 'b000011000;
    x_105 = 'b111101110;
    x_106 = 'b111110001;
    x_107 = 'b000011110;
    x_108 = 'b000000101;
    x_109 = 'b000011011;
    x_110 = 'b000011101;
    x_111 = 'b000011010;
    x_112 = 'b000001101;
    x_113 = 'b000001101;
    x_114 = 'b000000010;
    x_115 = 'b111110101;
    x_116 = 'b111110100;
    x_117 = 'b111111010;
    x_118 = 'b111111011;
    x_119 = 'b000010010;
    x_120 = 'b000010000;
    x_121 = 'b111111010;
    x_122 = 'b111101101;
    x_123 = 'b111111000;
    x_124 = 'b000001001;
    x_125 = 'b111111001;
    x_126 = 'b111100101;
    x_127 = 'b111110110;
    x_128 = 'b000001000;
    x_129 = 'b000001000;
    x_130 = 'b111111111;
    x_131 = 'b000000000;
    x_132 = 'b000000100;
    x_133 = 'b000000000;
    x_134 = 'b000000000;
    x_135 = 'b000000100;
    x_136 = 'b000000111;
    x_137 = 'b000001010;
    x_138 = 'b000010001;
    x_139 = 'b111111011;
    x_140 = 'b000000111;
    x_141 = 'b000001110;
    x_142 = 'b000010101;
    x_143 = 'b000010000;
    x_144 = 'b000001000;
    x_145 = 'b000000010;
    x_146 = 'b111111110;
    x_147 = 'b000000010;
    x_148 = 'b111111110;
    x_149 = 'b111111111;
    x_150 = 'b000000000;
    x_151 = 'b111111000;
    x_152 = 'b111110110;
    x_153 = 'b111110101;
    x_154 = 'b111110001;
    x_155 = 'b111111000;
    x_156 = 'b000000000;
    x_157 = 'b000000000;
    x_158 = 'b111110101;
    x_159 = 'b111110001;
    x_160 = 'b111111000;
    x_161 = 'b111110010;
    x_162 = 'b111101101;
    x_163 = 'b111110001;
    x_164 = 'b111110000;
    x_165 = 'b111110010;
    x_166 = 'b000000000;
    x_167 = 'b000001011;
    x_168 = 'b000011000;
    x_169 = 'b111101110;
    x_170 = 'b111110001;
    x_171 = 'b000011110;
    x_172 = 'b000000101;
    x_173 = 'b000011011;
    x_174 = 'b000011101;
    x_175 = 'b000011010;
    x_176 = 'b000001101;
    x_177 = 'b000001101;
    x_178 = 'b000000010;
    x_179 = 'b111110101;
    x_180 = 'b111110100;
    x_181 = 'b111111010;
    x_182 = 'b111111011;
    x_183 = 'b000010010;
    x_184 = 'b000010000;
    x_185 = 'b111111010;
    x_186 = 'b111101101;
    x_187 = 'b111111000;
    x_188 = 'b000001001;
    x_189 = 'b111111001;
    x_190 = 'b111100101;
    x_191 = 'b111110110;
    x_192 = 'b000001000;
    x_193 = 'b000001000;
    x_194 = 'b111111111;
    x_195 = 'b000000000;
    x_196 = 'b000000100;
    x_197 = 'b000000000;
    x_198 = 'b000000000;
    x_199 = 'b000000100;
    x_200 = 'b000000111;
    x_201 = 'b000001010;
    x_202 = 'b000010001;
    x_203 = 'b111111011;
    x_204 = 'b000000111;
    x_205 = 'b000001110;
    x_206 = 'b000010101;
    x_207 = 'b000010000;
    x_208 = 'b000001000;
    x_209 = 'b000000010;
    x_210 = 'b111111110;
    x_211 = 'b000000010;
    x_212 = 'b111111110;
    x_213 = 'b111111111;
    x_214 = 'b000000000;
    x_215 = 'b111111000;
    x_216 = 'b111110110;
    x_217 = 'b111110101;
    x_218 = 'b111110001;
    x_219 = 'b111111000;
    x_220 = 'b000000000;
    x_221 = 'b000000000;
    x_222 = 'b111110101;
    x_223 = 'b111110001;
    x_224 = 'b111111000;
    x_225 = 'b111110010;
    x_226 = 'b111101101;
    x_227 = 'b111110001;
    x_228 = 'b111110000;
    x_229 = 'b111110010;
    x_230 = 'b000000000;
    x_231 = 'b000001011;
    x_232 = 'b000011000;
    x_233 = 'b111101110;
    x_234 = 'b111110001;
    x_235 = 'b000011110;
    x_236 = 'b000000101;
    x_237 = 'b000011011;
    x_238 = 'b000011101;
    x_239 = 'b000011010;
    x_240 = 'b000001101;
    x_241 = 'b000001101;
    x_242 = 'b000000010;
    x_243 = 'b111110101;
    x_244 = 'b111110100;
    x_245 = 'b111111010;
    x_246 = 'b111111011;
    x_247 = 'b000010010;
    x_248 = 'b000010000;
    x_249 = 'b111111010;
    x_250 = 'b111101101;
    x_251 = 'b111111000;
    x_252 = 'b000001001;
    x_253 = 'b111111001;
    x_254 = 'b111100101;
    x_255 = 'b111110110;

    h_0 = 'b000001000;
    h_1 = 'b000001000;
    h_2 = 'b111111111;
    h_3 = 'b000000000;
    h_4 = 'b000000100;
    h_5 = 'b000000000;
    h_6 = 'b000000000;
    h_7 = 'b000000100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000001011;
    x_1 = 'b000001001;
    x_2 = 'b000000001;
    x_3 = 'b000000110;
    x_4 = 'b000001001;
    x_5 = 'b000000000;
    x_6 = 'b111110101;
    x_7 = 'b000001000;
    x_8 = 'b000000111;
    x_9 = 'b000001100;
    x_10 = 'b000010101;
    x_11 = 'b000000000;
    x_12 = 'b000001011;
    x_13 = 'b000001111;
    x_14 = 'b000010110;
    x_15 = 'b000001111;
    x_16 = 'b000001100;
    x_17 = 'b000001001;
    x_18 = 'b000000010;
    x_19 = 'b000000011;
    x_20 = 'b111111111;
    x_21 = 'b111111011;
    x_22 = 'b111111101;
    x_23 = 'b111110101;
    x_24 = 'b111110101;
    x_25 = 'b111110100;
    x_26 = 'b111110011;
    x_27 = 'b111110100;
    x_28 = 'b111111010;
    x_29 = 'b000000000;
    x_30 = 'b111110011;
    x_31 = 'b111110010;
    x_32 = 'b111111110;
    x_33 = 'b111111000;
    x_34 = 'b111110001;
    x_35 = 'b111110111;
    x_36 = 'b111101110;
    x_37 = 'b111101100;
    x_38 = 'b000000100;
    x_39 = 'b000000001;
    x_40 = 'b000001010;
    x_41 = 'b111011010;
    x_42 = 'b111110011;
    x_43 = 'b000010000;
    x_44 = 'b111110111;
    x_45 = 'b000001101;
    x_46 = 'b000001010;
    x_47 = 'b000001110;
    x_48 = 'b000000110;
    x_49 = 'b000001001;
    x_50 = 'b111111110;
    x_51 = 'b111101011;
    x_52 = 'b111101010;
    x_53 = 'b111100111;
    x_54 = 'b111100101;
    x_55 = 'b000000011;
    x_56 = 'b000000110;
    x_57 = 'b111101110;
    x_58 = 'b111010100;
    x_59 = 'b111010011;
    x_60 = 'b000000000;
    x_61 = 'b111100111;
    x_62 = 'b111000110;
    x_63 = 'b111100011;
    x_64 = 'b000001011;
    x_65 = 'b000001001;
    x_66 = 'b000000001;
    x_67 = 'b000000110;
    x_68 = 'b000001001;
    x_69 = 'b000000000;
    x_70 = 'b111110101;
    x_71 = 'b000001000;
    x_72 = 'b000000111;
    x_73 = 'b000001100;
    x_74 = 'b000010101;
    x_75 = 'b000000000;
    x_76 = 'b000001011;
    x_77 = 'b000001111;
    x_78 = 'b000010110;
    x_79 = 'b000001111;
    x_80 = 'b000001100;
    x_81 = 'b000001001;
    x_82 = 'b000000010;
    x_83 = 'b000000011;
    x_84 = 'b111111111;
    x_85 = 'b111111011;
    x_86 = 'b111111101;
    x_87 = 'b111110101;
    x_88 = 'b111110101;
    x_89 = 'b111110100;
    x_90 = 'b111110011;
    x_91 = 'b111110100;
    x_92 = 'b111111010;
    x_93 = 'b000000000;
    x_94 = 'b111110011;
    x_95 = 'b111110010;
    x_96 = 'b111111110;
    x_97 = 'b111111000;
    x_98 = 'b111110001;
    x_99 = 'b111110111;
    x_100 = 'b111101110;
    x_101 = 'b111101100;
    x_102 = 'b000000100;
    x_103 = 'b000000001;
    x_104 = 'b000001010;
    x_105 = 'b111011010;
    x_106 = 'b111110011;
    x_107 = 'b000010000;
    x_108 = 'b111110111;
    x_109 = 'b000001101;
    x_110 = 'b000001010;
    x_111 = 'b000001110;
    x_112 = 'b000000110;
    x_113 = 'b000001001;
    x_114 = 'b111111110;
    x_115 = 'b111101011;
    x_116 = 'b111101010;
    x_117 = 'b111100111;
    x_118 = 'b111100101;
    x_119 = 'b000000011;
    x_120 = 'b000000110;
    x_121 = 'b111101110;
    x_122 = 'b111010100;
    x_123 = 'b111010011;
    x_124 = 'b000000000;
    x_125 = 'b111100111;
    x_126 = 'b111000110;
    x_127 = 'b111100011;
    x_128 = 'b000001011;
    x_129 = 'b000001001;
    x_130 = 'b000000001;
    x_131 = 'b000000110;
    x_132 = 'b000001001;
    x_133 = 'b000000000;
    x_134 = 'b111110101;
    x_135 = 'b000001000;
    x_136 = 'b000000111;
    x_137 = 'b000001100;
    x_138 = 'b000010101;
    x_139 = 'b000000000;
    x_140 = 'b000001011;
    x_141 = 'b000001111;
    x_142 = 'b000010110;
    x_143 = 'b000001111;
    x_144 = 'b000001100;
    x_145 = 'b000001001;
    x_146 = 'b000000010;
    x_147 = 'b000000011;
    x_148 = 'b111111111;
    x_149 = 'b111111011;
    x_150 = 'b111111101;
    x_151 = 'b111110101;
    x_152 = 'b111110101;
    x_153 = 'b111110100;
    x_154 = 'b111110011;
    x_155 = 'b111110100;
    x_156 = 'b111111010;
    x_157 = 'b000000000;
    x_158 = 'b111110011;
    x_159 = 'b111110010;
    x_160 = 'b111111110;
    x_161 = 'b111111000;
    x_162 = 'b111110001;
    x_163 = 'b111110111;
    x_164 = 'b111101110;
    x_165 = 'b111101100;
    x_166 = 'b000000100;
    x_167 = 'b000000001;
    x_168 = 'b000001010;
    x_169 = 'b111011010;
    x_170 = 'b111110011;
    x_171 = 'b000010000;
    x_172 = 'b111110111;
    x_173 = 'b000001101;
    x_174 = 'b000001010;
    x_175 = 'b000001110;
    x_176 = 'b000000110;
    x_177 = 'b000001001;
    x_178 = 'b111111110;
    x_179 = 'b111101011;
    x_180 = 'b111101010;
    x_181 = 'b111100111;
    x_182 = 'b111100101;
    x_183 = 'b000000011;
    x_184 = 'b000000110;
    x_185 = 'b111101110;
    x_186 = 'b111010100;
    x_187 = 'b111010011;
    x_188 = 'b000000000;
    x_189 = 'b111100111;
    x_190 = 'b111000110;
    x_191 = 'b111100011;
    x_192 = 'b000001011;
    x_193 = 'b000001001;
    x_194 = 'b000000001;
    x_195 = 'b000000110;
    x_196 = 'b000001001;
    x_197 = 'b000000000;
    x_198 = 'b111110101;
    x_199 = 'b000001000;
    x_200 = 'b000000111;
    x_201 = 'b000001100;
    x_202 = 'b000010101;
    x_203 = 'b000000000;
    x_204 = 'b000001011;
    x_205 = 'b000001111;
    x_206 = 'b000010110;
    x_207 = 'b000001111;
    x_208 = 'b000001100;
    x_209 = 'b000001001;
    x_210 = 'b000000010;
    x_211 = 'b000000011;
    x_212 = 'b111111111;
    x_213 = 'b111111011;
    x_214 = 'b111111101;
    x_215 = 'b111110101;
    x_216 = 'b111110101;
    x_217 = 'b111110100;
    x_218 = 'b111110011;
    x_219 = 'b111110100;
    x_220 = 'b111111010;
    x_221 = 'b000000000;
    x_222 = 'b111110011;
    x_223 = 'b111110010;
    x_224 = 'b111111110;
    x_225 = 'b111111000;
    x_226 = 'b111110001;
    x_227 = 'b111110111;
    x_228 = 'b111101110;
    x_229 = 'b111101100;
    x_230 = 'b000000100;
    x_231 = 'b000000001;
    x_232 = 'b000001010;
    x_233 = 'b111011010;
    x_234 = 'b111110011;
    x_235 = 'b000010000;
    x_236 = 'b111110111;
    x_237 = 'b000001101;
    x_238 = 'b000001010;
    x_239 = 'b000001110;
    x_240 = 'b000000110;
    x_241 = 'b000001001;
    x_242 = 'b111111110;
    x_243 = 'b111101011;
    x_244 = 'b111101010;
    x_245 = 'b111100111;
    x_246 = 'b111100101;
    x_247 = 'b000000011;
    x_248 = 'b000000110;
    x_249 = 'b111101110;
    x_250 = 'b111010100;
    x_251 = 'b111010011;
    x_252 = 'b000000000;
    x_253 = 'b111100111;
    x_254 = 'b111000110;
    x_255 = 'b111100011;

    h_0 = 'b000001011;
    h_1 = 'b000001001;
    h_2 = 'b000000001;
    h_3 = 'b000000110;
    h_4 = 'b000001001;
    h_5 = 'b000000000;
    h_6 = 'b111110101;
    h_7 = 'b000001000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000001110;
    x_1 = 'b000001110;
    x_2 = 'b000001001;
    x_3 = 'b000001111;
    x_4 = 'b000010101;
    x_5 = 'b000001011;
    x_6 = 'b000000000;
    x_7 = 'b000000000;
    x_8 = 'b000000101;
    x_9 = 'b000001111;
    x_10 = 'b000011100;
    x_11 = 'b000001101;
    x_12 = 'b000001110;
    x_13 = 'b000001110;
    x_14 = 'b000000100;
    x_15 = 'b000000111;
    x_16 = 'b000001010;
    x_17 = 'b000001010;
    x_18 = 'b000000011;
    x_19 = 'b111111111;
    x_20 = 'b111111000;
    x_21 = 'b000000011;
    x_22 = 'b000000101;
    x_23 = 'b111111110;
    x_24 = 'b111111001;
    x_25 = 'b111111000;
    x_26 = 'b000000000;
    x_27 = 'b000000010;
    x_28 = 'b000000110;
    x_29 = 'b111111011;
    x_30 = 'b111111010;
    x_31 = 'b111111111;
    x_32 = 'b000001000;
    x_33 = 'b000001000;
    x_34 = 'b000000000;
    x_35 = 'b000000011;
    x_36 = 'b000000010;
    x_37 = 'b000000100;
    x_38 = 'b111111110;
    x_39 = 'b000011000;
    x_40 = 'b111111110;
    x_41 = 'b111100011;
    x_42 = 'b111100111;
    x_43 = 'b000000001;
    x_44 = 'b111100111;
    x_45 = 'b000000101;
    x_46 = 'b111110011;
    x_47 = 'b111111010;
    x_48 = 'b111110111;
    x_49 = 'b111111111;
    x_50 = 'b111111001;
    x_51 = 'b111100001;
    x_52 = 'b111011111;
    x_53 = 'b111010110;
    x_54 = 'b111010000;
    x_55 = 'b111101111;
    x_56 = 'b111110010;
    x_57 = 'b111100001;
    x_58 = 'b111000011;
    x_59 = 'b110110100;
    x_60 = 'b111101011;
    x_61 = 'b111001100;
    x_62 = 'b110100011;
    x_63 = 'b111000110;
    x_64 = 'b000001110;
    x_65 = 'b000001110;
    x_66 = 'b000001001;
    x_67 = 'b000001111;
    x_68 = 'b000010101;
    x_69 = 'b000001011;
    x_70 = 'b000000000;
    x_71 = 'b000000000;
    x_72 = 'b000000101;
    x_73 = 'b000001111;
    x_74 = 'b000011100;
    x_75 = 'b000001101;
    x_76 = 'b000001110;
    x_77 = 'b000001110;
    x_78 = 'b000000100;
    x_79 = 'b000000111;
    x_80 = 'b000001010;
    x_81 = 'b000001010;
    x_82 = 'b000000011;
    x_83 = 'b111111111;
    x_84 = 'b111111000;
    x_85 = 'b000000011;
    x_86 = 'b000000101;
    x_87 = 'b111111110;
    x_88 = 'b111111001;
    x_89 = 'b111111000;
    x_90 = 'b000000000;
    x_91 = 'b000000010;
    x_92 = 'b000000110;
    x_93 = 'b111111011;
    x_94 = 'b111111010;
    x_95 = 'b111111111;
    x_96 = 'b000001000;
    x_97 = 'b000001000;
    x_98 = 'b000000000;
    x_99 = 'b000000011;
    x_100 = 'b000000010;
    x_101 = 'b000000100;
    x_102 = 'b111111110;
    x_103 = 'b000011000;
    x_104 = 'b111111110;
    x_105 = 'b111100011;
    x_106 = 'b111100111;
    x_107 = 'b000000001;
    x_108 = 'b111100111;
    x_109 = 'b000000101;
    x_110 = 'b111110011;
    x_111 = 'b111111010;
    x_112 = 'b111110111;
    x_113 = 'b111111111;
    x_114 = 'b111111001;
    x_115 = 'b111100001;
    x_116 = 'b111011111;
    x_117 = 'b111010110;
    x_118 = 'b111010000;
    x_119 = 'b111101111;
    x_120 = 'b111110010;
    x_121 = 'b111100001;
    x_122 = 'b111000011;
    x_123 = 'b110110100;
    x_124 = 'b111101011;
    x_125 = 'b111001100;
    x_126 = 'b110100011;
    x_127 = 'b111000110;
    x_128 = 'b000001110;
    x_129 = 'b000001110;
    x_130 = 'b000001001;
    x_131 = 'b000001111;
    x_132 = 'b000010101;
    x_133 = 'b000001011;
    x_134 = 'b000000000;
    x_135 = 'b000000000;
    x_136 = 'b000000101;
    x_137 = 'b000001111;
    x_138 = 'b000011100;
    x_139 = 'b000001101;
    x_140 = 'b000001110;
    x_141 = 'b000001110;
    x_142 = 'b000000100;
    x_143 = 'b000000111;
    x_144 = 'b000001010;
    x_145 = 'b000001010;
    x_146 = 'b000000011;
    x_147 = 'b111111111;
    x_148 = 'b111111000;
    x_149 = 'b000000011;
    x_150 = 'b000000101;
    x_151 = 'b111111110;
    x_152 = 'b111111001;
    x_153 = 'b111111000;
    x_154 = 'b000000000;
    x_155 = 'b000000010;
    x_156 = 'b000000110;
    x_157 = 'b111111011;
    x_158 = 'b111111010;
    x_159 = 'b111111111;
    x_160 = 'b000001000;
    x_161 = 'b000001000;
    x_162 = 'b000000000;
    x_163 = 'b000000011;
    x_164 = 'b000000010;
    x_165 = 'b000000100;
    x_166 = 'b111111110;
    x_167 = 'b000011000;
    x_168 = 'b111111110;
    x_169 = 'b111100011;
    x_170 = 'b111100111;
    x_171 = 'b000000001;
    x_172 = 'b111100111;
    x_173 = 'b000000101;
    x_174 = 'b111110011;
    x_175 = 'b111111010;
    x_176 = 'b111110111;
    x_177 = 'b111111111;
    x_178 = 'b111111001;
    x_179 = 'b111100001;
    x_180 = 'b111011111;
    x_181 = 'b111010110;
    x_182 = 'b111010000;
    x_183 = 'b111101111;
    x_184 = 'b111110010;
    x_185 = 'b111100001;
    x_186 = 'b111000011;
    x_187 = 'b110110100;
    x_188 = 'b111101011;
    x_189 = 'b111001100;
    x_190 = 'b110100011;
    x_191 = 'b111000110;
    x_192 = 'b000001110;
    x_193 = 'b000001110;
    x_194 = 'b000001001;
    x_195 = 'b000001111;
    x_196 = 'b000010101;
    x_197 = 'b000001011;
    x_198 = 'b000000000;
    x_199 = 'b000000000;
    x_200 = 'b000000101;
    x_201 = 'b000001111;
    x_202 = 'b000011100;
    x_203 = 'b000001101;
    x_204 = 'b000001110;
    x_205 = 'b000001110;
    x_206 = 'b000000100;
    x_207 = 'b000000111;
    x_208 = 'b000001010;
    x_209 = 'b000001010;
    x_210 = 'b000000011;
    x_211 = 'b111111111;
    x_212 = 'b111111000;
    x_213 = 'b000000011;
    x_214 = 'b000000101;
    x_215 = 'b111111110;
    x_216 = 'b111111001;
    x_217 = 'b111111000;
    x_218 = 'b000000000;
    x_219 = 'b000000010;
    x_220 = 'b000000110;
    x_221 = 'b111111011;
    x_222 = 'b111111010;
    x_223 = 'b111111111;
    x_224 = 'b000001000;
    x_225 = 'b000001000;
    x_226 = 'b000000000;
    x_227 = 'b000000011;
    x_228 = 'b000000010;
    x_229 = 'b000000100;
    x_230 = 'b111111110;
    x_231 = 'b000011000;
    x_232 = 'b111111110;
    x_233 = 'b111100011;
    x_234 = 'b111100111;
    x_235 = 'b000000001;
    x_236 = 'b111100111;
    x_237 = 'b000000101;
    x_238 = 'b111110011;
    x_239 = 'b111111010;
    x_240 = 'b111110111;
    x_241 = 'b111111111;
    x_242 = 'b111111001;
    x_243 = 'b111100001;
    x_244 = 'b111011111;
    x_245 = 'b111010110;
    x_246 = 'b111010000;
    x_247 = 'b111101111;
    x_248 = 'b111110010;
    x_249 = 'b111100001;
    x_250 = 'b111000011;
    x_251 = 'b110110100;
    x_252 = 'b111101011;
    x_253 = 'b111001100;
    x_254 = 'b110100011;
    x_255 = 'b111000110;

    h_0 = 'b000001110;
    h_1 = 'b000001110;
    h_2 = 'b000001001;
    h_3 = 'b000001111;
    h_4 = 'b000010101;
    h_5 = 'b000001011;
    h_6 = 'b000000000;
    h_7 = 'b000000000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000001001;
    x_1 = 'b000010010;
    x_2 = 'b000010101;
    x_3 = 'b000011101;
    x_4 = 'b000011101;
    x_5 = 'b000010001;
    x_6 = 'b000001011;
    x_7 = 'b000000000;
    x_8 = 'b000001000;
    x_9 = 'b000011000;
    x_10 = 'b000100110;
    x_11 = 'b000001111;
    x_12 = 'b000001100;
    x_13 = 'b000001010;
    x_14 = 'b111111011;
    x_15 = 'b000001000;
    x_16 = 'b000001100;
    x_17 = 'b000001100;
    x_18 = 'b000000100;
    x_19 = 'b111111101;
    x_20 = 'b111110001;
    x_21 = 'b000000111;
    x_22 = 'b000001000;
    x_23 = 'b000000010;
    x_24 = 'b111111011;
    x_25 = 'b111111011;
    x_26 = 'b000000111;
    x_27 = 'b000000110;
    x_28 = 'b000001010;
    x_29 = 'b111111011;
    x_30 = 'b111111111;
    x_31 = 'b000000101;
    x_32 = 'b000010000;
    x_33 = 'b000010001;
    x_34 = 'b000001010;
    x_35 = 'b000001010;
    x_36 = 'b000000101;
    x_37 = 'b000000001;
    x_38 = 'b111111010;
    x_39 = 'b000011001;
    x_40 = 'b111110110;
    x_41 = 'b111111110;
    x_42 = 'b111110111;
    x_43 = 'b000011110;
    x_44 = 'b111110101;
    x_45 = 'b000000011;
    x_46 = 'b111110111;
    x_47 = 'b111111100;
    x_48 = 'b111111010;
    x_49 = 'b000000111;
    x_50 = 'b000000100;
    x_51 = 'b111101110;
    x_52 = 'b111101011;
    x_53 = 'b111100011;
    x_54 = 'b111011010;
    x_55 = 'b111110010;
    x_56 = 'b111110110;
    x_57 = 'b111101111;
    x_58 = 'b111010011;
    x_59 = 'b111000111;
    x_60 = 'b111011110;
    x_61 = 'b111000000;
    x_62 = 'b110010111;
    x_63 = 'b110111110;
    x_64 = 'b000001001;
    x_65 = 'b000010010;
    x_66 = 'b000010101;
    x_67 = 'b000011101;
    x_68 = 'b000011101;
    x_69 = 'b000010001;
    x_70 = 'b000001011;
    x_71 = 'b000000000;
    x_72 = 'b000001000;
    x_73 = 'b000011000;
    x_74 = 'b000100110;
    x_75 = 'b000001111;
    x_76 = 'b000001100;
    x_77 = 'b000001010;
    x_78 = 'b111111011;
    x_79 = 'b000001000;
    x_80 = 'b000001100;
    x_81 = 'b000001100;
    x_82 = 'b000000100;
    x_83 = 'b111111101;
    x_84 = 'b111110001;
    x_85 = 'b000000111;
    x_86 = 'b000001000;
    x_87 = 'b000000010;
    x_88 = 'b111111011;
    x_89 = 'b111111011;
    x_90 = 'b000000111;
    x_91 = 'b000000110;
    x_92 = 'b000001010;
    x_93 = 'b111111011;
    x_94 = 'b111111111;
    x_95 = 'b000000101;
    x_96 = 'b000010000;
    x_97 = 'b000010001;
    x_98 = 'b000001010;
    x_99 = 'b000001010;
    x_100 = 'b000000101;
    x_101 = 'b000000001;
    x_102 = 'b111111010;
    x_103 = 'b000011001;
    x_104 = 'b111110110;
    x_105 = 'b111111110;
    x_106 = 'b111110111;
    x_107 = 'b000011110;
    x_108 = 'b111110101;
    x_109 = 'b000000011;
    x_110 = 'b111110111;
    x_111 = 'b111111100;
    x_112 = 'b111111010;
    x_113 = 'b000000111;
    x_114 = 'b000000100;
    x_115 = 'b111101110;
    x_116 = 'b111101011;
    x_117 = 'b111100011;
    x_118 = 'b111011010;
    x_119 = 'b111110010;
    x_120 = 'b111110110;
    x_121 = 'b111101111;
    x_122 = 'b111010011;
    x_123 = 'b111000111;
    x_124 = 'b111011110;
    x_125 = 'b111000000;
    x_126 = 'b110010111;
    x_127 = 'b110111110;
    x_128 = 'b000001001;
    x_129 = 'b000010010;
    x_130 = 'b000010101;
    x_131 = 'b000011101;
    x_132 = 'b000011101;
    x_133 = 'b000010001;
    x_134 = 'b000001011;
    x_135 = 'b000000000;
    x_136 = 'b000001000;
    x_137 = 'b000011000;
    x_138 = 'b000100110;
    x_139 = 'b000001111;
    x_140 = 'b000001100;
    x_141 = 'b000001010;
    x_142 = 'b111111011;
    x_143 = 'b000001000;
    x_144 = 'b000001100;
    x_145 = 'b000001100;
    x_146 = 'b000000100;
    x_147 = 'b111111101;
    x_148 = 'b111110001;
    x_149 = 'b000000111;
    x_150 = 'b000001000;
    x_151 = 'b000000010;
    x_152 = 'b111111011;
    x_153 = 'b111111011;
    x_154 = 'b000000111;
    x_155 = 'b000000110;
    x_156 = 'b000001010;
    x_157 = 'b111111011;
    x_158 = 'b111111111;
    x_159 = 'b000000101;
    x_160 = 'b000010000;
    x_161 = 'b000010001;
    x_162 = 'b000001010;
    x_163 = 'b000001010;
    x_164 = 'b000000101;
    x_165 = 'b000000001;
    x_166 = 'b111111010;
    x_167 = 'b000011001;
    x_168 = 'b111110110;
    x_169 = 'b111111110;
    x_170 = 'b111110111;
    x_171 = 'b000011110;
    x_172 = 'b111110101;
    x_173 = 'b000000011;
    x_174 = 'b111110111;
    x_175 = 'b111111100;
    x_176 = 'b111111010;
    x_177 = 'b000000111;
    x_178 = 'b000000100;
    x_179 = 'b111101110;
    x_180 = 'b111101011;
    x_181 = 'b111100011;
    x_182 = 'b111011010;
    x_183 = 'b111110010;
    x_184 = 'b111110110;
    x_185 = 'b111101111;
    x_186 = 'b111010011;
    x_187 = 'b111000111;
    x_188 = 'b111011110;
    x_189 = 'b111000000;
    x_190 = 'b110010111;
    x_191 = 'b110111110;
    x_192 = 'b000001001;
    x_193 = 'b000010010;
    x_194 = 'b000010101;
    x_195 = 'b000011101;
    x_196 = 'b000011101;
    x_197 = 'b000010001;
    x_198 = 'b000001011;
    x_199 = 'b000000000;
    x_200 = 'b000001000;
    x_201 = 'b000011000;
    x_202 = 'b000100110;
    x_203 = 'b000001111;
    x_204 = 'b000001100;
    x_205 = 'b000001010;
    x_206 = 'b111111011;
    x_207 = 'b000001000;
    x_208 = 'b000001100;
    x_209 = 'b000001100;
    x_210 = 'b000000100;
    x_211 = 'b111111101;
    x_212 = 'b111110001;
    x_213 = 'b000000111;
    x_214 = 'b000001000;
    x_215 = 'b000000010;
    x_216 = 'b111111011;
    x_217 = 'b111111011;
    x_218 = 'b000000111;
    x_219 = 'b000000110;
    x_220 = 'b000001010;
    x_221 = 'b111111011;
    x_222 = 'b111111111;
    x_223 = 'b000000101;
    x_224 = 'b000010000;
    x_225 = 'b000010001;
    x_226 = 'b000001010;
    x_227 = 'b000001010;
    x_228 = 'b000000101;
    x_229 = 'b000000001;
    x_230 = 'b111111010;
    x_231 = 'b000011001;
    x_232 = 'b111110110;
    x_233 = 'b111111110;
    x_234 = 'b111110111;
    x_235 = 'b000011110;
    x_236 = 'b111110101;
    x_237 = 'b000000011;
    x_238 = 'b111110111;
    x_239 = 'b111111100;
    x_240 = 'b111111010;
    x_241 = 'b000000111;
    x_242 = 'b000000100;
    x_243 = 'b111101110;
    x_244 = 'b111101011;
    x_245 = 'b111100011;
    x_246 = 'b111011010;
    x_247 = 'b111110010;
    x_248 = 'b111110110;
    x_249 = 'b111101111;
    x_250 = 'b111010011;
    x_251 = 'b111000111;
    x_252 = 'b111011110;
    x_253 = 'b111000000;
    x_254 = 'b110010111;
    x_255 = 'b110111110;

    h_0 = 'b000001001;
    h_1 = 'b000010010;
    h_2 = 'b000010101;
    h_3 = 'b000011101;
    h_4 = 'b000011101;
    h_5 = 'b000010001;
    h_6 = 'b000001011;
    h_7 = 'b000000000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000001110;
    x_1 = 'b000011011;
    x_2 = 'b000011111;
    x_3 = 'b000100101;
    x_4 = 'b000100001;
    x_5 = 'b000010100;
    x_6 = 'b000001011;
    x_7 = 'b000000001;
    x_8 = 'b000010101;
    x_9 = 'b000100110;
    x_10 = 'b000110010;
    x_11 = 'b000010011;
    x_12 = 'b000010001;
    x_13 = 'b000010110;
    x_14 = 'b000000111;
    x_15 = 'b000010110;
    x_16 = 'b000011101;
    x_17 = 'b000011100;
    x_18 = 'b000010000;
    x_19 = 'b000000111;
    x_20 = 'b111111011;
    x_21 = 'b000001011;
    x_22 = 'b000001001;
    x_23 = 'b111111110;
    x_24 = 'b000000101;
    x_25 = 'b000000100;
    x_26 = 'b000000110;
    x_27 = 'b000000011;
    x_28 = 'b000000110;
    x_29 = 'b000010010;
    x_30 = 'b111111101;
    x_31 = 'b000000100;
    x_32 = 'b000010001;
    x_33 = 'b000001111;
    x_34 = 'b000001011;
    x_35 = 'b000001011;
    x_36 = 'b000000010;
    x_37 = 'b111110101;
    x_38 = 'b000001110;
    x_39 = 'b000011001;
    x_40 = 'b000010101;
    x_41 = 'b111111100;
    x_42 = 'b000010001;
    x_43 = 'b000001000;
    x_44 = 'b000000110;
    x_45 = 'b000000011;
    x_46 = 'b000000101;
    x_47 = 'b000001010;
    x_48 = 'b000000101;
    x_49 = 'b000010100;
    x_50 = 'b000010101;
    x_51 = 'b000000000;
    x_52 = 'b111111011;
    x_53 = 'b111110000;
    x_54 = 'b111100011;
    x_55 = 'b111111001;
    x_56 = 'b000000000;
    x_57 = 'b000000001;
    x_58 = 'b111101001;
    x_59 = 'b111011100;
    x_60 = 'b111100001;
    x_61 = 'b111001101;
    x_62 = 'b110100111;
    x_63 = 'b110111111;
    x_64 = 'b000001110;
    x_65 = 'b000011011;
    x_66 = 'b000011111;
    x_67 = 'b000100101;
    x_68 = 'b000100001;
    x_69 = 'b000010100;
    x_70 = 'b000001011;
    x_71 = 'b000000001;
    x_72 = 'b000010101;
    x_73 = 'b000100110;
    x_74 = 'b000110010;
    x_75 = 'b000010011;
    x_76 = 'b000010001;
    x_77 = 'b000010110;
    x_78 = 'b000000111;
    x_79 = 'b000010110;
    x_80 = 'b000011101;
    x_81 = 'b000011100;
    x_82 = 'b000010000;
    x_83 = 'b000000111;
    x_84 = 'b111111011;
    x_85 = 'b000001011;
    x_86 = 'b000001001;
    x_87 = 'b111111110;
    x_88 = 'b000000101;
    x_89 = 'b000000100;
    x_90 = 'b000000110;
    x_91 = 'b000000011;
    x_92 = 'b000000110;
    x_93 = 'b000010010;
    x_94 = 'b111111101;
    x_95 = 'b000000100;
    x_96 = 'b000010001;
    x_97 = 'b000001111;
    x_98 = 'b000001011;
    x_99 = 'b000001011;
    x_100 = 'b000000010;
    x_101 = 'b111110101;
    x_102 = 'b000001110;
    x_103 = 'b000011001;
    x_104 = 'b000010101;
    x_105 = 'b111111100;
    x_106 = 'b000010001;
    x_107 = 'b000001000;
    x_108 = 'b000000110;
    x_109 = 'b000000011;
    x_110 = 'b000000101;
    x_111 = 'b000001010;
    x_112 = 'b000000101;
    x_113 = 'b000010100;
    x_114 = 'b000010101;
    x_115 = 'b000000000;
    x_116 = 'b111111011;
    x_117 = 'b111110000;
    x_118 = 'b111100011;
    x_119 = 'b111111001;
    x_120 = 'b000000000;
    x_121 = 'b000000001;
    x_122 = 'b111101001;
    x_123 = 'b111011100;
    x_124 = 'b111100001;
    x_125 = 'b111001101;
    x_126 = 'b110100111;
    x_127 = 'b110111111;
    x_128 = 'b000001110;
    x_129 = 'b000011011;
    x_130 = 'b000011111;
    x_131 = 'b000100101;
    x_132 = 'b000100001;
    x_133 = 'b000010100;
    x_134 = 'b000001011;
    x_135 = 'b000000001;
    x_136 = 'b000010101;
    x_137 = 'b000100110;
    x_138 = 'b000110010;
    x_139 = 'b000010011;
    x_140 = 'b000010001;
    x_141 = 'b000010110;
    x_142 = 'b000000111;
    x_143 = 'b000010110;
    x_144 = 'b000011101;
    x_145 = 'b000011100;
    x_146 = 'b000010000;
    x_147 = 'b000000111;
    x_148 = 'b111111011;
    x_149 = 'b000001011;
    x_150 = 'b000001001;
    x_151 = 'b111111110;
    x_152 = 'b000000101;
    x_153 = 'b000000100;
    x_154 = 'b000000110;
    x_155 = 'b000000011;
    x_156 = 'b000000110;
    x_157 = 'b000010010;
    x_158 = 'b111111101;
    x_159 = 'b000000100;
    x_160 = 'b000010001;
    x_161 = 'b000001111;
    x_162 = 'b000001011;
    x_163 = 'b000001011;
    x_164 = 'b000000010;
    x_165 = 'b111110101;
    x_166 = 'b000001110;
    x_167 = 'b000011001;
    x_168 = 'b000010101;
    x_169 = 'b111111100;
    x_170 = 'b000010001;
    x_171 = 'b000001000;
    x_172 = 'b000000110;
    x_173 = 'b000000011;
    x_174 = 'b000000101;
    x_175 = 'b000001010;
    x_176 = 'b000000101;
    x_177 = 'b000010100;
    x_178 = 'b000010101;
    x_179 = 'b000000000;
    x_180 = 'b111111011;
    x_181 = 'b111110000;
    x_182 = 'b111100011;
    x_183 = 'b111111001;
    x_184 = 'b000000000;
    x_185 = 'b000000001;
    x_186 = 'b111101001;
    x_187 = 'b111011100;
    x_188 = 'b111100001;
    x_189 = 'b111001101;
    x_190 = 'b110100111;
    x_191 = 'b110111111;
    x_192 = 'b000001110;
    x_193 = 'b000011011;
    x_194 = 'b000011111;
    x_195 = 'b000100101;
    x_196 = 'b000100001;
    x_197 = 'b000010100;
    x_198 = 'b000001011;
    x_199 = 'b000000001;
    x_200 = 'b000010101;
    x_201 = 'b000100110;
    x_202 = 'b000110010;
    x_203 = 'b000010011;
    x_204 = 'b000010001;
    x_205 = 'b000010110;
    x_206 = 'b000000111;
    x_207 = 'b000010110;
    x_208 = 'b000011101;
    x_209 = 'b000011100;
    x_210 = 'b000010000;
    x_211 = 'b000000111;
    x_212 = 'b111111011;
    x_213 = 'b000001011;
    x_214 = 'b000001001;
    x_215 = 'b111111110;
    x_216 = 'b000000101;
    x_217 = 'b000000100;
    x_218 = 'b000000110;
    x_219 = 'b000000011;
    x_220 = 'b000000110;
    x_221 = 'b000010010;
    x_222 = 'b111111101;
    x_223 = 'b000000100;
    x_224 = 'b000010001;
    x_225 = 'b000001111;
    x_226 = 'b000001011;
    x_227 = 'b000001011;
    x_228 = 'b000000010;
    x_229 = 'b111110101;
    x_230 = 'b000001110;
    x_231 = 'b000011001;
    x_232 = 'b000010101;
    x_233 = 'b111111100;
    x_234 = 'b000010001;
    x_235 = 'b000001000;
    x_236 = 'b000000110;
    x_237 = 'b000000011;
    x_238 = 'b000000101;
    x_239 = 'b000001010;
    x_240 = 'b000000101;
    x_241 = 'b000010100;
    x_242 = 'b000010101;
    x_243 = 'b000000000;
    x_244 = 'b111111011;
    x_245 = 'b111110000;
    x_246 = 'b111100011;
    x_247 = 'b111111001;
    x_248 = 'b000000000;
    x_249 = 'b000000001;
    x_250 = 'b111101001;
    x_251 = 'b111011100;
    x_252 = 'b111100001;
    x_253 = 'b111001101;
    x_254 = 'b110100111;
    x_255 = 'b110111111;

    h_0 = 'b000001110;
    h_1 = 'b000011011;
    h_2 = 'b000011111;
    h_3 = 'b000100101;
    h_4 = 'b000100001;
    h_5 = 'b000010100;
    h_6 = 'b000001011;
    h_7 = 'b000000001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000011010;
    x_1 = 'b000100110;
    x_2 = 'b000100111;
    x_3 = 'b000101011;
    x_4 = 'b000100111;
    x_5 = 'b000011011;
    x_6 = 'b000010010;
    x_7 = 'b000010110;
    x_8 = 'b000100111;
    x_9 = 'b000110101;
    x_10 = 'b001000010;
    x_11 = 'b000100110;
    x_12 = 'b000011101;
    x_13 = 'b000011100;
    x_14 = 'b000100000;
    x_15 = 'b000101101;
    x_16 = 'b000110011;
    x_17 = 'b000110001;
    x_18 = 'b000100111;
    x_19 = 'b000011110;
    x_20 = 'b000001100;
    x_21 = 'b000010011;
    x_22 = 'b000010000;
    x_23 = 'b000000110;
    x_24 = 'b000001100;
    x_25 = 'b000001011;
    x_26 = 'b000001111;
    x_27 = 'b000001111;
    x_28 = 'b000001111;
    x_29 = 'b000011001;
    x_30 = 'b000000101;
    x_31 = 'b000010001;
    x_32 = 'b000011100;
    x_33 = 'b000011010;
    x_34 = 'b000010101;
    x_35 = 'b000010111;
    x_36 = 'b000010001;
    x_37 = 'b000000001;
    x_38 = 'b000011101;
    x_39 = 'b000100001;
    x_40 = 'b000101110;
    x_41 = 'b000000011;
    x_42 = 'b000010010;
    x_43 = 'b111111001;
    x_44 = 'b000011111;
    x_45 = 'b000011001;
    x_46 = 'b000011100;
    x_47 = 'b000100011;
    x_48 = 'b000011101;
    x_49 = 'b000101010;
    x_50 = 'b000101100;
    x_51 = 'b000100000;
    x_52 = 'b000011011;
    x_53 = 'b000001110;
    x_54 = 'b000000011;
    x_55 = 'b000001110;
    x_56 = 'b000010101;
    x_57 = 'b000011001;
    x_58 = 'b000001010;
    x_59 = 'b111111101;
    x_60 = 'b111110111;
    x_61 = 'b111101011;
    x_62 = 'b111001110;
    x_63 = 'b111001111;
    x_64 = 'b000011010;
    x_65 = 'b000100110;
    x_66 = 'b000100111;
    x_67 = 'b000101011;
    x_68 = 'b000100111;
    x_69 = 'b000011011;
    x_70 = 'b000010010;
    x_71 = 'b000010110;
    x_72 = 'b000100111;
    x_73 = 'b000110101;
    x_74 = 'b001000010;
    x_75 = 'b000100110;
    x_76 = 'b000011101;
    x_77 = 'b000011100;
    x_78 = 'b000100000;
    x_79 = 'b000101101;
    x_80 = 'b000110011;
    x_81 = 'b000110001;
    x_82 = 'b000100111;
    x_83 = 'b000011110;
    x_84 = 'b000001100;
    x_85 = 'b000010011;
    x_86 = 'b000010000;
    x_87 = 'b000000110;
    x_88 = 'b000001100;
    x_89 = 'b000001011;
    x_90 = 'b000001111;
    x_91 = 'b000001111;
    x_92 = 'b000001111;
    x_93 = 'b000011001;
    x_94 = 'b000000101;
    x_95 = 'b000010001;
    x_96 = 'b000011100;
    x_97 = 'b000011010;
    x_98 = 'b000010101;
    x_99 = 'b000010111;
    x_100 = 'b000010001;
    x_101 = 'b000000001;
    x_102 = 'b000011101;
    x_103 = 'b000100001;
    x_104 = 'b000101110;
    x_105 = 'b000000011;
    x_106 = 'b000010010;
    x_107 = 'b111111001;
    x_108 = 'b000011111;
    x_109 = 'b000011001;
    x_110 = 'b000011100;
    x_111 = 'b000100011;
    x_112 = 'b000011101;
    x_113 = 'b000101010;
    x_114 = 'b000101100;
    x_115 = 'b000100000;
    x_116 = 'b000011011;
    x_117 = 'b000001110;
    x_118 = 'b000000011;
    x_119 = 'b000001110;
    x_120 = 'b000010101;
    x_121 = 'b000011001;
    x_122 = 'b000001010;
    x_123 = 'b111111101;
    x_124 = 'b111110111;
    x_125 = 'b111101011;
    x_126 = 'b111001110;
    x_127 = 'b111001111;
    x_128 = 'b000011010;
    x_129 = 'b000100110;
    x_130 = 'b000100111;
    x_131 = 'b000101011;
    x_132 = 'b000100111;
    x_133 = 'b000011011;
    x_134 = 'b000010010;
    x_135 = 'b000010110;
    x_136 = 'b000100111;
    x_137 = 'b000110101;
    x_138 = 'b001000010;
    x_139 = 'b000100110;
    x_140 = 'b000011101;
    x_141 = 'b000011100;
    x_142 = 'b000100000;
    x_143 = 'b000101101;
    x_144 = 'b000110011;
    x_145 = 'b000110001;
    x_146 = 'b000100111;
    x_147 = 'b000011110;
    x_148 = 'b000001100;
    x_149 = 'b000010011;
    x_150 = 'b000010000;
    x_151 = 'b000000110;
    x_152 = 'b000001100;
    x_153 = 'b000001011;
    x_154 = 'b000001111;
    x_155 = 'b000001111;
    x_156 = 'b000001111;
    x_157 = 'b000011001;
    x_158 = 'b000000101;
    x_159 = 'b000010001;
    x_160 = 'b000011100;
    x_161 = 'b000011010;
    x_162 = 'b000010101;
    x_163 = 'b000010111;
    x_164 = 'b000010001;
    x_165 = 'b000000001;
    x_166 = 'b000011101;
    x_167 = 'b000100001;
    x_168 = 'b000101110;
    x_169 = 'b000000011;
    x_170 = 'b000010010;
    x_171 = 'b111111001;
    x_172 = 'b000011111;
    x_173 = 'b000011001;
    x_174 = 'b000011100;
    x_175 = 'b000100011;
    x_176 = 'b000011101;
    x_177 = 'b000101010;
    x_178 = 'b000101100;
    x_179 = 'b000100000;
    x_180 = 'b000011011;
    x_181 = 'b000001110;
    x_182 = 'b000000011;
    x_183 = 'b000001110;
    x_184 = 'b000010101;
    x_185 = 'b000011001;
    x_186 = 'b000001010;
    x_187 = 'b111111101;
    x_188 = 'b111110111;
    x_189 = 'b111101011;
    x_190 = 'b111001110;
    x_191 = 'b111001111;
    x_192 = 'b000011010;
    x_193 = 'b000100110;
    x_194 = 'b000100111;
    x_195 = 'b000101011;
    x_196 = 'b000100111;
    x_197 = 'b000011011;
    x_198 = 'b000010010;
    x_199 = 'b000010110;
    x_200 = 'b000100111;
    x_201 = 'b000110101;
    x_202 = 'b001000010;
    x_203 = 'b000100110;
    x_204 = 'b000011101;
    x_205 = 'b000011100;
    x_206 = 'b000100000;
    x_207 = 'b000101101;
    x_208 = 'b000110011;
    x_209 = 'b000110001;
    x_210 = 'b000100111;
    x_211 = 'b000011110;
    x_212 = 'b000001100;
    x_213 = 'b000010011;
    x_214 = 'b000010000;
    x_215 = 'b000000110;
    x_216 = 'b000001100;
    x_217 = 'b000001011;
    x_218 = 'b000001111;
    x_219 = 'b000001111;
    x_220 = 'b000001111;
    x_221 = 'b000011001;
    x_222 = 'b000000101;
    x_223 = 'b000010001;
    x_224 = 'b000011100;
    x_225 = 'b000011010;
    x_226 = 'b000010101;
    x_227 = 'b000010111;
    x_228 = 'b000010001;
    x_229 = 'b000000001;
    x_230 = 'b000011101;
    x_231 = 'b000100001;
    x_232 = 'b000101110;
    x_233 = 'b000000011;
    x_234 = 'b000010010;
    x_235 = 'b111111001;
    x_236 = 'b000011111;
    x_237 = 'b000011001;
    x_238 = 'b000011100;
    x_239 = 'b000100011;
    x_240 = 'b000011101;
    x_241 = 'b000101010;
    x_242 = 'b000101100;
    x_243 = 'b000100000;
    x_244 = 'b000011011;
    x_245 = 'b000001110;
    x_246 = 'b000000011;
    x_247 = 'b000001110;
    x_248 = 'b000010101;
    x_249 = 'b000011001;
    x_250 = 'b000001010;
    x_251 = 'b111111101;
    x_252 = 'b111110111;
    x_253 = 'b111101011;
    x_254 = 'b111001110;
    x_255 = 'b111001111;

    h_0 = 'b000011010;
    h_1 = 'b000100110;
    h_2 = 'b000100111;
    h_3 = 'b000101011;
    h_4 = 'b000100111;
    h_5 = 'b000011011;
    h_6 = 'b000010010;
    h_7 = 'b000010110;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000100100;
    x_1 = 'b000101111;
    x_2 = 'b000101111;
    x_3 = 'b000110001;
    x_4 = 'b000101110;
    x_5 = 'b000100010;
    x_6 = 'b000011000;
    x_7 = 'b000100001;
    x_8 = 'b000110000;
    x_9 = 'b000111001;
    x_10 = 'b001000001;
    x_11 = 'b000101110;
    x_12 = 'b000101000;
    x_13 = 'b000100111;
    x_14 = 'b000101000;
    x_15 = 'b000110001;
    x_16 = 'b000110101;
    x_17 = 'b000110000;
    x_18 = 'b000101101;
    x_19 = 'b000101011;
    x_20 = 'b000011010;
    x_21 = 'b000001101;
    x_22 = 'b000001010;
    x_23 = 'b111111101;
    x_24 = 'b000000010;
    x_25 = 'b000000010;
    x_26 = 'b000000111;
    x_27 = 'b000000100;
    x_28 = 'b111111110;
    x_29 = 'b000001100;
    x_30 = 'b000000000;
    x_31 = 'b000000111;
    x_32 = 'b000010010;
    x_33 = 'b000001111;
    x_34 = 'b000001000;
    x_35 = 'b000001001;
    x_36 = 'b111111101;
    x_37 = 'b111110100;
    x_38 = 'b000010010;
    x_39 = 'b000010101;
    x_40 = 'b000011101;
    x_41 = 'b111111000;
    x_42 = 'b000000001;
    x_43 = 'b111011111;
    x_44 = 'b000001110;
    x_45 = 'b000010010;
    x_46 = 'b000010110;
    x_47 = 'b000011100;
    x_48 = 'b000010100;
    x_49 = 'b000100000;
    x_50 = 'b000011111;
    x_51 = 'b000011110;
    x_52 = 'b000011010;
    x_53 = 'b000010001;
    x_54 = 'b000000100;
    x_55 = 'b000001100;
    x_56 = 'b000001111;
    x_57 = 'b000011000;
    x_58 = 'b000010010;
    x_59 = 'b000001010;
    x_60 = 'b000001010;
    x_61 = 'b000000101;
    x_62 = 'b111110010;
    x_63 = 'b111100011;
    x_64 = 'b000100100;
    x_65 = 'b000101111;
    x_66 = 'b000101111;
    x_67 = 'b000110001;
    x_68 = 'b000101110;
    x_69 = 'b000100010;
    x_70 = 'b000011000;
    x_71 = 'b000100001;
    x_72 = 'b000110000;
    x_73 = 'b000111001;
    x_74 = 'b001000001;
    x_75 = 'b000101110;
    x_76 = 'b000101000;
    x_77 = 'b000100111;
    x_78 = 'b000101000;
    x_79 = 'b000110001;
    x_80 = 'b000110101;
    x_81 = 'b000110000;
    x_82 = 'b000101101;
    x_83 = 'b000101011;
    x_84 = 'b000011010;
    x_85 = 'b000001101;
    x_86 = 'b000001010;
    x_87 = 'b111111101;
    x_88 = 'b000000010;
    x_89 = 'b000000010;
    x_90 = 'b000000111;
    x_91 = 'b000000100;
    x_92 = 'b111111110;
    x_93 = 'b000001100;
    x_94 = 'b000000000;
    x_95 = 'b000000111;
    x_96 = 'b000010010;
    x_97 = 'b000001111;
    x_98 = 'b000001000;
    x_99 = 'b000001001;
    x_100 = 'b111111101;
    x_101 = 'b111110100;
    x_102 = 'b000010010;
    x_103 = 'b000010101;
    x_104 = 'b000011101;
    x_105 = 'b111111000;
    x_106 = 'b000000001;
    x_107 = 'b111011111;
    x_108 = 'b000001110;
    x_109 = 'b000010010;
    x_110 = 'b000010110;
    x_111 = 'b000011100;
    x_112 = 'b000010100;
    x_113 = 'b000100000;
    x_114 = 'b000011111;
    x_115 = 'b000011110;
    x_116 = 'b000011010;
    x_117 = 'b000010001;
    x_118 = 'b000000100;
    x_119 = 'b000001100;
    x_120 = 'b000001111;
    x_121 = 'b000011000;
    x_122 = 'b000010010;
    x_123 = 'b000001010;
    x_124 = 'b000001010;
    x_125 = 'b000000101;
    x_126 = 'b111110010;
    x_127 = 'b111100011;
    x_128 = 'b000100100;
    x_129 = 'b000101111;
    x_130 = 'b000101111;
    x_131 = 'b000110001;
    x_132 = 'b000101110;
    x_133 = 'b000100010;
    x_134 = 'b000011000;
    x_135 = 'b000100001;
    x_136 = 'b000110000;
    x_137 = 'b000111001;
    x_138 = 'b001000001;
    x_139 = 'b000101110;
    x_140 = 'b000101000;
    x_141 = 'b000100111;
    x_142 = 'b000101000;
    x_143 = 'b000110001;
    x_144 = 'b000110101;
    x_145 = 'b000110000;
    x_146 = 'b000101101;
    x_147 = 'b000101011;
    x_148 = 'b000011010;
    x_149 = 'b000001101;
    x_150 = 'b000001010;
    x_151 = 'b111111101;
    x_152 = 'b000000010;
    x_153 = 'b000000010;
    x_154 = 'b000000111;
    x_155 = 'b000000100;
    x_156 = 'b111111110;
    x_157 = 'b000001100;
    x_158 = 'b000000000;
    x_159 = 'b000000111;
    x_160 = 'b000010010;
    x_161 = 'b000001111;
    x_162 = 'b000001000;
    x_163 = 'b000001001;
    x_164 = 'b111111101;
    x_165 = 'b111110100;
    x_166 = 'b000010010;
    x_167 = 'b000010101;
    x_168 = 'b000011101;
    x_169 = 'b111111000;
    x_170 = 'b000000001;
    x_171 = 'b111011111;
    x_172 = 'b000001110;
    x_173 = 'b000010010;
    x_174 = 'b000010110;
    x_175 = 'b000011100;
    x_176 = 'b000010100;
    x_177 = 'b000100000;
    x_178 = 'b000011111;
    x_179 = 'b000011110;
    x_180 = 'b000011010;
    x_181 = 'b000010001;
    x_182 = 'b000000100;
    x_183 = 'b000001100;
    x_184 = 'b000001111;
    x_185 = 'b000011000;
    x_186 = 'b000010010;
    x_187 = 'b000001010;
    x_188 = 'b000001010;
    x_189 = 'b000000101;
    x_190 = 'b111110010;
    x_191 = 'b111100011;
    x_192 = 'b000100100;
    x_193 = 'b000101111;
    x_194 = 'b000101111;
    x_195 = 'b000110001;
    x_196 = 'b000101110;
    x_197 = 'b000100010;
    x_198 = 'b000011000;
    x_199 = 'b000100001;
    x_200 = 'b000110000;
    x_201 = 'b000111001;
    x_202 = 'b001000001;
    x_203 = 'b000101110;
    x_204 = 'b000101000;
    x_205 = 'b000100111;
    x_206 = 'b000101000;
    x_207 = 'b000110001;
    x_208 = 'b000110101;
    x_209 = 'b000110000;
    x_210 = 'b000101101;
    x_211 = 'b000101011;
    x_212 = 'b000011010;
    x_213 = 'b000001101;
    x_214 = 'b000001010;
    x_215 = 'b111111101;
    x_216 = 'b000000010;
    x_217 = 'b000000010;
    x_218 = 'b000000111;
    x_219 = 'b000000100;
    x_220 = 'b111111110;
    x_221 = 'b000001100;
    x_222 = 'b000000000;
    x_223 = 'b000000111;
    x_224 = 'b000010010;
    x_225 = 'b000001111;
    x_226 = 'b000001000;
    x_227 = 'b000001001;
    x_228 = 'b111111101;
    x_229 = 'b111110100;
    x_230 = 'b000010010;
    x_231 = 'b000010101;
    x_232 = 'b000011101;
    x_233 = 'b111111000;
    x_234 = 'b000000001;
    x_235 = 'b111011111;
    x_236 = 'b000001110;
    x_237 = 'b000010010;
    x_238 = 'b000010110;
    x_239 = 'b000011100;
    x_240 = 'b000010100;
    x_241 = 'b000100000;
    x_242 = 'b000011111;
    x_243 = 'b000011110;
    x_244 = 'b000011010;
    x_245 = 'b000010001;
    x_246 = 'b000000100;
    x_247 = 'b000001100;
    x_248 = 'b000001111;
    x_249 = 'b000011000;
    x_250 = 'b000010010;
    x_251 = 'b000001010;
    x_252 = 'b000001010;
    x_253 = 'b000000101;
    x_254 = 'b111110010;
    x_255 = 'b111100011;

    h_0 = 'b000100100;
    h_1 = 'b000101111;
    h_2 = 'b000101111;
    h_3 = 'b000110001;
    h_4 = 'b000101110;
    h_5 = 'b000100010;
    h_6 = 'b000011000;
    h_7 = 'b000100001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000010010;
    x_1 = 'b000011010;
    x_2 = 'b000010110;
    x_3 = 'b000010101;
    x_4 = 'b000010001;
    x_5 = 'b000000011;
    x_6 = 'b111110100;
    x_7 = 'b000001111;
    x_8 = 'b000011101;
    x_9 = 'b000100000;
    x_10 = 'b000100111;
    x_11 = 'b000010110;
    x_12 = 'b000010100;
    x_13 = 'b000001101;
    x_14 = 'b000011000;
    x_15 = 'b000100001;
    x_16 = 'b000100011;
    x_17 = 'b000011110;
    x_18 = 'b000011111;
    x_19 = 'b000011111;
    x_20 = 'b000010001;
    x_21 = 'b111111011;
    x_22 = 'b111111010;
    x_23 = 'b111110001;
    x_24 = 'b111110010;
    x_25 = 'b111110010;
    x_26 = 'b111110010;
    x_27 = 'b111110001;
    x_28 = 'b111111100;
    x_29 = 'b111111100;
    x_30 = 'b111110010;
    x_31 = 'b111101111;
    x_32 = 'b111111111;
    x_33 = 'b111110111;
    x_34 = 'b111101111;
    x_35 = 'b111110011;
    x_36 = 'b111100111;
    x_37 = 'b111101010;
    x_38 = 'b000000000;
    x_39 = 'b000000000;
    x_40 = 'b000000111;
    x_41 = 'b111010111;
    x_42 = 'b000000001;
    x_43 = 'b000010110;
    x_44 = 'b000000111;
    x_45 = 'b000011010;
    x_46 = 'b000011011;
    x_47 = 'b000011100;
    x_48 = 'b000011000;
    x_49 = 'b000100101;
    x_50 = 'b000100011;
    x_51 = 'b000101000;
    x_52 = 'b000100101;
    x_53 = 'b000100000;
    x_54 = 'b000011001;
    x_55 = 'b000011001;
    x_56 = 'b000011101;
    x_57 = 'b000101000;
    x_58 = 'b000100111;
    x_59 = 'b000100101;
    x_60 = 'b000011011;
    x_61 = 'b000011110;
    x_62 = 'b000001101;
    x_63 = 'b111111110;
    x_64 = 'b000010010;
    x_65 = 'b000011010;
    x_66 = 'b000010110;
    x_67 = 'b000010101;
    x_68 = 'b000010001;
    x_69 = 'b000000011;
    x_70 = 'b111110100;
    x_71 = 'b000001111;
    x_72 = 'b000011101;
    x_73 = 'b000100000;
    x_74 = 'b000100111;
    x_75 = 'b000010110;
    x_76 = 'b000010100;
    x_77 = 'b000001101;
    x_78 = 'b000011000;
    x_79 = 'b000100001;
    x_80 = 'b000100011;
    x_81 = 'b000011110;
    x_82 = 'b000011111;
    x_83 = 'b000011111;
    x_84 = 'b000010001;
    x_85 = 'b111111011;
    x_86 = 'b111111010;
    x_87 = 'b111110001;
    x_88 = 'b111110010;
    x_89 = 'b111110010;
    x_90 = 'b111110010;
    x_91 = 'b111110001;
    x_92 = 'b111111100;
    x_93 = 'b111111100;
    x_94 = 'b111110010;
    x_95 = 'b111101111;
    x_96 = 'b111111111;
    x_97 = 'b111110111;
    x_98 = 'b111101111;
    x_99 = 'b111110011;
    x_100 = 'b111100111;
    x_101 = 'b111101010;
    x_102 = 'b000000000;
    x_103 = 'b000000000;
    x_104 = 'b000000111;
    x_105 = 'b111010111;
    x_106 = 'b000000001;
    x_107 = 'b000010110;
    x_108 = 'b000000111;
    x_109 = 'b000011010;
    x_110 = 'b000011011;
    x_111 = 'b000011100;
    x_112 = 'b000011000;
    x_113 = 'b000100101;
    x_114 = 'b000100011;
    x_115 = 'b000101000;
    x_116 = 'b000100101;
    x_117 = 'b000100000;
    x_118 = 'b000011001;
    x_119 = 'b000011001;
    x_120 = 'b000011101;
    x_121 = 'b000101000;
    x_122 = 'b000100111;
    x_123 = 'b000100101;
    x_124 = 'b000011011;
    x_125 = 'b000011110;
    x_126 = 'b000001101;
    x_127 = 'b111111110;
    x_128 = 'b000010010;
    x_129 = 'b000011010;
    x_130 = 'b000010110;
    x_131 = 'b000010101;
    x_132 = 'b000010001;
    x_133 = 'b000000011;
    x_134 = 'b111110100;
    x_135 = 'b000001111;
    x_136 = 'b000011101;
    x_137 = 'b000100000;
    x_138 = 'b000100111;
    x_139 = 'b000010110;
    x_140 = 'b000010100;
    x_141 = 'b000001101;
    x_142 = 'b000011000;
    x_143 = 'b000100001;
    x_144 = 'b000100011;
    x_145 = 'b000011110;
    x_146 = 'b000011111;
    x_147 = 'b000011111;
    x_148 = 'b000010001;
    x_149 = 'b111111011;
    x_150 = 'b111111010;
    x_151 = 'b111110001;
    x_152 = 'b111110010;
    x_153 = 'b111110010;
    x_154 = 'b111110010;
    x_155 = 'b111110001;
    x_156 = 'b111111100;
    x_157 = 'b111111100;
    x_158 = 'b111110010;
    x_159 = 'b111101111;
    x_160 = 'b111111111;
    x_161 = 'b111110111;
    x_162 = 'b111101111;
    x_163 = 'b111110011;
    x_164 = 'b111100111;
    x_165 = 'b111101010;
    x_166 = 'b000000000;
    x_167 = 'b000000000;
    x_168 = 'b000000111;
    x_169 = 'b111010111;
    x_170 = 'b000000001;
    x_171 = 'b000010110;
    x_172 = 'b000000111;
    x_173 = 'b000011010;
    x_174 = 'b000011011;
    x_175 = 'b000011100;
    x_176 = 'b000011000;
    x_177 = 'b000100101;
    x_178 = 'b000100011;
    x_179 = 'b000101000;
    x_180 = 'b000100101;
    x_181 = 'b000100000;
    x_182 = 'b000011001;
    x_183 = 'b000011001;
    x_184 = 'b000011101;
    x_185 = 'b000101000;
    x_186 = 'b000100111;
    x_187 = 'b000100101;
    x_188 = 'b000011011;
    x_189 = 'b000011110;
    x_190 = 'b000001101;
    x_191 = 'b111111110;
    x_192 = 'b000010010;
    x_193 = 'b000011010;
    x_194 = 'b000010110;
    x_195 = 'b000010101;
    x_196 = 'b000010001;
    x_197 = 'b000000011;
    x_198 = 'b111110100;
    x_199 = 'b000001111;
    x_200 = 'b000011101;
    x_201 = 'b000100000;
    x_202 = 'b000100111;
    x_203 = 'b000010110;
    x_204 = 'b000010100;
    x_205 = 'b000001101;
    x_206 = 'b000011000;
    x_207 = 'b000100001;
    x_208 = 'b000100011;
    x_209 = 'b000011110;
    x_210 = 'b000011111;
    x_211 = 'b000011111;
    x_212 = 'b000010001;
    x_213 = 'b111111011;
    x_214 = 'b111111010;
    x_215 = 'b111110001;
    x_216 = 'b111110010;
    x_217 = 'b111110010;
    x_218 = 'b111110010;
    x_219 = 'b111110001;
    x_220 = 'b111111100;
    x_221 = 'b111111100;
    x_222 = 'b111110010;
    x_223 = 'b111101111;
    x_224 = 'b111111111;
    x_225 = 'b111110111;
    x_226 = 'b111101111;
    x_227 = 'b111110011;
    x_228 = 'b111100111;
    x_229 = 'b111101010;
    x_230 = 'b000000000;
    x_231 = 'b000000000;
    x_232 = 'b000000111;
    x_233 = 'b111010111;
    x_234 = 'b000000001;
    x_235 = 'b000010110;
    x_236 = 'b000000111;
    x_237 = 'b000011010;
    x_238 = 'b000011011;
    x_239 = 'b000011100;
    x_240 = 'b000011000;
    x_241 = 'b000100101;
    x_242 = 'b000100011;
    x_243 = 'b000101000;
    x_244 = 'b000100101;
    x_245 = 'b000100000;
    x_246 = 'b000011001;
    x_247 = 'b000011001;
    x_248 = 'b000011101;
    x_249 = 'b000101000;
    x_250 = 'b000100111;
    x_251 = 'b000100101;
    x_252 = 'b000011011;
    x_253 = 'b000011110;
    x_254 = 'b000001101;
    x_255 = 'b111111110;

    h_0 = 'b000010010;
    h_1 = 'b000011010;
    h_2 = 'b000010110;
    h_3 = 'b000010101;
    h_4 = 'b000010001;
    h_5 = 'b000000011;
    h_6 = 'b111110100;
    h_7 = 'b000001111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000001001;
    x_1 = 'b000010000;
    x_2 = 'b000001011;
    x_3 = 'b000001011;
    x_4 = 'b000000110;
    x_5 = 'b111111001;
    x_6 = 'b111101110;
    x_7 = 'b000001001;
    x_8 = 'b000010100;
    x_9 = 'b000011010;
    x_10 = 'b000100100;
    x_11 = 'b000010011;
    x_12 = 'b000010010;
    x_13 = 'b000001010;
    x_14 = 'b000010101;
    x_15 = 'b000011110;
    x_16 = 'b000100000;
    x_17 = 'b000100001;
    x_18 = 'b000100011;
    x_19 = 'b000100100;
    x_20 = 'b000010111;
    x_21 = 'b111110111;
    x_22 = 'b111110100;
    x_23 = 'b111101100;
    x_24 = 'b111101111;
    x_25 = 'b111110000;
    x_26 = 'b111101011;
    x_27 = 'b111101100;
    x_28 = 'b111111011;
    x_29 = 'b111111101;
    x_30 = 'b111110001;
    x_31 = 'b111101110;
    x_32 = 'b111111010;
    x_33 = 'b111110100;
    x_34 = 'b111101011;
    x_35 = 'b111101101;
    x_36 = 'b111100110;
    x_37 = 'b111100111;
    x_38 = 'b111111111;
    x_39 = 'b111110111;
    x_40 = 'b000001000;
    x_41 = 'b111001111;
    x_42 = 'b000001000;
    x_43 = 'b000011110;
    x_44 = 'b111111101;
    x_45 = 'b000101001;
    x_46 = 'b000010010;
    x_47 = 'b000011001;
    x_48 = 'b000010110;
    x_49 = 'b000100110;
    x_50 = 'b000101000;
    x_51 = 'b000101101;
    x_52 = 'b000101001;
    x_53 = 'b000100111;
    x_54 = 'b000100110;
    x_55 = 'b000011101;
    x_56 = 'b000011110;
    x_57 = 'b000110000;
    x_58 = 'b000101110;
    x_59 = 'b000110000;
    x_60 = 'b000101001;
    x_61 = 'b000110011;
    x_62 = 'b000011111;
    x_63 = 'b000011001;
    x_64 = 'b000001001;
    x_65 = 'b000010000;
    x_66 = 'b000001011;
    x_67 = 'b000001011;
    x_68 = 'b000000110;
    x_69 = 'b111111001;
    x_70 = 'b111101110;
    x_71 = 'b000001001;
    x_72 = 'b000010100;
    x_73 = 'b000011010;
    x_74 = 'b000100100;
    x_75 = 'b000010011;
    x_76 = 'b000010010;
    x_77 = 'b000001010;
    x_78 = 'b000010101;
    x_79 = 'b000011110;
    x_80 = 'b000100000;
    x_81 = 'b000100001;
    x_82 = 'b000100011;
    x_83 = 'b000100100;
    x_84 = 'b000010111;
    x_85 = 'b111110111;
    x_86 = 'b111110100;
    x_87 = 'b111101100;
    x_88 = 'b111101111;
    x_89 = 'b111110000;
    x_90 = 'b111101011;
    x_91 = 'b111101100;
    x_92 = 'b111111011;
    x_93 = 'b111111101;
    x_94 = 'b111110001;
    x_95 = 'b111101110;
    x_96 = 'b111111010;
    x_97 = 'b111110100;
    x_98 = 'b111101011;
    x_99 = 'b111101101;
    x_100 = 'b111100110;
    x_101 = 'b111100111;
    x_102 = 'b111111111;
    x_103 = 'b111110111;
    x_104 = 'b000001000;
    x_105 = 'b111001111;
    x_106 = 'b000001000;
    x_107 = 'b000011110;
    x_108 = 'b111111101;
    x_109 = 'b000101001;
    x_110 = 'b000010010;
    x_111 = 'b000011001;
    x_112 = 'b000010110;
    x_113 = 'b000100110;
    x_114 = 'b000101000;
    x_115 = 'b000101101;
    x_116 = 'b000101001;
    x_117 = 'b000100111;
    x_118 = 'b000100110;
    x_119 = 'b000011101;
    x_120 = 'b000011110;
    x_121 = 'b000110000;
    x_122 = 'b000101110;
    x_123 = 'b000110000;
    x_124 = 'b000101001;
    x_125 = 'b000110011;
    x_126 = 'b000011111;
    x_127 = 'b000011001;
    x_128 = 'b000001001;
    x_129 = 'b000010000;
    x_130 = 'b000001011;
    x_131 = 'b000001011;
    x_132 = 'b000000110;
    x_133 = 'b111111001;
    x_134 = 'b111101110;
    x_135 = 'b000001001;
    x_136 = 'b000010100;
    x_137 = 'b000011010;
    x_138 = 'b000100100;
    x_139 = 'b000010011;
    x_140 = 'b000010010;
    x_141 = 'b000001010;
    x_142 = 'b000010101;
    x_143 = 'b000011110;
    x_144 = 'b000100000;
    x_145 = 'b000100001;
    x_146 = 'b000100011;
    x_147 = 'b000100100;
    x_148 = 'b000010111;
    x_149 = 'b111110111;
    x_150 = 'b111110100;
    x_151 = 'b111101100;
    x_152 = 'b111101111;
    x_153 = 'b111110000;
    x_154 = 'b111101011;
    x_155 = 'b111101100;
    x_156 = 'b111111011;
    x_157 = 'b111111101;
    x_158 = 'b111110001;
    x_159 = 'b111101110;
    x_160 = 'b111111010;
    x_161 = 'b111110100;
    x_162 = 'b111101011;
    x_163 = 'b111101101;
    x_164 = 'b111100110;
    x_165 = 'b111100111;
    x_166 = 'b111111111;
    x_167 = 'b111110111;
    x_168 = 'b000001000;
    x_169 = 'b111001111;
    x_170 = 'b000001000;
    x_171 = 'b000011110;
    x_172 = 'b111111101;
    x_173 = 'b000101001;
    x_174 = 'b000010010;
    x_175 = 'b000011001;
    x_176 = 'b000010110;
    x_177 = 'b000100110;
    x_178 = 'b000101000;
    x_179 = 'b000101101;
    x_180 = 'b000101001;
    x_181 = 'b000100111;
    x_182 = 'b000100110;
    x_183 = 'b000011101;
    x_184 = 'b000011110;
    x_185 = 'b000110000;
    x_186 = 'b000101110;
    x_187 = 'b000110000;
    x_188 = 'b000101001;
    x_189 = 'b000110011;
    x_190 = 'b000011111;
    x_191 = 'b000011001;
    x_192 = 'b000001001;
    x_193 = 'b000010000;
    x_194 = 'b000001011;
    x_195 = 'b000001011;
    x_196 = 'b000000110;
    x_197 = 'b111111001;
    x_198 = 'b111101110;
    x_199 = 'b000001001;
    x_200 = 'b000010100;
    x_201 = 'b000011010;
    x_202 = 'b000100100;
    x_203 = 'b000010011;
    x_204 = 'b000010010;
    x_205 = 'b000001010;
    x_206 = 'b000010101;
    x_207 = 'b000011110;
    x_208 = 'b000100000;
    x_209 = 'b000100001;
    x_210 = 'b000100011;
    x_211 = 'b000100100;
    x_212 = 'b000010111;
    x_213 = 'b111110111;
    x_214 = 'b111110100;
    x_215 = 'b111101100;
    x_216 = 'b111101111;
    x_217 = 'b111110000;
    x_218 = 'b111101011;
    x_219 = 'b111101100;
    x_220 = 'b111111011;
    x_221 = 'b111111101;
    x_222 = 'b111110001;
    x_223 = 'b111101110;
    x_224 = 'b111111010;
    x_225 = 'b111110100;
    x_226 = 'b111101011;
    x_227 = 'b111101101;
    x_228 = 'b111100110;
    x_229 = 'b111100111;
    x_230 = 'b111111111;
    x_231 = 'b111110111;
    x_232 = 'b000001000;
    x_233 = 'b111001111;
    x_234 = 'b000001000;
    x_235 = 'b000011110;
    x_236 = 'b111111101;
    x_237 = 'b000101001;
    x_238 = 'b000010010;
    x_239 = 'b000011001;
    x_240 = 'b000010110;
    x_241 = 'b000100110;
    x_242 = 'b000101000;
    x_243 = 'b000101101;
    x_244 = 'b000101001;
    x_245 = 'b000100111;
    x_246 = 'b000100110;
    x_247 = 'b000011101;
    x_248 = 'b000011110;
    x_249 = 'b000110000;
    x_250 = 'b000101110;
    x_251 = 'b000110000;
    x_252 = 'b000101001;
    x_253 = 'b000110011;
    x_254 = 'b000011111;
    x_255 = 'b000011001;

    h_0 = 'b000001001;
    h_1 = 'b000010000;
    h_2 = 'b000001011;
    h_3 = 'b000001011;
    h_4 = 'b000000110;
    h_5 = 'b111111001;
    h_6 = 'b111101110;
    h_7 = 'b000001001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111111001;
    x_1 = 'b111111001;
    x_2 = 'b111101111;
    x_3 = 'b111110101;
    x_4 = 'b111111000;
    x_5 = 'b111110100;
    x_6 = 'b111111001;
    x_7 = 'b111111111;
    x_8 = 'b111110010;
    x_9 = 'b111101011;
    x_10 = 'b111101110;
    x_11 = 'b111101101;
    x_12 = 'b111111000;
    x_13 = 'b000000101;
    x_14 = 'b111110010;
    x_15 = 'b111110011;
    x_16 = 'b111101110;
    x_17 = 'b111101100;
    x_18 = 'b111110101;
    x_19 = 'b111110001;
    x_20 = 'b000000110;
    x_21 = 'b000001100;
    x_22 = 'b000001100;
    x_23 = 'b000000111;
    x_24 = 'b000000111;
    x_25 = 'b000000111;
    x_26 = 'b000000011;
    x_27 = 'b111111011;
    x_28 = 'b111110111;
    x_29 = 'b000000010;
    x_30 = 'b000001000;
    x_31 = 'b111111101;
    x_32 = 'b000000010;
    x_33 = 'b111111010;
    x_34 = 'b111111010;
    x_35 = 'b111111100;
    x_36 = 'b111111000;
    x_37 = 'b111111001;
    x_38 = 'b000000000;
    x_39 = 'b000010010;
    x_40 = 'b111111110;
    x_41 = 'b000110001;
    x_42 = 'b111111010;
    x_43 = 'b000010000;
    x_44 = 'b111110000;
    x_45 = 'b000010101;
    x_46 = 'b111101000;
    x_47 = 'b111110011;
    x_48 = 'b111110011;
    x_49 = 'b111110101;
    x_50 = 'b111110011;
    x_51 = 'b111110111;
    x_52 = 'b111110111;
    x_53 = 'b111111110;
    x_54 = 'b000000110;
    x_55 = 'b111101010;
    x_56 = 'b111110101;
    x_57 = 'b111111000;
    x_58 = 'b111111010;
    x_59 = 'b111111001;
    x_60 = 'b111111001;
    x_61 = 'b111110100;
    x_62 = 'b111110101;
    x_63 = 'b000000010;
    x_64 = 'b111111001;
    x_65 = 'b111111001;
    x_66 = 'b111101111;
    x_67 = 'b111110101;
    x_68 = 'b111111000;
    x_69 = 'b111110100;
    x_70 = 'b111111001;
    x_71 = 'b111111111;
    x_72 = 'b111110010;
    x_73 = 'b111101011;
    x_74 = 'b111101110;
    x_75 = 'b111101101;
    x_76 = 'b111111000;
    x_77 = 'b000000101;
    x_78 = 'b111110010;
    x_79 = 'b111110011;
    x_80 = 'b111101110;
    x_81 = 'b111101100;
    x_82 = 'b111110101;
    x_83 = 'b111110001;
    x_84 = 'b000000110;
    x_85 = 'b000001100;
    x_86 = 'b000001100;
    x_87 = 'b000000111;
    x_88 = 'b000000111;
    x_89 = 'b000000111;
    x_90 = 'b000000011;
    x_91 = 'b111111011;
    x_92 = 'b111110111;
    x_93 = 'b000000010;
    x_94 = 'b000001000;
    x_95 = 'b111111101;
    x_96 = 'b000000010;
    x_97 = 'b111111010;
    x_98 = 'b111111010;
    x_99 = 'b111111100;
    x_100 = 'b111111000;
    x_101 = 'b111111001;
    x_102 = 'b000000000;
    x_103 = 'b000010010;
    x_104 = 'b111111110;
    x_105 = 'b000110001;
    x_106 = 'b111111010;
    x_107 = 'b000010000;
    x_108 = 'b111110000;
    x_109 = 'b000010101;
    x_110 = 'b111101000;
    x_111 = 'b111110011;
    x_112 = 'b111110011;
    x_113 = 'b111110101;
    x_114 = 'b111110011;
    x_115 = 'b111110111;
    x_116 = 'b111110111;
    x_117 = 'b111111110;
    x_118 = 'b000000110;
    x_119 = 'b111101010;
    x_120 = 'b111110101;
    x_121 = 'b111111000;
    x_122 = 'b111111010;
    x_123 = 'b111111001;
    x_124 = 'b111111001;
    x_125 = 'b111110100;
    x_126 = 'b111110101;
    x_127 = 'b000000010;
    x_128 = 'b111111001;
    x_129 = 'b111111001;
    x_130 = 'b111101111;
    x_131 = 'b111110101;
    x_132 = 'b111111000;
    x_133 = 'b111110100;
    x_134 = 'b111111001;
    x_135 = 'b111111111;
    x_136 = 'b111110010;
    x_137 = 'b111101011;
    x_138 = 'b111101110;
    x_139 = 'b111101101;
    x_140 = 'b111111000;
    x_141 = 'b000000101;
    x_142 = 'b111110010;
    x_143 = 'b111110011;
    x_144 = 'b111101110;
    x_145 = 'b111101100;
    x_146 = 'b111110101;
    x_147 = 'b111110001;
    x_148 = 'b000000110;
    x_149 = 'b000001100;
    x_150 = 'b000001100;
    x_151 = 'b000000111;
    x_152 = 'b000000111;
    x_153 = 'b000000111;
    x_154 = 'b000000011;
    x_155 = 'b111111011;
    x_156 = 'b111110111;
    x_157 = 'b000000010;
    x_158 = 'b000001000;
    x_159 = 'b111111101;
    x_160 = 'b000000010;
    x_161 = 'b111111010;
    x_162 = 'b111111010;
    x_163 = 'b111111100;
    x_164 = 'b111111000;
    x_165 = 'b111111001;
    x_166 = 'b000000000;
    x_167 = 'b000010010;
    x_168 = 'b111111110;
    x_169 = 'b000110001;
    x_170 = 'b111111010;
    x_171 = 'b000010000;
    x_172 = 'b111110000;
    x_173 = 'b000010101;
    x_174 = 'b111101000;
    x_175 = 'b111110011;
    x_176 = 'b111110011;
    x_177 = 'b111110101;
    x_178 = 'b111110011;
    x_179 = 'b111110111;
    x_180 = 'b111110111;
    x_181 = 'b111111110;
    x_182 = 'b000000110;
    x_183 = 'b111101010;
    x_184 = 'b111110101;
    x_185 = 'b111111000;
    x_186 = 'b111111010;
    x_187 = 'b111111001;
    x_188 = 'b111111001;
    x_189 = 'b111110100;
    x_190 = 'b111110101;
    x_191 = 'b000000010;
    x_192 = 'b111111001;
    x_193 = 'b111111001;
    x_194 = 'b111101111;
    x_195 = 'b111110101;
    x_196 = 'b111111000;
    x_197 = 'b111110100;
    x_198 = 'b111111001;
    x_199 = 'b111111111;
    x_200 = 'b111110010;
    x_201 = 'b111101011;
    x_202 = 'b111101110;
    x_203 = 'b111101101;
    x_204 = 'b111111000;
    x_205 = 'b000000101;
    x_206 = 'b111110010;
    x_207 = 'b111110011;
    x_208 = 'b111101110;
    x_209 = 'b111101100;
    x_210 = 'b111110101;
    x_211 = 'b111110001;
    x_212 = 'b000000110;
    x_213 = 'b000001100;
    x_214 = 'b000001100;
    x_215 = 'b000000111;
    x_216 = 'b000000111;
    x_217 = 'b000000111;
    x_218 = 'b000000011;
    x_219 = 'b111111011;
    x_220 = 'b111110111;
    x_221 = 'b000000010;
    x_222 = 'b000001000;
    x_223 = 'b111111101;
    x_224 = 'b000000010;
    x_225 = 'b111111010;
    x_226 = 'b111111010;
    x_227 = 'b111111100;
    x_228 = 'b111111000;
    x_229 = 'b111111001;
    x_230 = 'b000000000;
    x_231 = 'b000010010;
    x_232 = 'b111111110;
    x_233 = 'b000110001;
    x_234 = 'b111111010;
    x_235 = 'b000010000;
    x_236 = 'b111110000;
    x_237 = 'b000010101;
    x_238 = 'b111101000;
    x_239 = 'b111110011;
    x_240 = 'b111110011;
    x_241 = 'b111110101;
    x_242 = 'b111110011;
    x_243 = 'b111110111;
    x_244 = 'b111110111;
    x_245 = 'b111111110;
    x_246 = 'b000000110;
    x_247 = 'b111101010;
    x_248 = 'b111110101;
    x_249 = 'b111111000;
    x_250 = 'b111111010;
    x_251 = 'b111111001;
    x_252 = 'b111111001;
    x_253 = 'b111110100;
    x_254 = 'b111110101;
    x_255 = 'b000000010;

    h_0 = 'b111111001;
    h_1 = 'b111111001;
    h_2 = 'b111101111;
    h_3 = 'b111110101;
    h_4 = 'b111111000;
    h_5 = 'b111110100;
    h_6 = 'b111111001;
    h_7 = 'b111111111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b000000001;
    x_1 = 'b000000000;
    x_2 = 'b111110101;
    x_3 = 'b111111101;
    x_4 = 'b111111100;
    x_5 = 'b111110111;
    x_6 = 'b111111010;
    x_7 = 'b000000011;
    x_8 = 'b111110100;
    x_9 = 'b111101110;
    x_10 = 'b111110011;
    x_11 = 'b111110011;
    x_12 = 'b111111010;
    x_13 = 'b000001011;
    x_14 = 'b111110011;
    x_15 = 'b111110000;
    x_16 = 'b111101110;
    x_17 = 'b111101110;
    x_18 = 'b111110101;
    x_19 = 'b111101111;
    x_20 = 'b000000011;
    x_21 = 'b000001101;
    x_22 = 'b000001011;
    x_23 = 'b000000110;
    x_24 = 'b000001000;
    x_25 = 'b000000111;
    x_26 = 'b000000010;
    x_27 = 'b111111100;
    x_28 = 'b111110101;
    x_29 = 'b000000010;
    x_30 = 'b000001000;
    x_31 = 'b111111110;
    x_32 = 'b000000010;
    x_33 = 'b111111001;
    x_34 = 'b111111001;
    x_35 = 'b111111001;
    x_36 = 'b111110111;
    x_37 = 'b111110100;
    x_38 = 'b111111111;
    x_39 = 'b000001001;
    x_40 = 'b111110111;
    x_41 = 'b000000101;
    x_42 = 'b111110011;
    x_43 = 'b000001001;
    x_44 = 'b111101000;
    x_45 = 'b000001010;
    x_46 = 'b111100001;
    x_47 = 'b111101010;
    x_48 = 'b111101011;
    x_49 = 'b111101110;
    x_50 = 'b111101101;
    x_51 = 'b111110000;
    x_52 = 'b111110000;
    x_53 = 'b111110100;
    x_54 = 'b111110111;
    x_55 = 'b111011111;
    x_56 = 'b111101010;
    x_57 = 'b111101111;
    x_58 = 'b111110011;
    x_59 = 'b111110100;
    x_60 = 'b111110010;
    x_61 = 'b111110000;
    x_62 = 'b111110100;
    x_63 = 'b111111101;
    x_64 = 'b000000001;
    x_65 = 'b000000000;
    x_66 = 'b111110101;
    x_67 = 'b111111101;
    x_68 = 'b111111100;
    x_69 = 'b111110111;
    x_70 = 'b111111010;
    x_71 = 'b000000011;
    x_72 = 'b111110100;
    x_73 = 'b111101110;
    x_74 = 'b111110011;
    x_75 = 'b111110011;
    x_76 = 'b111111010;
    x_77 = 'b000001011;
    x_78 = 'b111110011;
    x_79 = 'b111110000;
    x_80 = 'b111101110;
    x_81 = 'b111101110;
    x_82 = 'b111110101;
    x_83 = 'b111101111;
    x_84 = 'b000000011;
    x_85 = 'b000001101;
    x_86 = 'b000001011;
    x_87 = 'b000000110;
    x_88 = 'b000001000;
    x_89 = 'b000000111;
    x_90 = 'b000000010;
    x_91 = 'b111111100;
    x_92 = 'b111110101;
    x_93 = 'b000000010;
    x_94 = 'b000001000;
    x_95 = 'b111111110;
    x_96 = 'b000000010;
    x_97 = 'b111111001;
    x_98 = 'b111111001;
    x_99 = 'b111111001;
    x_100 = 'b111110111;
    x_101 = 'b111110100;
    x_102 = 'b111111111;
    x_103 = 'b000001001;
    x_104 = 'b111110111;
    x_105 = 'b000000101;
    x_106 = 'b111110011;
    x_107 = 'b000001001;
    x_108 = 'b111101000;
    x_109 = 'b000001010;
    x_110 = 'b111100001;
    x_111 = 'b111101010;
    x_112 = 'b111101011;
    x_113 = 'b111101110;
    x_114 = 'b111101101;
    x_115 = 'b111110000;
    x_116 = 'b111110000;
    x_117 = 'b111110100;
    x_118 = 'b111110111;
    x_119 = 'b111011111;
    x_120 = 'b111101010;
    x_121 = 'b111101111;
    x_122 = 'b111110011;
    x_123 = 'b111110100;
    x_124 = 'b111110010;
    x_125 = 'b111110000;
    x_126 = 'b111110100;
    x_127 = 'b111111101;
    x_128 = 'b000000001;
    x_129 = 'b000000000;
    x_130 = 'b111110101;
    x_131 = 'b111111101;
    x_132 = 'b111111100;
    x_133 = 'b111110111;
    x_134 = 'b111111010;
    x_135 = 'b000000011;
    x_136 = 'b111110100;
    x_137 = 'b111101110;
    x_138 = 'b111110011;
    x_139 = 'b111110011;
    x_140 = 'b111111010;
    x_141 = 'b000001011;
    x_142 = 'b111110011;
    x_143 = 'b111110000;
    x_144 = 'b111101110;
    x_145 = 'b111101110;
    x_146 = 'b111110101;
    x_147 = 'b111101111;
    x_148 = 'b000000011;
    x_149 = 'b000001101;
    x_150 = 'b000001011;
    x_151 = 'b000000110;
    x_152 = 'b000001000;
    x_153 = 'b000000111;
    x_154 = 'b000000010;
    x_155 = 'b111111100;
    x_156 = 'b111110101;
    x_157 = 'b000000010;
    x_158 = 'b000001000;
    x_159 = 'b111111110;
    x_160 = 'b000000010;
    x_161 = 'b111111001;
    x_162 = 'b111111001;
    x_163 = 'b111111001;
    x_164 = 'b111110111;
    x_165 = 'b111110100;
    x_166 = 'b111111111;
    x_167 = 'b000001001;
    x_168 = 'b111110111;
    x_169 = 'b000000101;
    x_170 = 'b111110011;
    x_171 = 'b000001001;
    x_172 = 'b111101000;
    x_173 = 'b000001010;
    x_174 = 'b111100001;
    x_175 = 'b111101010;
    x_176 = 'b111101011;
    x_177 = 'b111101110;
    x_178 = 'b111101101;
    x_179 = 'b111110000;
    x_180 = 'b111110000;
    x_181 = 'b111110100;
    x_182 = 'b111110111;
    x_183 = 'b111011111;
    x_184 = 'b111101010;
    x_185 = 'b111101111;
    x_186 = 'b111110011;
    x_187 = 'b111110100;
    x_188 = 'b111110010;
    x_189 = 'b111110000;
    x_190 = 'b111110100;
    x_191 = 'b111111101;
    x_192 = 'b000000001;
    x_193 = 'b000000000;
    x_194 = 'b111110101;
    x_195 = 'b111111101;
    x_196 = 'b111111100;
    x_197 = 'b111110111;
    x_198 = 'b111111010;
    x_199 = 'b000000011;
    x_200 = 'b111110100;
    x_201 = 'b111101110;
    x_202 = 'b111110011;
    x_203 = 'b111110011;
    x_204 = 'b111111010;
    x_205 = 'b000001011;
    x_206 = 'b111110011;
    x_207 = 'b111110000;
    x_208 = 'b111101110;
    x_209 = 'b111101110;
    x_210 = 'b111110101;
    x_211 = 'b111101111;
    x_212 = 'b000000011;
    x_213 = 'b000001101;
    x_214 = 'b000001011;
    x_215 = 'b000000110;
    x_216 = 'b000001000;
    x_217 = 'b000000111;
    x_218 = 'b000000010;
    x_219 = 'b111111100;
    x_220 = 'b111110101;
    x_221 = 'b000000010;
    x_222 = 'b000001000;
    x_223 = 'b111111110;
    x_224 = 'b000000010;
    x_225 = 'b111111001;
    x_226 = 'b111111001;
    x_227 = 'b111111001;
    x_228 = 'b111110111;
    x_229 = 'b111110100;
    x_230 = 'b111111111;
    x_231 = 'b000001001;
    x_232 = 'b111110111;
    x_233 = 'b000000101;
    x_234 = 'b111110011;
    x_235 = 'b000001001;
    x_236 = 'b111101000;
    x_237 = 'b000001010;
    x_238 = 'b111100001;
    x_239 = 'b111101010;
    x_240 = 'b111101011;
    x_241 = 'b111101110;
    x_242 = 'b111101101;
    x_243 = 'b111110000;
    x_244 = 'b111110000;
    x_245 = 'b111110100;
    x_246 = 'b111110111;
    x_247 = 'b111011111;
    x_248 = 'b111101010;
    x_249 = 'b111101111;
    x_250 = 'b111110011;
    x_251 = 'b111110100;
    x_252 = 'b111110010;
    x_253 = 'b111110000;
    x_254 = 'b111110100;
    x_255 = 'b111111101;

    h_0 = 'b000000001;
    h_1 = 'b000000000;
    h_2 = 'b111110101;
    h_3 = 'b111111101;
    h_4 = 'b111111100;
    h_5 = 'b111110111;
    h_6 = 'b111111010;
    h_7 = 'b000000011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111110111;
    x_1 = 'b111110101;
    x_2 = 'b111101100;
    x_3 = 'b111110100;
    x_4 = 'b111110011;
    x_5 = 'b111101110;
    x_6 = 'b111101110;
    x_7 = 'b111110101;
    x_8 = 'b111100101;
    x_9 = 'b111100000;
    x_10 = 'b111100110;
    x_11 = 'b111100100;
    x_12 = 'b111101000;
    x_13 = 'b111110010;
    x_14 = 'b111100110;
    x_15 = 'b111011111;
    x_16 = 'b111011100;
    x_17 = 'b111011111;
    x_18 = 'b111100011;
    x_19 = 'b111011010;
    x_20 = 'b111100110;
    x_21 = 'b000001001;
    x_22 = 'b000000111;
    x_23 = 'b000000011;
    x_24 = 'b000000001;
    x_25 = 'b000000001;
    x_26 = 'b111111010;
    x_27 = 'b111110101;
    x_28 = 'b111110000;
    x_29 = 'b111111011;
    x_30 = 'b000000001;
    x_31 = 'b111110101;
    x_32 = 'b111110111;
    x_33 = 'b111101111;
    x_34 = 'b111110000;
    x_35 = 'b111110001;
    x_36 = 'b111101100;
    x_37 = 'b111101100;
    x_38 = 'b111111000;
    x_39 = 'b111110010;
    x_40 = 'b111110001;
    x_41 = 'b111100011;
    x_42 = 'b111101110;
    x_43 = 'b111110110;
    x_44 = 'b111100010;
    x_45 = 'b111100001;
    x_46 = 'b111011001;
    x_47 = 'b111011100;
    x_48 = 'b111011010;
    x_49 = 'b111011001;
    x_50 = 'b111011001;
    x_51 = 'b111011000;
    x_52 = 'b111010101;
    x_53 = 'b111010011;
    x_54 = 'b111001110;
    x_55 = 'b111010011;
    x_56 = 'b111011010;
    x_57 = 'b111011100;
    x_58 = 'b111011100;
    x_59 = 'b111011001;
    x_60 = 'b111100111;
    x_61 = 'b111100011;
    x_62 = 'b111101001;
    x_63 = 'b111110000;
    x_64 = 'b111110111;
    x_65 = 'b111110101;
    x_66 = 'b111101100;
    x_67 = 'b111110100;
    x_68 = 'b111110011;
    x_69 = 'b111101110;
    x_70 = 'b111101110;
    x_71 = 'b111110101;
    x_72 = 'b111100101;
    x_73 = 'b111100000;
    x_74 = 'b111100110;
    x_75 = 'b111100100;
    x_76 = 'b111101000;
    x_77 = 'b111110010;
    x_78 = 'b111100110;
    x_79 = 'b111011111;
    x_80 = 'b111011100;
    x_81 = 'b111011111;
    x_82 = 'b111100011;
    x_83 = 'b111011010;
    x_84 = 'b111100110;
    x_85 = 'b000001001;
    x_86 = 'b000000111;
    x_87 = 'b000000011;
    x_88 = 'b000000001;
    x_89 = 'b000000001;
    x_90 = 'b111111010;
    x_91 = 'b111110101;
    x_92 = 'b111110000;
    x_93 = 'b111111011;
    x_94 = 'b000000001;
    x_95 = 'b111110101;
    x_96 = 'b111110111;
    x_97 = 'b111101111;
    x_98 = 'b111110000;
    x_99 = 'b111110001;
    x_100 = 'b111101100;
    x_101 = 'b111101100;
    x_102 = 'b111111000;
    x_103 = 'b111110010;
    x_104 = 'b111110001;
    x_105 = 'b111100011;
    x_106 = 'b111101110;
    x_107 = 'b111110110;
    x_108 = 'b111100010;
    x_109 = 'b111100001;
    x_110 = 'b111011001;
    x_111 = 'b111011100;
    x_112 = 'b111011010;
    x_113 = 'b111011001;
    x_114 = 'b111011001;
    x_115 = 'b111011000;
    x_116 = 'b111010101;
    x_117 = 'b111010011;
    x_118 = 'b111001110;
    x_119 = 'b111010011;
    x_120 = 'b111011010;
    x_121 = 'b111011100;
    x_122 = 'b111011100;
    x_123 = 'b111011001;
    x_124 = 'b111100111;
    x_125 = 'b111100011;
    x_126 = 'b111101001;
    x_127 = 'b111110000;
    x_128 = 'b111110111;
    x_129 = 'b111110101;
    x_130 = 'b111101100;
    x_131 = 'b111110100;
    x_132 = 'b111110011;
    x_133 = 'b111101110;
    x_134 = 'b111101110;
    x_135 = 'b111110101;
    x_136 = 'b111100101;
    x_137 = 'b111100000;
    x_138 = 'b111100110;
    x_139 = 'b111100100;
    x_140 = 'b111101000;
    x_141 = 'b111110010;
    x_142 = 'b111100110;
    x_143 = 'b111011111;
    x_144 = 'b111011100;
    x_145 = 'b111011111;
    x_146 = 'b111100011;
    x_147 = 'b111011010;
    x_148 = 'b111100110;
    x_149 = 'b000001001;
    x_150 = 'b000000111;
    x_151 = 'b000000011;
    x_152 = 'b000000001;
    x_153 = 'b000000001;
    x_154 = 'b111111010;
    x_155 = 'b111110101;
    x_156 = 'b111110000;
    x_157 = 'b111111011;
    x_158 = 'b000000001;
    x_159 = 'b111110101;
    x_160 = 'b111110111;
    x_161 = 'b111101111;
    x_162 = 'b111110000;
    x_163 = 'b111110001;
    x_164 = 'b111101100;
    x_165 = 'b111101100;
    x_166 = 'b111111000;
    x_167 = 'b111110010;
    x_168 = 'b111110001;
    x_169 = 'b111100011;
    x_170 = 'b111101110;
    x_171 = 'b111110110;
    x_172 = 'b111100010;
    x_173 = 'b111100001;
    x_174 = 'b111011001;
    x_175 = 'b111011100;
    x_176 = 'b111011010;
    x_177 = 'b111011001;
    x_178 = 'b111011001;
    x_179 = 'b111011000;
    x_180 = 'b111010101;
    x_181 = 'b111010011;
    x_182 = 'b111001110;
    x_183 = 'b111010011;
    x_184 = 'b111011010;
    x_185 = 'b111011100;
    x_186 = 'b111011100;
    x_187 = 'b111011001;
    x_188 = 'b111100111;
    x_189 = 'b111100011;
    x_190 = 'b111101001;
    x_191 = 'b111110000;
    x_192 = 'b111110111;
    x_193 = 'b111110101;
    x_194 = 'b111101100;
    x_195 = 'b111110100;
    x_196 = 'b111110011;
    x_197 = 'b111101110;
    x_198 = 'b111101110;
    x_199 = 'b111110101;
    x_200 = 'b111100101;
    x_201 = 'b111100000;
    x_202 = 'b111100110;
    x_203 = 'b111100100;
    x_204 = 'b111101000;
    x_205 = 'b111110010;
    x_206 = 'b111100110;
    x_207 = 'b111011111;
    x_208 = 'b111011100;
    x_209 = 'b111011111;
    x_210 = 'b111100011;
    x_211 = 'b111011010;
    x_212 = 'b111100110;
    x_213 = 'b000001001;
    x_214 = 'b000000111;
    x_215 = 'b000000011;
    x_216 = 'b000000001;
    x_217 = 'b000000001;
    x_218 = 'b111111010;
    x_219 = 'b111110101;
    x_220 = 'b111110000;
    x_221 = 'b111111011;
    x_222 = 'b000000001;
    x_223 = 'b111110101;
    x_224 = 'b111110111;
    x_225 = 'b111101111;
    x_226 = 'b111110000;
    x_227 = 'b111110001;
    x_228 = 'b111101100;
    x_229 = 'b111101100;
    x_230 = 'b111111000;
    x_231 = 'b111110010;
    x_232 = 'b111110001;
    x_233 = 'b111100011;
    x_234 = 'b111101110;
    x_235 = 'b111110110;
    x_236 = 'b111100010;
    x_237 = 'b111100001;
    x_238 = 'b111011001;
    x_239 = 'b111011100;
    x_240 = 'b111011010;
    x_241 = 'b111011001;
    x_242 = 'b111011001;
    x_243 = 'b111011000;
    x_244 = 'b111010101;
    x_245 = 'b111010011;
    x_246 = 'b111001110;
    x_247 = 'b111010011;
    x_248 = 'b111011010;
    x_249 = 'b111011100;
    x_250 = 'b111011100;
    x_251 = 'b111011001;
    x_252 = 'b111100111;
    x_253 = 'b111100011;
    x_254 = 'b111101001;
    x_255 = 'b111110000;

    h_0 = 'b111110111;
    h_1 = 'b111110101;
    h_2 = 'b111101100;
    h_3 = 'b111110100;
    h_4 = 'b111110011;
    h_5 = 'b111101110;
    h_6 = 'b111101110;
    h_7 = 'b111110101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b111110111;
    x_1 = 'b111110010;
    x_2 = 'b111100101;
    x_3 = 'b111101111;
    x_4 = 'b111101111;
    x_5 = 'b111101001;
    x_6 = 'b111101100;
    x_7 = 'b111111001;
    x_8 = 'b111011111;
    x_9 = 'b111011000;
    x_10 = 'b111011011;
    x_11 = 'b111011000;
    x_12 = 'b111011001;
    x_13 = 'b111100010;
    x_14 = 'b111100111;
    x_15 = 'b111011011;
    x_16 = 'b111010010;
    x_17 = 'b111010011;
    x_18 = 'b111011000;
    x_19 = 'b111001001;
    x_20 = 'b111010010;
    x_21 = 'b000010001;
    x_22 = 'b000010010;
    x_23 = 'b000001101;
    x_24 = 'b000001011;
    x_25 = 'b000001010;
    x_26 = 'b000000110;
    x_27 = 'b000000001;
    x_28 = 'b111111001;
    x_29 = 'b000001001;
    x_30 = 'b000001001;
    x_31 = 'b111111110;
    x_32 = 'b111111110;
    x_33 = 'b111111011;
    x_34 = 'b111111101;
    x_35 = 'b111111101;
    x_36 = 'b111111011;
    x_37 = 'b111111010;
    x_38 = 'b000000110;
    x_39 = 'b111111101;
    x_40 = 'b000000011;
    x_41 = 'b111111000;
    x_42 = 'b000000100;
    x_43 = 'b111011011;
    x_44 = 'b111101001;
    x_45 = 'b111000100;
    x_46 = 'b111011101;
    x_47 = 'b111011100;
    x_48 = 'b111010111;
    x_49 = 'b111010010;
    x_50 = 'b111010000;
    x_51 = 'b111001111;
    x_52 = 'b111001110;
    x_53 = 'b111001000;
    x_54 = 'b111000010;
    x_55 = 'b111001111;
    x_56 = 'b111010010;
    x_57 = 'b111010100;
    x_58 = 'b111010011;
    x_59 = 'b111010000;
    x_60 = 'b111011110;
    x_61 = 'b111011000;
    x_62 = 'b111011110;
    x_63 = 'b111101011;
    x_64 = 'b111110111;
    x_65 = 'b111110010;
    x_66 = 'b111100101;
    x_67 = 'b111101111;
    x_68 = 'b111101111;
    x_69 = 'b111101001;
    x_70 = 'b111101100;
    x_71 = 'b111111001;
    x_72 = 'b111011111;
    x_73 = 'b111011000;
    x_74 = 'b111011011;
    x_75 = 'b111011000;
    x_76 = 'b111011001;
    x_77 = 'b111100010;
    x_78 = 'b111100111;
    x_79 = 'b111011011;
    x_80 = 'b111010010;
    x_81 = 'b111010011;
    x_82 = 'b111011000;
    x_83 = 'b111001001;
    x_84 = 'b111010010;
    x_85 = 'b000010001;
    x_86 = 'b000010010;
    x_87 = 'b000001101;
    x_88 = 'b000001011;
    x_89 = 'b000001010;
    x_90 = 'b000000110;
    x_91 = 'b000000001;
    x_92 = 'b111111001;
    x_93 = 'b000001001;
    x_94 = 'b000001001;
    x_95 = 'b111111110;
    x_96 = 'b111111110;
    x_97 = 'b111111011;
    x_98 = 'b111111101;
    x_99 = 'b111111101;
    x_100 = 'b111111011;
    x_101 = 'b111111010;
    x_102 = 'b000000110;
    x_103 = 'b111111101;
    x_104 = 'b000000011;
    x_105 = 'b111111000;
    x_106 = 'b000000100;
    x_107 = 'b111011011;
    x_108 = 'b111101001;
    x_109 = 'b111000100;
    x_110 = 'b111011101;
    x_111 = 'b111011100;
    x_112 = 'b111010111;
    x_113 = 'b111010010;
    x_114 = 'b111010000;
    x_115 = 'b111001111;
    x_116 = 'b111001110;
    x_117 = 'b111001000;
    x_118 = 'b111000010;
    x_119 = 'b111001111;
    x_120 = 'b111010010;
    x_121 = 'b111010100;
    x_122 = 'b111010011;
    x_123 = 'b111010000;
    x_124 = 'b111011110;
    x_125 = 'b111011000;
    x_126 = 'b111011110;
    x_127 = 'b111101011;
    x_128 = 'b111110111;
    x_129 = 'b111110010;
    x_130 = 'b111100101;
    x_131 = 'b111101111;
    x_132 = 'b111101111;
    x_133 = 'b111101001;
    x_134 = 'b111101100;
    x_135 = 'b111111001;
    x_136 = 'b111011111;
    x_137 = 'b111011000;
    x_138 = 'b111011011;
    x_139 = 'b111011000;
    x_140 = 'b111011001;
    x_141 = 'b111100010;
    x_142 = 'b111100111;
    x_143 = 'b111011011;
    x_144 = 'b111010010;
    x_145 = 'b111010011;
    x_146 = 'b111011000;
    x_147 = 'b111001001;
    x_148 = 'b111010010;
    x_149 = 'b000010001;
    x_150 = 'b000010010;
    x_151 = 'b000001101;
    x_152 = 'b000001011;
    x_153 = 'b000001010;
    x_154 = 'b000000110;
    x_155 = 'b000000001;
    x_156 = 'b111111001;
    x_157 = 'b000001001;
    x_158 = 'b000001001;
    x_159 = 'b111111110;
    x_160 = 'b111111110;
    x_161 = 'b111111011;
    x_162 = 'b111111101;
    x_163 = 'b111111101;
    x_164 = 'b111111011;
    x_165 = 'b111111010;
    x_166 = 'b000000110;
    x_167 = 'b111111101;
    x_168 = 'b000000011;
    x_169 = 'b111111000;
    x_170 = 'b000000100;
    x_171 = 'b111011011;
    x_172 = 'b111101001;
    x_173 = 'b111000100;
    x_174 = 'b111011101;
    x_175 = 'b111011100;
    x_176 = 'b111010111;
    x_177 = 'b111010010;
    x_178 = 'b111010000;
    x_179 = 'b111001111;
    x_180 = 'b111001110;
    x_181 = 'b111001000;
    x_182 = 'b111000010;
    x_183 = 'b111001111;
    x_184 = 'b111010010;
    x_185 = 'b111010100;
    x_186 = 'b111010011;
    x_187 = 'b111010000;
    x_188 = 'b111011110;
    x_189 = 'b111011000;
    x_190 = 'b111011110;
    x_191 = 'b111101011;
    x_192 = 'b111110111;
    x_193 = 'b111110010;
    x_194 = 'b111100101;
    x_195 = 'b111101111;
    x_196 = 'b111101111;
    x_197 = 'b111101001;
    x_198 = 'b111101100;
    x_199 = 'b111111001;
    x_200 = 'b111011111;
    x_201 = 'b111011000;
    x_202 = 'b111011011;
    x_203 = 'b111011000;
    x_204 = 'b111011001;
    x_205 = 'b111100010;
    x_206 = 'b111100111;
    x_207 = 'b111011011;
    x_208 = 'b111010010;
    x_209 = 'b111010011;
    x_210 = 'b111011000;
    x_211 = 'b111001001;
    x_212 = 'b111010010;
    x_213 = 'b000010001;
    x_214 = 'b000010010;
    x_215 = 'b000001101;
    x_216 = 'b000001011;
    x_217 = 'b000001010;
    x_218 = 'b000000110;
    x_219 = 'b000000001;
    x_220 = 'b111111001;
    x_221 = 'b000001001;
    x_222 = 'b000001001;
    x_223 = 'b111111110;
    x_224 = 'b111111110;
    x_225 = 'b111111011;
    x_226 = 'b111111101;
    x_227 = 'b111111101;
    x_228 = 'b111111011;
    x_229 = 'b111111010;
    x_230 = 'b000000110;
    x_231 = 'b111111101;
    x_232 = 'b000000011;
    x_233 = 'b111111000;
    x_234 = 'b000000100;
    x_235 = 'b111011011;
    x_236 = 'b111101001;
    x_237 = 'b111000100;
    x_238 = 'b111011101;
    x_239 = 'b111011100;
    x_240 = 'b111010111;
    x_241 = 'b111010010;
    x_242 = 'b111010000;
    x_243 = 'b111001111;
    x_244 = 'b111001110;
    x_245 = 'b111001000;
    x_246 = 'b111000010;
    x_247 = 'b111001111;
    x_248 = 'b111010010;
    x_249 = 'b111010100;
    x_250 = 'b111010011;
    x_251 = 'b111010000;
    x_252 = 'b111011110;
    x_253 = 'b111011000;
    x_254 = 'b111011110;
    x_255 = 'b111101011;

    h_0 = 'b111110111;
    h_1 = 'b111110010;
    h_2 = 'b111100101;
    h_3 = 'b111101111;
    h_4 = 'b111101111;
    h_5 = 'b111101001;
    h_6 = 'b111101100;
    h_7 = 'b111111001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b %09b %09b %09b %09b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    $fclose(fd);    
$finish;
    end
endmodule