`timescale 1ns / 1ps

module gru_tb;

// Parameters
parameter int D          = 64;
parameter int H          = 16;
parameter int DATA_WIDTH = 26;
parameter int FRAC_BITS  = 16;
parameter int NUM_PARALLEL = 16;
parameter real CLK_PERIOD = 10.0;

// Clock and reset
logic clk;
logic rst_n;
logic start;
logic done;

// Cycle counter
int cycle_count = 0;
int test_start_cycle = 0;
int test_cycles = 0;
int total_cycles = 0;
bit test_timeout = 0;

// Input arrays
logic signed [DATA_WIDTH-1:0] x_t [D-1:0];
logic signed [DATA_WIDTH-1:0] h_t_prev [H-1:0];
logic signed [DATA_WIDTH-1:0] h_t [H-1:0];

// Weight matrices
logic signed [DATA_WIDTH-1:0] W_ir [H-1:0][D-1:0];
logic signed [DATA_WIDTH-1:0] W_hr [H-1:0][H-1:0];
logic signed [DATA_WIDTH-1:0] b_ir [H-1:0];
logic signed [DATA_WIDTH-1:0] b_hr [H-1:0];

logic signed [DATA_WIDTH-1:0] W_iz [H-1:0][D-1:0];
logic signed [DATA_WIDTH-1:0] W_hz [H-1:0][H-1:0];
logic signed [DATA_WIDTH-1:0] b_iz [H-1:0];
logic signed [DATA_WIDTH-1:0] b_hz [H-1:0];

logic signed [DATA_WIDTH-1:0] W_in [H-1:0][D-1:0];
logic signed [DATA_WIDTH-1:0] W_hn [H-1:0][H-1:0];
logic signed [DATA_WIDTH-1:0] b_in [H-1:0];
logic signed [DATA_WIDTH-1:0] b_hn [H-1:0];

// DUT instantiation
gru_cell_parallel #(
    .D(D),
    .H(H),
    .DATA_WIDTH(DATA_WIDTH),
    .FRAC_BITS(FRAC_BITS),
    .NUM_PARALLEL(NUM_PARALLEL)
) dut (
    .clk(clk),
    .rst_n(rst_n),
    .start(start),
    .x_t(x_t),
    .h_t_prev(h_t_prev),
    .W_ir(W_ir),
    .W_hr(W_hr),
    .b_ir(b_ir),
    .b_hr(b_hr),
    .W_iz(W_iz),
    .W_hz(W_hz),
    .b_iz(b_iz),
    .b_hz(b_hz),
    .W_in(W_in),
    .W_hn(W_hn),
    .b_in(b_in),
    .b_hn(b_hn),
    .h_t(h_t),
    .done(done)
);

// Clock generation
initial begin
    clk = 0;
    forever #5 clk = ~clk; // 100MHz clock
end

// Cycle counter
always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        cycle_count <= 0;
    end else begin
        cycle_count <= cycle_count + 1;
    end
end

initial begin
    // Open files for writing
    integer fd_output;
    integer fd_cycles;
    
    fd_output = $fopen("../../../../../output_d64_h16_dw26_fb16_np16.txt", "w+");
    if (fd_output == 0) begin
        $display("ERROR: Failed to open output file!");
        $finish;
    end
    
    fd_cycles = $fopen("../../../../../cycles_d64_h16_dw26_fb16_np16.txt", "w+");
    if (fd_cycles == 0) begin
        $display("ERROR: Failed to open cycles file!");
        $fclose(fd_output);
        $finish;
    end
    
    // Write header to cycles file
    $fdisplay(fd_cycles, "==========================================================");
    $fdisplay(fd_cycles, "GRU Cell Parallel Cycle Count Results");
    $fdisplay(fd_cycles, "==========================================================");
    $fdisplay(fd_cycles, "Parameters:");
    $fdisplay(fd_cycles, "  D (Input Dimension):     64");
    $fdisplay(fd_cycles, "  H (Hidden Dimension):    16");
    $fdisplay(fd_cycles, "  DATA_WIDTH:              26");
    $fdisplay(fd_cycles, "  FRAC_BITS:               16");
    $fdisplay(fd_cycles, "  NUM_PARALLEL:            16");
    $fdisplay(fd_cycles, "  Total Test Vectors:      100");
    $fdisplay(fd_cycles, "==========================================================");
    $fdisplay(fd_cycles, "");
    
    // Initialize weights
    // Initialize W_ir weights
    W_ir[0][0] = 26'b00000000000001010010011110;
    W_ir[0][1] = 26'b00000000000010011100011000;
    W_ir[0][2] = 26'b00000000000001110111001110;
    W_ir[0][3] = 26'b00000000000010001100110010;
    W_ir[0][4] = 26'b11111111111110110100110100;
    W_ir[0][5] = 26'b11111111111101010101000001;
    W_ir[0][6] = 26'b00000000000001110011010001;
    W_ir[0][7] = 26'b00000000000000111101101110;
    W_ir[0][8] = 26'b11111111111100100000101110;
    W_ir[0][9] = 26'b00000000000000010110011000;
    W_ir[0][10] = 26'b00000000000011111010111111;
    W_ir[0][11] = 26'b11111111111111111110101100;
    W_ir[0][12] = 26'b00000000000010011111111001;
    W_ir[0][13] = 26'b00000000000000101100000000;
    W_ir[0][14] = 26'b00000000000000100111011101;
    W_ir[0][15] = 26'b00000000000010111001011010;
    W_ir[0][16] = 26'b11111111111111100000000101;
    W_ir[0][17] = 26'b00000000000011011100110111;
    W_ir[0][18] = 26'b11111111111111100011001001;
    W_ir[0][19] = 26'b00000000000010010001001011;
    W_ir[0][20] = 26'b11111111111111100001111100;
    W_ir[0][21] = 26'b00000000000010000111001000;
    W_ir[0][22] = 26'b00000000000001100001111111;
    W_ir[0][23] = 26'b00000000000001100011100000;
    W_ir[0][24] = 26'b11111111111101011110111110;
    W_ir[0][25] = 26'b00000000000001111000001100;
    W_ir[0][26] = 26'b00000000000010001011100110;
    W_ir[0][27] = 26'b00000000000001011011010101;
    W_ir[0][28] = 26'b00000000000011100010100110;
    W_ir[0][29] = 26'b11111111111100101100001011;
    W_ir[0][30] = 26'b11111111111110110101100001;
    W_ir[0][31] = 26'b00000000000001100111000001;
    W_ir[0][32] = 26'b00000000000000110001101110;
    W_ir[0][33] = 26'b00000000000001111010001100;
    W_ir[0][34] = 26'b00000000000001111010011110;
    W_ir[0][35] = 26'b00000000000000011010111101;
    W_ir[0][36] = 26'b00000000000011111110101101;
    W_ir[0][37] = 26'b00000000000001010001000000;
    W_ir[0][38] = 26'b11111111111110111011001110;
    W_ir[0][39] = 26'b00000000000000111101100110;
    W_ir[0][40] = 26'b00000000000010010101101000;
    W_ir[0][41] = 26'b11111111111101000000111011;
    W_ir[0][42] = 26'b00000000000000111100111010;
    W_ir[0][43] = 26'b11111111111110100001001011;
    W_ir[0][44] = 26'b11111111111111111001001101;
    W_ir[0][45] = 26'b11111111111101110010100010;
    W_ir[0][46] = 26'b11111111111100111001111111;
    W_ir[0][47] = 26'b00000000000011011110110000;
    W_ir[0][48] = 26'b11111111111111000101001111;
    W_ir[0][49] = 26'b11111111111110011100100001;
    W_ir[0][50] = 26'b11111111111111100110010101;
    W_ir[0][51] = 26'b00000000000000000001001000;
    W_ir[0][52] = 26'b11111111111100011011000001;
    W_ir[0][53] = 26'b11111111111110101001001010;
    W_ir[0][54] = 26'b00000000000001000011001101;
    W_ir[0][55] = 26'b11111111111110011111000000;
    W_ir[0][56] = 26'b00000000000010011001010000;
    W_ir[0][57] = 26'b11111111111110010101100110;
    W_ir[0][58] = 26'b11111111111110101101100110;
    W_ir[0][59] = 26'b00000000000010000111111111;
    W_ir[0][60] = 26'b11111111111101010100000101;
    W_ir[0][61] = 26'b11111111111100110111101111;
    W_ir[0][62] = 26'b11111111111100110001111110;
    W_ir[0][63] = 26'b00000000000010000101110100;
    W_ir[1][0] = 26'b11111111111110001011100101;
    W_ir[1][1] = 26'b11111111111110011001011110;
    W_ir[1][2] = 26'b00000000000010111111010101;
    W_ir[1][3] = 26'b00000000000010010110010001;
    W_ir[1][4] = 26'b00000000000000010100010110;
    W_ir[1][5] = 26'b00000000000000111110001011;
    W_ir[1][6] = 26'b00000000000000110100100011;
    W_ir[1][7] = 26'b00000000000000100000111100;
    W_ir[1][8] = 26'b00000000000000101000000110;
    W_ir[1][9] = 26'b00000000000000100101000110;
    W_ir[1][10] = 26'b11111111111111100001110010;
    W_ir[1][11] = 26'b11111111111111111110110000;
    W_ir[1][12] = 26'b00000000000000101110101111;
    W_ir[1][13] = 26'b00000000000001110000000010;
    W_ir[1][14] = 26'b11111111111101010110100001;
    W_ir[1][15] = 26'b00000000000000100010000110;
    W_ir[1][16] = 26'b11111111111111111111010101;
    W_ir[1][17] = 26'b11111111111111111100011011;
    W_ir[1][18] = 26'b11111111111111110010001110;
    W_ir[1][19] = 26'b11111111111110101111110011;
    W_ir[1][20] = 26'b11111111111111110000001110;
    W_ir[1][21] = 26'b00000000000000101101101100;
    W_ir[1][22] = 26'b11111111111111000000000101;
    W_ir[1][23] = 26'b11111111111110100000000011;
    W_ir[1][24] = 26'b00000000000000000001010010;
    W_ir[1][25] = 26'b00000000000010111010010000;
    W_ir[1][26] = 26'b11111111111100110010100110;
    W_ir[1][27] = 26'b11111111111100111010100001;
    W_ir[1][28] = 26'b00000000000011010110011111;
    W_ir[1][29] = 26'b00000000000001000001001111;
    W_ir[1][30] = 26'b00000000000000001110100011;
    W_ir[1][31] = 26'b11111111111111111101101000;
    W_ir[1][32] = 26'b11111111111110000101001001;
    W_ir[1][33] = 26'b11111111111111110100011111;
    W_ir[1][34] = 26'b11111111111111101101010000;
    W_ir[1][35] = 26'b00000000000000001111000011;
    W_ir[1][36] = 26'b00000000000000111110110001;
    W_ir[1][37] = 26'b00000000000000100100010101;
    W_ir[1][38] = 26'b00000000000000110010010010;
    W_ir[1][39] = 26'b00000000000010000000010101;
    W_ir[1][40] = 26'b00000000000001001101001111;
    W_ir[1][41] = 26'b00000000000000000001100100;
    W_ir[1][42] = 26'b11111111111111110101010000;
    W_ir[1][43] = 26'b00000000000001000000110101;
    W_ir[1][44] = 26'b00000000000000011000101010;
    W_ir[1][45] = 26'b00000000000000110010011110;
    W_ir[1][46] = 26'b11111111111111110011101111;
    W_ir[1][47] = 26'b11111111111111011100010110;
    W_ir[1][48] = 26'b11111111111111011011011100;
    W_ir[1][49] = 26'b11111111111100101011101001;
    W_ir[1][50] = 26'b00000000000001111010010100;
    W_ir[1][51] = 26'b00000000000010101010101011;
    W_ir[1][52] = 26'b11111111111111001110000110;
    W_ir[1][53] = 26'b11111111111110011101101001;
    W_ir[1][54] = 26'b11111111111110100000000001;
    W_ir[1][55] = 26'b11111111111110010011011010;
    W_ir[1][56] = 26'b11111111111111000001100011;
    W_ir[1][57] = 26'b00000000000011001011011010;
    W_ir[1][58] = 26'b00000000000001110111010000;
    W_ir[1][59] = 26'b11111111111101111100010111;
    W_ir[1][60] = 26'b11111111111111011110011011;
    W_ir[1][61] = 26'b11111111111111001001101000;
    W_ir[1][62] = 26'b00000000000010101100001010;
    W_ir[1][63] = 26'b11111111111110011110111110;
    W_ir[2][0] = 26'b11111111111110100100011111;
    W_ir[2][1] = 26'b11111111111111000000011100;
    W_ir[2][2] = 26'b11111111111100100110000011;
    W_ir[2][3] = 26'b11111111111101111000110111;
    W_ir[2][4] = 26'b11111111111110110101100100;
    W_ir[2][5] = 26'b11111111111111011101011011;
    W_ir[2][6] = 26'b00000000000000010111100001;
    W_ir[2][7] = 26'b11111111111101011101100010;
    W_ir[2][8] = 26'b11111111111111010100001101;
    W_ir[2][9] = 26'b11111111111111010110000101;
    W_ir[2][10] = 26'b11111111111111010000011101;
    W_ir[2][11] = 26'b11111111111100010110011101;
    W_ir[2][12] = 26'b11111111111111011010111101;
    W_ir[2][13] = 26'b00000000000000110111100010;
    W_ir[2][14] = 26'b11111111111111010100001001;
    W_ir[2][15] = 26'b00000000000001010111110110;
    W_ir[2][16] = 26'b11111111111101011001111110;
    W_ir[2][17] = 26'b00000000000011100101011000;
    W_ir[2][18] = 26'b00000000000000001100000001;
    W_ir[2][19] = 26'b00000000000001001011110100;
    W_ir[2][20] = 26'b00000000000000110111101110;
    W_ir[2][21] = 26'b11111111111110110111111000;
    W_ir[2][22] = 26'b00000000000001110111110011;
    W_ir[2][23] = 26'b00000000000011010011111011;
    W_ir[2][24] = 26'b00000000000001101100000010;
    W_ir[2][25] = 26'b00000000000000100011010011;
    W_ir[2][26] = 26'b11111111111111110000001111;
    W_ir[2][27] = 26'b11111111111100101101101100;
    W_ir[2][28] = 26'b11111111111111000011110001;
    W_ir[2][29] = 26'b00000000000011110001010100;
    W_ir[2][30] = 26'b11111111111110011111111010;
    W_ir[2][31] = 26'b11111111111110100001000010;
    W_ir[2][32] = 26'b00000000000000001010110100;
    W_ir[2][33] = 26'b00000000000001011011110101;
    W_ir[2][34] = 26'b11111111111111010001001101;
    W_ir[2][35] = 26'b11111111111111001001110111;
    W_ir[2][36] = 26'b00000000000000001100001111;
    W_ir[2][37] = 26'b00000000000000101010010111;
    W_ir[2][38] = 26'b00000000000010000000001100;
    W_ir[2][39] = 26'b11111111111111111110101010;
    W_ir[2][40] = 26'b00000000000001110001111000;
    W_ir[2][41] = 26'b11111111111111001010101010;
    W_ir[2][42] = 26'b00000000000001110110010111;
    W_ir[2][43] = 26'b11111111111111110011001010;
    W_ir[2][44] = 26'b00000000000000101100111111;
    W_ir[2][45] = 26'b00000000000000111111010011;
    W_ir[2][46] = 26'b00000000000000110001111000;
    W_ir[2][47] = 26'b00000000000000011001111101;
    W_ir[2][48] = 26'b00000000000000110011100010;
    W_ir[2][49] = 26'b00000000000000101011010101;
    W_ir[2][50] = 26'b11111111111110000101111111;
    W_ir[2][51] = 26'b00000000000001010111000001;
    W_ir[2][52] = 26'b00000000000001010001111110;
    W_ir[2][53] = 26'b00000000000000111001000101;
    W_ir[2][54] = 26'b11111111111100100101001000;
    W_ir[2][55] = 26'b00000000000001001011001000;
    W_ir[2][56] = 26'b00000000000000110010000111;
    W_ir[2][57] = 26'b11111111111101011100111010;
    W_ir[2][58] = 26'b11111111111110000111101110;
    W_ir[2][59] = 26'b11111111111110010110010101;
    W_ir[2][60] = 26'b00000000000010011001011000;
    W_ir[2][61] = 26'b00000000000001000110001101;
    W_ir[2][62] = 26'b00000000000010011111001000;
    W_ir[2][63] = 26'b00000000000100011010010100;
    W_ir[3][0] = 26'b11111111111111110111011110;
    W_ir[3][1] = 26'b00000000000011111101100001;
    W_ir[3][2] = 26'b00000000000000000000100000;
    W_ir[3][3] = 26'b00000000000011001010011110;
    W_ir[3][4] = 26'b11111111111101001000000010;
    W_ir[3][5] = 26'b00000000000000101001011000;
    W_ir[3][6] = 26'b00000000000000011110100000;
    W_ir[3][7] = 26'b11111111111110110011010110;
    W_ir[3][8] = 26'b11111111111111100011001101;
    W_ir[3][9] = 26'b00000000000010100110101101;
    W_ir[3][10] = 26'b11111111111110001001101000;
    W_ir[3][11] = 26'b11111111111111101001111110;
    W_ir[3][12] = 26'b11111111111101111110100110;
    W_ir[3][13] = 26'b11111111111111010100101010;
    W_ir[3][14] = 26'b11111111111111000111101011;
    W_ir[3][15] = 26'b11111111111111100011000101;
    W_ir[3][16] = 26'b00000000000000001001101100;
    W_ir[3][17] = 26'b00000000000000101010110110;
    W_ir[3][18] = 26'b11111111111110100111000111;
    W_ir[3][19] = 26'b00000000000010000001111100;
    W_ir[3][20] = 26'b11111111111111001100000011;
    W_ir[3][21] = 26'b00000000000000110011010100;
    W_ir[3][22] = 26'b00000000000001010100011010;
    W_ir[3][23] = 26'b00000000000000110110011111;
    W_ir[3][24] = 26'b00000000000011010100010011;
    W_ir[3][25] = 26'b00000000000000101110100101;
    W_ir[3][26] = 26'b11111111111111100010000100;
    W_ir[3][27] = 26'b11111111111110110010101011;
    W_ir[3][28] = 26'b00000000000000101101010001;
    W_ir[3][29] = 26'b00000000000000100110001010;
    W_ir[3][30] = 26'b11111111111101111000000011;
    W_ir[3][31] = 26'b00000000000100001000111101;
    W_ir[3][32] = 26'b00000000000010000111110010;
    W_ir[3][33] = 26'b11111111111101100010011101;
    W_ir[3][34] = 26'b00000000000001000000001100;
    W_ir[3][35] = 26'b00000000000000100100110100;
    W_ir[3][36] = 26'b00000000000000101110111111;
    W_ir[3][37] = 26'b11111111111100011111101010;
    W_ir[3][38] = 26'b00000000000001100010010000;
    W_ir[3][39] = 26'b00000000000000001110011010;
    W_ir[3][40] = 26'b11111111111111111011010001;
    W_ir[3][41] = 26'b00000000000010010101010100;
    W_ir[3][42] = 26'b11111111111101011000110011;
    W_ir[3][43] = 26'b00000000000000011000001110;
    W_ir[3][44] = 26'b11111111111110100111111100;
    W_ir[3][45] = 26'b11111111111110111000100101;
    W_ir[3][46] = 26'b00000000000011000101110111;
    W_ir[3][47] = 26'b11111111111110100011100010;
    W_ir[3][48] = 26'b11111111111111001010000110;
    W_ir[3][49] = 26'b11111111111111011001100010;
    W_ir[3][50] = 26'b11111111111110001111111010;
    W_ir[3][51] = 26'b11111111111110100000010011;
    W_ir[3][52] = 26'b11111111111110010111100111;
    W_ir[3][53] = 26'b11111111111110001011010010;
    W_ir[3][54] = 26'b11111111111110111101100001;
    W_ir[3][55] = 26'b11111111111100011000001000;
    W_ir[3][56] = 26'b11111111111110010011001000;
    W_ir[3][57] = 26'b00000000000001111100111001;
    W_ir[3][58] = 26'b11111111111101110011100010;
    W_ir[3][59] = 26'b11111111111110011100011110;
    W_ir[3][60] = 26'b11111111111110011111111101;
    W_ir[3][61] = 26'b11111111111110101101010110;
    W_ir[3][62] = 26'b11111111111101000001000110;
    W_ir[3][63] = 26'b11111111111110110000001010;
    W_ir[4][0] = 26'b11111111111111110010000001;
    W_ir[4][1] = 26'b11111111111111001101101000;
    W_ir[4][2] = 26'b11111111111111011010110110;
    W_ir[4][3] = 26'b11111111111110011100111100;
    W_ir[4][4] = 26'b00000000000000000101000010;
    W_ir[4][5] = 26'b00000000000001011100011001;
    W_ir[4][6] = 26'b11111111111110001101011110;
    W_ir[4][7] = 26'b11111111111101011101000111;
    W_ir[4][8] = 26'b11111111111100010100000010;
    W_ir[4][9] = 26'b11111111111110100101100101;
    W_ir[4][10] = 26'b11111111111100101110000101;
    W_ir[4][11] = 26'b11111111111110111100001000;
    W_ir[4][12] = 26'b11111111111111011010011000;
    W_ir[4][13] = 26'b00000000000001011100001011;
    W_ir[4][14] = 26'b00000000000000011001001001;
    W_ir[4][15] = 26'b11111111111111011010010100;
    W_ir[4][16] = 26'b11111111111110000011001110;
    W_ir[4][17] = 26'b11111111111110100010010111;
    W_ir[4][18] = 26'b11111111111110000110011001;
    W_ir[4][19] = 26'b11111111111101101010011010;
    W_ir[4][20] = 26'b11111111111111011100100001;
    W_ir[4][21] = 26'b00000000000001101011001101;
    W_ir[4][22] = 26'b00000000000100001110110100;
    W_ir[4][23] = 26'b00000000000010010101111110;
    W_ir[4][24] = 26'b11111111111100100000100101;
    W_ir[4][25] = 26'b11111111111101001011010011;
    W_ir[4][26] = 26'b00000000000000001110100110;
    W_ir[4][27] = 26'b11111111111100100000010111;
    W_ir[4][28] = 26'b00000000000010111110010001;
    W_ir[4][29] = 26'b11111111111111110110101110;
    W_ir[4][30] = 26'b00000000000010110101110111;
    W_ir[4][31] = 26'b11111111111110000100100100;
    W_ir[4][32] = 26'b11111111111100101111111111;
    W_ir[4][33] = 26'b11111111111101001010101110;
    W_ir[4][34] = 26'b11111111111110000110001111;
    W_ir[4][35] = 26'b11111111111101111011100100;
    W_ir[4][36] = 26'b11111111111100110110011101;
    W_ir[4][37] = 26'b11111111111101010101011100;
    W_ir[4][38] = 26'b11111111111110010010000110;
    W_ir[4][39] = 26'b00000000000001000100110110;
    W_ir[4][40] = 26'b00000000000000101111111011;
    W_ir[4][41] = 26'b11111111111110001100011101;
    W_ir[4][42] = 26'b11111111111111101111100111;
    W_ir[4][43] = 26'b11111111111110100111101001;
    W_ir[4][44] = 26'b11111111111100001000111000;
    W_ir[4][45] = 26'b11111111111111010101111011;
    W_ir[4][46] = 26'b11111111111111010101001001;
    W_ir[4][47] = 26'b11111111111111100001011001;
    W_ir[4][48] = 26'b00000000000000000000100110;
    W_ir[4][49] = 26'b11111111111111001001110110;
    W_ir[4][50] = 26'b00000000000010100111001011;
    W_ir[4][51] = 26'b11111111111110011011111001;
    W_ir[4][52] = 26'b00000000000011101010001011;
    W_ir[4][53] = 26'b00000000000001110001010000;
    W_ir[4][54] = 26'b00000000000011110110001001;
    W_ir[4][55] = 26'b00000000000011001101011001;
    W_ir[4][56] = 26'b00000000000001010000010001;
    W_ir[4][57] = 26'b11111111111100100001110111;
    W_ir[4][58] = 26'b00000000000010000011010101;
    W_ir[4][59] = 26'b00000000000110111011010000;
    W_ir[4][60] = 26'b00000000000101001011001100;
    W_ir[4][61] = 26'b00000000000101011101011000;
    W_ir[4][62] = 26'b00000000000110011100100010;
    W_ir[4][63] = 26'b00000000000101110000001010;
    W_ir[5][0] = 26'b00000000000000101010000111;
    W_ir[5][1] = 26'b00000000000000101101010100;
    W_ir[5][2] = 26'b00000000000000110101100001;
    W_ir[5][3] = 26'b11111111111111100000111000;
    W_ir[5][4] = 26'b11111111111111011101011111;
    W_ir[5][5] = 26'b11111111111101101100001000;
    W_ir[5][6] = 26'b00000000000011000111010101;
    W_ir[5][7] = 26'b11111111111100010101001110;
    W_ir[5][8] = 26'b11111111111101001001110110;
    W_ir[5][9] = 26'b11111111111110111101100010;
    W_ir[5][10] = 26'b11111111111111111010100011;
    W_ir[5][11] = 26'b11111111111111011010011110;
    W_ir[5][12] = 26'b11111111111101110000101010;
    W_ir[5][13] = 26'b11111111111111010110000100;
    W_ir[5][14] = 26'b11111111111110000011110001;
    W_ir[5][15] = 26'b11111111111101111111011000;
    W_ir[5][16] = 26'b00000000000010010011111000;
    W_ir[5][17] = 26'b11111111111101011111000101;
    W_ir[5][18] = 26'b00000000000000011110111101;
    W_ir[5][19] = 26'b11111111111100110111101110;
    W_ir[5][20] = 26'b11111111111111011000000100;
    W_ir[5][21] = 26'b00000000000000000101011010;
    W_ir[5][22] = 26'b00000000000001010010011110;
    W_ir[5][23] = 26'b00000000000000110011011011;
    W_ir[5][24] = 26'b11111111111111101011111101;
    W_ir[5][25] = 26'b11111111111110011110011011;
    W_ir[5][26] = 26'b11111111111111101100111100;
    W_ir[5][27] = 26'b00000000000001011100110100;
    W_ir[5][28] = 26'b00000000000000010100000001;
    W_ir[5][29] = 26'b11111111111110001010000010;
    W_ir[5][30] = 26'b11111111111111000100001110;
    W_ir[5][31] = 26'b11111111111100100010000100;
    W_ir[5][32] = 26'b11111111111111110001011001;
    W_ir[5][33] = 26'b11111111111100000000010010;
    W_ir[5][34] = 26'b11111111111110111111011000;
    W_ir[5][35] = 26'b00000000000001111100100101;
    W_ir[5][36] = 26'b11111111111110000001111110;
    W_ir[5][37] = 26'b11111111111101000100011101;
    W_ir[5][38] = 26'b11111111111011101001010010;
    W_ir[5][39] = 26'b00000000000010100011011110;
    W_ir[5][40] = 26'b11111111111110101110101000;
    W_ir[5][41] = 26'b11111111111111011111111101;
    W_ir[5][42] = 26'b00000000000000001101101101;
    W_ir[5][43] = 26'b11111111111110100110001100;
    W_ir[5][44] = 26'b00000000000000100001000111;
    W_ir[5][45] = 26'b11111111111110101001111111;
    W_ir[5][46] = 26'b11111111111111011011001100;
    W_ir[5][47] = 26'b00000000000001111010001001;
    W_ir[5][48] = 26'b00000000000000111100110111;
    W_ir[5][49] = 26'b00000000000000110010000100;
    W_ir[5][50] = 26'b00000000000000101010101010;
    W_ir[5][51] = 26'b00000000000000101100011101;
    W_ir[5][52] = 26'b11111111111110111011001001;
    W_ir[5][53] = 26'b11111111111110101101110111;
    W_ir[5][54] = 26'b00000000000000111010100100;
    W_ir[5][55] = 26'b00000000000000000000101010;
    W_ir[5][56] = 26'b00000000000000101100001011;
    W_ir[5][57] = 26'b11111111111101101111011110;
    W_ir[5][58] = 26'b11111111111101111001100110;
    W_ir[5][59] = 26'b11111111111110110110001001;
    W_ir[5][60] = 26'b00000000000011101110101010;
    W_ir[5][61] = 26'b00000000000010100001110101;
    W_ir[5][62] = 26'b11111111111110110000001100;
    W_ir[5][63] = 26'b00000000000010010000110110;
    W_ir[6][0] = 26'b00000000000010111010101011;
    W_ir[6][1] = 26'b11111111111111001110101111;
    W_ir[6][2] = 26'b00000000000100101011010000;
    W_ir[6][3] = 26'b11111111111110110011011101;
    W_ir[6][4] = 26'b00000000000010100111110011;
    W_ir[6][5] = 26'b00000000000000100111010110;
    W_ir[6][6] = 26'b11111111111100101100000111;
    W_ir[6][7] = 26'b00000000000100101100001101;
    W_ir[6][8] = 26'b00000000000101011000111110;
    W_ir[6][9] = 26'b00000000000011001010011111;
    W_ir[6][10] = 26'b00000000000011110110101100;
    W_ir[6][11] = 26'b11111111111111111010000001;
    W_ir[6][12] = 26'b00000000000000000011010001;
    W_ir[6][13] = 26'b00000000000001001010011001;
    W_ir[6][14] = 26'b11111111111110110111110100;
    W_ir[6][15] = 26'b11111111111100101110000111;
    W_ir[6][16] = 26'b11111111111110101001000111;
    W_ir[6][17] = 26'b00000000000010011101100000;
    W_ir[6][18] = 26'b11111111111111111010010001;
    W_ir[6][19] = 26'b11111111111111110100101100;
    W_ir[6][20] = 26'b11111111111111010001011000;
    W_ir[6][21] = 26'b11111111111101010101011001;
    W_ir[6][22] = 26'b00000000000100010110000011;
    W_ir[6][23] = 26'b11111111111111110101110100;
    W_ir[6][24] = 26'b11111111111101011101001010;
    W_ir[6][25] = 26'b00000000000001010000101100;
    W_ir[6][26] = 26'b11111111111101001111000100;
    W_ir[6][27] = 26'b11111111111101111000000010;
    W_ir[6][28] = 26'b00000000000011000011010010;
    W_ir[6][29] = 26'b00000000000010101000111011;
    W_ir[6][30] = 26'b11111111111101011000001111;
    W_ir[6][31] = 26'b00000000000010011001111111;
    W_ir[6][32] = 26'b00000000000000001101011100;
    W_ir[6][33] = 26'b00000000000001010000110010;
    W_ir[6][34] = 26'b00000000000011010110101011;
    W_ir[6][35] = 26'b00000000000100000001010000;
    W_ir[6][36] = 26'b11111111111111101100010001;
    W_ir[6][37] = 26'b00000000000000111110101110;
    W_ir[6][38] = 26'b11111111111100000101101011;
    W_ir[6][39] = 26'b11111111111111100110101101;
    W_ir[6][40] = 26'b00000000000001111111101000;
    W_ir[6][41] = 26'b11111111111110011101111111;
    W_ir[6][42] = 26'b00000000000100011011110001;
    W_ir[6][43] = 26'b00000000000001000011110111;
    W_ir[6][44] = 26'b00000000000010001000010001;
    W_ir[6][45] = 26'b11111111111110001010001111;
    W_ir[6][46] = 26'b11111111111100101110011001;
    W_ir[6][47] = 26'b00000000000011111111110000;
    W_ir[6][48] = 26'b11111111111101000000100001;
    W_ir[6][49] = 26'b11111111111110001001000011;
    W_ir[6][50] = 26'b00000000000010000000110001;
    W_ir[6][51] = 26'b11111111111111101101011001;
    W_ir[6][52] = 26'b00000000000010001000001110;
    W_ir[6][53] = 26'b11111111111001001011110000;
    W_ir[6][54] = 26'b11111111111111000101010110;
    W_ir[6][55] = 26'b00000000000000100110010010;
    W_ir[6][56] = 26'b11111111111101100101010011;
    W_ir[6][57] = 26'b11111111111110111000010100;
    W_ir[6][58] = 26'b11111111111101011100000011;
    W_ir[6][59] = 26'b11111111111101000001111101;
    W_ir[6][60] = 26'b11111111111111000101011100;
    W_ir[6][61] = 26'b11111111111001110111111000;
    W_ir[6][62] = 26'b11111111111000100111111011;
    W_ir[6][63] = 26'b11111111111000001011111000;
    W_ir[7][0] = 26'b11111111111010100101000101;
    W_ir[7][1] = 26'b11111111111010011000010011;
    W_ir[7][2] = 26'b00000000000001100011101001;
    W_ir[7][3] = 26'b11111111111111001100010011;
    W_ir[7][4] = 26'b00000000000011000110100010;
    W_ir[7][5] = 26'b00000000000100001111001011;
    W_ir[7][6] = 26'b11111111111100100101011000;
    W_ir[7][7] = 26'b00000000000000110100001001;
    W_ir[7][8] = 26'b11111111111101011101100010;
    W_ir[7][9] = 26'b11111111111001110010100100;
    W_ir[7][10] = 26'b11111111111101110111010100;
    W_ir[7][11] = 26'b00000000000010011110010110;
    W_ir[7][12] = 26'b00000000000010111111000111;
    W_ir[7][13] = 26'b11111111111101001101010100;
    W_ir[7][14] = 26'b00000000000011000001110011;
    W_ir[7][15] = 26'b11111111111111111111011001;
    W_ir[7][16] = 26'b00000000000000100111100110;
    W_ir[7][17] = 26'b11111111111110011111111101;
    W_ir[7][18] = 26'b00000000000000100110111101;
    W_ir[7][19] = 26'b00000000000011101011001011;
    W_ir[7][20] = 26'b11111111111110001111101111;
    W_ir[7][21] = 26'b11111111111110100010011001;
    W_ir[7][22] = 26'b00000000000011111101010101;
    W_ir[7][23] = 26'b11111111111110010100110100;
    W_ir[7][24] = 26'b00000000000011100100001111;
    W_ir[7][25] = 26'b00000000000001101110001100;
    W_ir[7][26] = 26'b00000000000010001010100010;
    W_ir[7][27] = 26'b11111111111111000111000010;
    W_ir[7][28] = 26'b00000000000010110101010000;
    W_ir[7][29] = 26'b00000000000100010000111110;
    W_ir[7][30] = 26'b00000000000010110010010001;
    W_ir[7][31] = 26'b00000000000001011111110010;
    W_ir[7][32] = 26'b11111111111101011100110010;
    W_ir[7][33] = 26'b11111111111110011101100110;
    W_ir[7][34] = 26'b11111111111010001110110110;
    W_ir[7][35] = 26'b11111111111100110100101001;
    W_ir[7][36] = 26'b00000000000011110010010010;
    W_ir[7][37] = 26'b00000000000000000010001101;
    W_ir[7][38] = 26'b00000000000011001100111110;
    W_ir[7][39] = 26'b11111111111011101111101011;
    W_ir[7][40] = 26'b11111111111111110110110001;
    W_ir[7][41] = 26'b11111111111011110111111001;
    W_ir[7][42] = 26'b11111111111011100110100100;
    W_ir[7][43] = 26'b11111111111011011100000110;
    W_ir[7][44] = 26'b11111111111101101010000110;
    W_ir[7][45] = 26'b00000000000000100110011110;
    W_ir[7][46] = 26'b00000000001000110000011011;
    W_ir[7][47] = 26'b11111111111101101001010101;
    W_ir[7][48] = 26'b11111111111111100110110011;
    W_ir[7][49] = 26'b11111111111101011001110101;
    W_ir[7][50] = 26'b11111111111100001001111100;
    W_ir[7][51] = 26'b00000000000101110110001100;
    W_ir[7][52] = 26'b11111111111011101001101110;
    W_ir[7][53] = 26'b00000000000001011000101100;
    W_ir[7][54] = 26'b00000000000100011011111011;
    W_ir[7][55] = 26'b00000000000000101101000100;
    W_ir[7][56] = 26'b00000000001001000101101110;
    W_ir[7][57] = 26'b00000000000001001001101001;
    W_ir[7][58] = 26'b00000000001001010001010100;
    W_ir[7][59] = 26'b00000000000001011110100011;
    W_ir[7][60] = 26'b11111111111100001001110101;
    W_ir[7][61] = 26'b00000000000100011100000101;
    W_ir[7][62] = 26'b00000000000110000001100100;
    W_ir[7][63] = 26'b11111111111100001001111000;
    W_ir[8][0] = 26'b11111111111110001110100011;
    W_ir[8][1] = 26'b00000000000000111101111100;
    W_ir[8][2] = 26'b11111111111111001100010000;
    W_ir[8][3] = 26'b00000000000010001101110100;
    W_ir[8][4] = 26'b11111111111111011001001100;
    W_ir[8][5] = 26'b11111111111110111001011101;
    W_ir[8][6] = 26'b11111111111100100000000111;
    W_ir[8][7] = 26'b11111111111110000110100000;
    W_ir[8][8] = 26'b11111111111110111010010110;
    W_ir[8][9] = 26'b00000000000010010110010110;
    W_ir[8][10] = 26'b00000000000001000101101010;
    W_ir[8][11] = 26'b00000000000011011101110110;
    W_ir[8][12] = 26'b11111111111111000100010000;
    W_ir[8][13] = 26'b00000000000001110011000110;
    W_ir[8][14] = 26'b00000000000001110001111010;
    W_ir[8][15] = 26'b00000000000000110000101010;
    W_ir[8][16] = 26'b11111111111111010110011010;
    W_ir[8][17] = 26'b00000000000010101110101111;
    W_ir[8][18] = 26'b00000000000011111111000010;
    W_ir[8][19] = 26'b00000000000010001101110110;
    W_ir[8][20] = 26'b11111111111111100110101111;
    W_ir[8][21] = 26'b00000000000000101110110100;
    W_ir[8][22] = 26'b00000000000010110001101110;
    W_ir[8][23] = 26'b00000000000000101000000010;
    W_ir[8][24] = 26'b00000000000000001111011101;
    W_ir[8][25] = 26'b11111111111111010100011000;
    W_ir[8][26] = 26'b11111111111100010011001011;
    W_ir[8][27] = 26'b00000000000000110101111110;
    W_ir[8][28] = 26'b00000000000001111100110010;
    W_ir[8][29] = 26'b00000000000000001010111011;
    W_ir[8][30] = 26'b00000000000010011110011010;
    W_ir[8][31] = 26'b00000000000010000111010100;
    W_ir[8][32] = 26'b11111111111111011011000101;
    W_ir[8][33] = 26'b11111111111101101111100111;
    W_ir[8][34] = 26'b11111111111100111000000100;
    W_ir[8][35] = 26'b11111111111110011101101011;
    W_ir[8][36] = 26'b11111111111110010001001110;
    W_ir[8][37] = 26'b11111111111010110100100100;
    W_ir[8][38] = 26'b00000000000000111000111111;
    W_ir[8][39] = 26'b11111111111111101110010000;
    W_ir[8][40] = 26'b11111111111111010010111011;
    W_ir[8][41] = 26'b00000000000011011010111011;
    W_ir[8][42] = 26'b11111111111101010111001111;
    W_ir[8][43] = 26'b00000000000010001010111000;
    W_ir[8][44] = 26'b00000000000000000001011110;
    W_ir[8][45] = 26'b11111111111110000001111011;
    W_ir[8][46] = 26'b11111111111101101010011100;
    W_ir[8][47] = 26'b00000000000010101011101110;
    W_ir[8][48] = 26'b00000000000001000110010011;
    W_ir[8][49] = 26'b00000000000100101110100101;
    W_ir[8][50] = 26'b11111111111111111111000110;
    W_ir[8][51] = 26'b00000000000000111101101001;
    W_ir[8][52] = 26'b11111111111110110101000101;
    W_ir[8][53] = 26'b11111111111101000111100011;
    W_ir[8][54] = 26'b11111111111100101100100011;
    W_ir[8][55] = 26'b11111111111110010110111011;
    W_ir[8][56] = 26'b00000000000011101100000001;
    W_ir[8][57] = 26'b11111111111110110100110100;
    W_ir[8][58] = 26'b00000000000011110011100011;
    W_ir[8][59] = 26'b11111111111111001000010111;
    W_ir[8][60] = 26'b11111111111011101000101001;
    W_ir[8][61] = 26'b11111111111001000111111100;
    W_ir[8][62] = 26'b11111111111000000011011110;
    W_ir[8][63] = 26'b00000000000001101111011100;
    W_ir[9][0] = 26'b00000000000011001011001011;
    W_ir[9][1] = 26'b00000000000001000110010100;
    W_ir[9][2] = 26'b00000000000000101101100111;
    W_ir[9][3] = 26'b00000000000000000011001001;
    W_ir[9][4] = 26'b00000000000000011110111010;
    W_ir[9][5] = 26'b00000000000010011010001010;
    W_ir[9][6] = 26'b11111111111100110100011101;
    W_ir[9][7] = 26'b11111111111101011010001101;
    W_ir[9][8] = 26'b00000000000000000100111010;
    W_ir[9][9] = 26'b00000000000100000010001010;
    W_ir[9][10] = 26'b00000000000010000100111110;
    W_ir[9][11] = 26'b11111111111011110010010001;
    W_ir[9][12] = 26'b11111111111101011011110011;
    W_ir[9][13] = 26'b00000000000010101110000101;
    W_ir[9][14] = 26'b11111111111111001010110010;
    W_ir[9][15] = 26'b00000000000011001101001011;
    W_ir[9][16] = 26'b11111111111100001110001001;
    W_ir[9][17] = 26'b00000000000001110110101110;
    W_ir[9][18] = 26'b00000000000100100010000101;
    W_ir[9][19] = 26'b11111111111101010000110110;
    W_ir[9][20] = 26'b11111111111101100110010111;
    W_ir[9][21] = 26'b11111111111100010000011111;
    W_ir[9][22] = 26'b00000000000010001101100001;
    W_ir[9][23] = 26'b00000000000101001111010111;
    W_ir[9][24] = 26'b00000000000001111011111000;
    W_ir[9][25] = 26'b11111111111110000101010011;
    W_ir[9][26] = 26'b11111111111110011000000111;
    W_ir[9][27] = 26'b11111111111101111010111001;
    W_ir[9][28] = 26'b11111111111110101001110010;
    W_ir[9][29] = 26'b11111111111100110110000111;
    W_ir[9][30] = 26'b11111111111111000111010000;
    W_ir[9][31] = 26'b11111111111100110011011011;
    W_ir[9][32] = 26'b00000000000010011100111000;
    W_ir[9][33] = 26'b11111111111110111110010111;
    W_ir[9][34] = 26'b11111111111101111110001100;
    W_ir[9][35] = 26'b00000000000010100101101001;
    W_ir[9][36] = 26'b11111111111011011011011111;
    W_ir[9][37] = 26'b00000000000000101001110101;
    W_ir[9][38] = 26'b11111111111111111000110010;
    W_ir[9][39] = 26'b11111111111101111110000000;
    W_ir[9][40] = 26'b00000000000010110110011011;
    W_ir[9][41] = 26'b00000000000001011011111100;
    W_ir[9][42] = 26'b00000000000011101111110000;
    W_ir[9][43] = 26'b00000000000011001101101111;
    W_ir[9][44] = 26'b00000000000000001100010111;
    W_ir[9][45] = 26'b00000000000011101010100001;
    W_ir[9][46] = 26'b00000000000001000001010000;
    W_ir[9][47] = 26'b11111111111111001001011100;
    W_ir[9][48] = 26'b11111111111101000101000100;
    W_ir[9][49] = 26'b11111111111111011010111110;
    W_ir[9][50] = 26'b11111111111110010100101101;
    W_ir[9][51] = 26'b00000000000001110100100011;
    W_ir[9][52] = 26'b00000000000010101110000101;
    W_ir[9][53] = 26'b00000000000001100010000010;
    W_ir[9][54] = 26'b11111111111100001011111111;
    W_ir[9][55] = 26'b00000000000100110010111100;
    W_ir[9][56] = 26'b00000000000010011010001101;
    W_ir[9][57] = 26'b11111111111111000010100101;
    W_ir[9][58] = 26'b11111111111111101101111110;
    W_ir[9][59] = 26'b00000000000011011111000010;
    W_ir[9][60] = 26'b11111111111011101110001111;
    W_ir[9][61] = 26'b11111111111111110011001001;
    W_ir[9][62] = 26'b11111111111110010010000011;
    W_ir[9][63] = 26'b11111111111110100000000111;
    W_ir[10][0] = 26'b00000000000001011011101000;
    W_ir[10][1] = 26'b00000000000001111110011000;
    W_ir[10][2] = 26'b11111111111111010000100000;
    W_ir[10][3] = 26'b00000000000000110001101001;
    W_ir[10][4] = 26'b00000000000011001101001101;
    W_ir[10][5] = 26'b00000000000001011001000111;
    W_ir[10][6] = 26'b11111111111011011001111100;
    W_ir[10][7] = 26'b00000000000001011100100011;
    W_ir[10][8] = 26'b11111111111010000011000101;
    W_ir[10][9] = 26'b11111111111111001100110111;
    W_ir[10][10] = 26'b11111111111111111011010111;
    W_ir[10][11] = 26'b11111111111110001111010101;
    W_ir[10][12] = 26'b11111111111100100001110101;
    W_ir[10][13] = 26'b00000000000001100100110110;
    W_ir[10][14] = 26'b11111111111111110010000101;
    W_ir[10][15] = 26'b11111111111010100110100111;
    W_ir[10][16] = 26'b00000000000010000100010011;
    W_ir[10][17] = 26'b00000000000010010100011110;
    W_ir[10][18] = 26'b11111111111010000100000010;
    W_ir[10][19] = 26'b11111111111011110011011000;
    W_ir[10][20] = 26'b00000000000011010011010011;
    W_ir[10][21] = 26'b11111111111100110111101000;
    W_ir[10][22] = 26'b00000000000001010110100000;
    W_ir[10][23] = 26'b11111111111101000001100010;
    W_ir[10][24] = 26'b00000000000001100101010001;
    W_ir[10][25] = 26'b11111111111101010011011100;
    W_ir[10][26] = 26'b00000000000100101011101000;
    W_ir[10][27] = 26'b11111111111111001111100111;
    W_ir[10][28] = 26'b00000000000010110011111101;
    W_ir[10][29] = 26'b00000000000100011011101011;
    W_ir[10][30] = 26'b11111111111111011000010001;
    W_ir[10][31] = 26'b00000000000000000001001010;
    W_ir[10][32] = 26'b00000000000101011011111011;
    W_ir[10][33] = 26'b11111111111011111001110010;
    W_ir[10][34] = 26'b11111111111100001011101101;
    W_ir[10][35] = 26'b11111111111110001011000000;
    W_ir[10][36] = 26'b00000000000101000010111001;
    W_ir[10][37] = 26'b00000000000100001011011101;
    W_ir[10][38] = 26'b11111111111101011010000111;
    W_ir[10][39] = 26'b11111111111010101110101100;
    W_ir[10][40] = 26'b00000000000010001101110001;
    W_ir[10][41] = 26'b11111111111111101100110101;
    W_ir[10][42] = 26'b11111111111100001110011010;
    W_ir[10][43] = 26'b00000000000000101100100000;
    W_ir[10][44] = 26'b11111111111110101101101100;
    W_ir[10][45] = 26'b00000000000010011001111110;
    W_ir[10][46] = 26'b11111111111111000111001111;
    W_ir[10][47] = 26'b11111111111111000110001101;
    W_ir[10][48] = 26'b11111111111110011111100100;
    W_ir[10][49] = 26'b11111111111111111100010100;
    W_ir[10][50] = 26'b11111111111100001110000101;
    W_ir[10][51] = 26'b11111111111110011010011110;
    W_ir[10][52] = 26'b11111111111011111011111011;
    W_ir[10][53] = 26'b00000000000011011010011011;
    W_ir[10][54] = 26'b11111111111111011111111010;
    W_ir[10][55] = 26'b11111111111110001110001000;
    W_ir[10][56] = 26'b11111111111110010010100100;
    W_ir[10][57] = 26'b00000000000011100110100100;
    W_ir[10][58] = 26'b00000000000011110111001010;
    W_ir[10][59] = 26'b00000000000100110110011110;
    W_ir[10][60] = 26'b00000000000111100101011010;
    W_ir[10][61] = 26'b00000000000101000101101000;
    W_ir[10][62] = 26'b00000000001000101110110110;
    W_ir[10][63] = 26'b00000000000110011110011110;
    W_ir[11][0] = 26'b11111111111010011000111100;
    W_ir[11][1] = 26'b00000000000100000101101011;
    W_ir[11][2] = 26'b00000000000000010011010110;
    W_ir[11][3] = 26'b00000000000100011011110010;
    W_ir[11][4] = 26'b11111111111010111001000111;
    W_ir[11][5] = 26'b00000000000001000110101110;
    W_ir[11][6] = 26'b11111111111011100001000110;
    W_ir[11][7] = 26'b00000000000010011110011111;
    W_ir[11][8] = 26'b11111111111001000110111001;
    W_ir[11][9] = 26'b11111111111010011000001111;
    W_ir[11][10] = 26'b00000000000100101000010100;
    W_ir[11][11] = 26'b11111111111010011000101011;
    W_ir[11][12] = 26'b11111111111010100011011100;
    W_ir[11][13] = 26'b00000000000010010100100010;
    W_ir[11][14] = 26'b00000000000001111110100100;
    W_ir[11][15] = 26'b00000000000001111111010000;
    W_ir[11][16] = 26'b00000000000101010100010001;
    W_ir[11][17] = 26'b11111111111110111000110110;
    W_ir[11][18] = 26'b11111111111111111110100111;
    W_ir[11][19] = 26'b00000000000110010110001100;
    W_ir[11][20] = 26'b11111111111111000001111100;
    W_ir[11][21] = 26'b11111111111100001110001100;
    W_ir[11][22] = 26'b11111111111110100101010101;
    W_ir[11][23] = 26'b11111111111110001011010100;
    W_ir[11][24] = 26'b11111111111011000010110001;
    W_ir[11][25] = 26'b11111111111111000101100011;
    W_ir[11][26] = 26'b11111111111011111101100111;
    W_ir[11][27] = 26'b11111111111010111111100110;
    W_ir[11][28] = 26'b00000000000110100110110010;
    W_ir[11][29] = 26'b00000000000010001101101001;
    W_ir[11][30] = 26'b00000000000000011001101000;
    W_ir[11][31] = 26'b00000000000011101010100011;
    W_ir[11][32] = 26'b00000000000010001001111100;
    W_ir[11][33] = 26'b11111111111111000000100100;
    W_ir[11][34] = 26'b00000000000011100100111101;
    W_ir[11][35] = 26'b00000000000001110011010000;
    W_ir[11][36] = 26'b11111111111011101111001000;
    W_ir[11][37] = 26'b11111111111010110110110111;
    W_ir[11][38] = 26'b00000000000010001001011100;
    W_ir[11][39] = 26'b11111111111111110100110110;
    W_ir[11][40] = 26'b11111111111010000010010101;
    W_ir[11][41] = 26'b11111111111010110011000110;
    W_ir[11][42] = 26'b00000000000100000101011001;
    W_ir[11][43] = 26'b00000000000000010111101011;
    W_ir[11][44] = 26'b00000000000001011000101011;
    W_ir[11][45] = 26'b00000000000110001110001011;
    W_ir[11][46] = 26'b11111111111111011011111101;
    W_ir[11][47] = 26'b00000000000101000000101000;
    W_ir[11][48] = 26'b00000000000000100110000000;
    W_ir[11][49] = 26'b11111111111111011010110100;
    W_ir[11][50] = 26'b11111111111101010011011110;
    W_ir[11][51] = 26'b00000000000010110011000101;
    W_ir[11][52] = 26'b11111111111110110000100011;
    W_ir[11][53] = 26'b11111111111010111100011101;
    W_ir[11][54] = 26'b00000000000110001000111110;
    W_ir[11][55] = 26'b00000000000000111100101001;
    W_ir[11][56] = 26'b11111111111101000110100001;
    W_ir[11][57] = 26'b00000000000010110101111011;
    W_ir[11][58] = 26'b11111111111101100111011111;
    W_ir[11][59] = 26'b00000000000101100010100110;
    W_ir[11][60] = 26'b00000000000101011101001011;
    W_ir[11][61] = 26'b00000000000001010011010000;
    W_ir[11][62] = 26'b00000000000000011100100101;
    W_ir[11][63] = 26'b00000000000100101111011110;
    W_ir[12][0] = 26'b00000000000001010010011110;
    W_ir[12][1] = 26'b00000000000010011100011000;
    W_ir[12][2] = 26'b00000000000001110111001110;
    W_ir[12][3] = 26'b00000000000010001100110010;
    W_ir[12][4] = 26'b11111111111110110100110100;
    W_ir[12][5] = 26'b11111111111101010101000001;
    W_ir[12][6] = 26'b00000000000001110011010001;
    W_ir[12][7] = 26'b00000000000000111101101110;
    W_ir[12][8] = 26'b11111111111100100000101110;
    W_ir[12][9] = 26'b00000000000000010110011000;
    W_ir[12][10] = 26'b00000000000011111010111111;
    W_ir[12][11] = 26'b11111111111111111110101100;
    W_ir[12][12] = 26'b00000000000010011111111001;
    W_ir[12][13] = 26'b00000000000000101100000000;
    W_ir[12][14] = 26'b00000000000000100111011101;
    W_ir[12][15] = 26'b00000000000010111001011010;
    W_ir[12][16] = 26'b11111111111111100000000101;
    W_ir[12][17] = 26'b00000000000011011100110111;
    W_ir[12][18] = 26'b11111111111111100011001001;
    W_ir[12][19] = 26'b00000000000010010001001011;
    W_ir[12][20] = 26'b11111111111111100001111100;
    W_ir[12][21] = 26'b00000000000010000111001000;
    W_ir[12][22] = 26'b00000000000001100001111111;
    W_ir[12][23] = 26'b00000000000001100011100000;
    W_ir[12][24] = 26'b11111111111101011110111110;
    W_ir[12][25] = 26'b00000000000001111000001100;
    W_ir[12][26] = 26'b00000000000010001011100110;
    W_ir[12][27] = 26'b00000000000001011011010101;
    W_ir[12][28] = 26'b00000000000011100010100110;
    W_ir[12][29] = 26'b11111111111100101100001011;
    W_ir[12][30] = 26'b11111111111110110101100001;
    W_ir[12][31] = 26'b00000000000001100111000001;
    W_ir[12][32] = 26'b00000000000000110001101110;
    W_ir[12][33] = 26'b00000000000001111010001100;
    W_ir[12][34] = 26'b00000000000001111010011110;
    W_ir[12][35] = 26'b00000000000000011010111101;
    W_ir[12][36] = 26'b00000000000011111110101101;
    W_ir[12][37] = 26'b00000000000001010001000000;
    W_ir[12][38] = 26'b11111111111110111011001110;
    W_ir[12][39] = 26'b00000000000000111101100110;
    W_ir[12][40] = 26'b00000000000010010101101000;
    W_ir[12][41] = 26'b11111111111101000000111011;
    W_ir[12][42] = 26'b00000000000000111100111010;
    W_ir[12][43] = 26'b11111111111110100001001011;
    W_ir[12][44] = 26'b11111111111111111001001101;
    W_ir[12][45] = 26'b11111111111101110010100010;
    W_ir[12][46] = 26'b11111111111100111001111111;
    W_ir[12][47] = 26'b00000000000011011110110000;
    W_ir[12][48] = 26'b11111111111111000101001111;
    W_ir[12][49] = 26'b11111111111110011100100001;
    W_ir[12][50] = 26'b11111111111111100110010101;
    W_ir[12][51] = 26'b00000000000000000001001000;
    W_ir[12][52] = 26'b11111111111100011011000001;
    W_ir[12][53] = 26'b11111111111110101001001010;
    W_ir[12][54] = 26'b00000000000001000011001101;
    W_ir[12][55] = 26'b11111111111110011111000000;
    W_ir[12][56] = 26'b00000000000010011001010000;
    W_ir[12][57] = 26'b11111111111110010101100110;
    W_ir[12][58] = 26'b11111111111110101101100110;
    W_ir[12][59] = 26'b00000000000010000111111111;
    W_ir[12][60] = 26'b11111111111101010100000101;
    W_ir[12][61] = 26'b11111111111100110111101111;
    W_ir[12][62] = 26'b11111111111100110001111110;
    W_ir[12][63] = 26'b00000000000010000101110100;
    W_ir[13][0] = 26'b11111111111110001011100101;
    W_ir[13][1] = 26'b11111111111110011001011110;
    W_ir[13][2] = 26'b00000000000010111111010101;
    W_ir[13][3] = 26'b00000000000010010110010001;
    W_ir[13][4] = 26'b00000000000000010100010110;
    W_ir[13][5] = 26'b00000000000000111110001011;
    W_ir[13][6] = 26'b00000000000000110100100011;
    W_ir[13][7] = 26'b00000000000000100000111100;
    W_ir[13][8] = 26'b00000000000000101000000110;
    W_ir[13][9] = 26'b00000000000000100101000110;
    W_ir[13][10] = 26'b11111111111111100001110010;
    W_ir[13][11] = 26'b11111111111111111110110000;
    W_ir[13][12] = 26'b00000000000000101110101111;
    W_ir[13][13] = 26'b00000000000001110000000010;
    W_ir[13][14] = 26'b11111111111101010110100001;
    W_ir[13][15] = 26'b00000000000000100010000110;
    W_ir[13][16] = 26'b11111111111111111111010101;
    W_ir[13][17] = 26'b11111111111111111100011011;
    W_ir[13][18] = 26'b11111111111111110010001110;
    W_ir[13][19] = 26'b11111111111110101111110011;
    W_ir[13][20] = 26'b11111111111111110000001110;
    W_ir[13][21] = 26'b00000000000000101101101100;
    W_ir[13][22] = 26'b11111111111111000000000101;
    W_ir[13][23] = 26'b11111111111110100000000011;
    W_ir[13][24] = 26'b00000000000000000001010010;
    W_ir[13][25] = 26'b00000000000010111010010000;
    W_ir[13][26] = 26'b11111111111100110010100110;
    W_ir[13][27] = 26'b11111111111100111010100001;
    W_ir[13][28] = 26'b00000000000011010110011111;
    W_ir[13][29] = 26'b00000000000001000001001111;
    W_ir[13][30] = 26'b00000000000000001110100011;
    W_ir[13][31] = 26'b11111111111111111101101000;
    W_ir[13][32] = 26'b11111111111110000101001001;
    W_ir[13][33] = 26'b11111111111111110100011111;
    W_ir[13][34] = 26'b11111111111111101101010000;
    W_ir[13][35] = 26'b00000000000000001111000011;
    W_ir[13][36] = 26'b00000000000000111110110001;
    W_ir[13][37] = 26'b00000000000000100100010101;
    W_ir[13][38] = 26'b00000000000000110010010010;
    W_ir[13][39] = 26'b00000000000010000000010101;
    W_ir[13][40] = 26'b00000000000001001101001111;
    W_ir[13][41] = 26'b00000000000000000001100100;
    W_ir[13][42] = 26'b11111111111111110101010000;
    W_ir[13][43] = 26'b00000000000001000000110101;
    W_ir[13][44] = 26'b00000000000000011000101010;
    W_ir[13][45] = 26'b00000000000000110010011110;
    W_ir[13][46] = 26'b11111111111111110011101111;
    W_ir[13][47] = 26'b11111111111111011100010110;
    W_ir[13][48] = 26'b11111111111111011011011100;
    W_ir[13][49] = 26'b11111111111100101011101001;
    W_ir[13][50] = 26'b00000000000001111010010100;
    W_ir[13][51] = 26'b00000000000010101010101011;
    W_ir[13][52] = 26'b11111111111111001110000110;
    W_ir[13][53] = 26'b11111111111110011101101001;
    W_ir[13][54] = 26'b11111111111110100000000001;
    W_ir[13][55] = 26'b11111111111110010011011010;
    W_ir[13][56] = 26'b11111111111111000001100011;
    W_ir[13][57] = 26'b00000000000011001011011010;
    W_ir[13][58] = 26'b00000000000001110111010000;
    W_ir[13][59] = 26'b11111111111101111100010111;
    W_ir[13][60] = 26'b11111111111111011110011011;
    W_ir[13][61] = 26'b11111111111111001001101000;
    W_ir[13][62] = 26'b00000000000010101100001010;
    W_ir[13][63] = 26'b11111111111110011110111110;
    W_ir[14][0] = 26'b11111111111110100100011111;
    W_ir[14][1] = 26'b11111111111111000000011100;
    W_ir[14][2] = 26'b11111111111100100110000011;
    W_ir[14][3] = 26'b11111111111101111000110111;
    W_ir[14][4] = 26'b11111111111110110101100100;
    W_ir[14][5] = 26'b11111111111111011101011011;
    W_ir[14][6] = 26'b00000000000000010111100001;
    W_ir[14][7] = 26'b11111111111101011101100010;
    W_ir[14][8] = 26'b11111111111111010100001101;
    W_ir[14][9] = 26'b11111111111111010110000101;
    W_ir[14][10] = 26'b11111111111111010000011101;
    W_ir[14][11] = 26'b11111111111100010110011101;
    W_ir[14][12] = 26'b11111111111111011010111101;
    W_ir[14][13] = 26'b00000000000000110111100010;
    W_ir[14][14] = 26'b11111111111111010100001001;
    W_ir[14][15] = 26'b00000000000001010111110110;
    W_ir[14][16] = 26'b11111111111101011001111110;
    W_ir[14][17] = 26'b00000000000011100101011000;
    W_ir[14][18] = 26'b00000000000000001100000001;
    W_ir[14][19] = 26'b00000000000001001011110100;
    W_ir[14][20] = 26'b00000000000000110111101110;
    W_ir[14][21] = 26'b11111111111110110111111000;
    W_ir[14][22] = 26'b00000000000001110111110011;
    W_ir[14][23] = 26'b00000000000011010011111011;
    W_ir[14][24] = 26'b00000000000001101100000010;
    W_ir[14][25] = 26'b00000000000000100011010011;
    W_ir[14][26] = 26'b11111111111111110000001111;
    W_ir[14][27] = 26'b11111111111100101101101100;
    W_ir[14][28] = 26'b11111111111111000011110001;
    W_ir[14][29] = 26'b00000000000011110001010100;
    W_ir[14][30] = 26'b11111111111110011111111010;
    W_ir[14][31] = 26'b11111111111110100001000010;
    W_ir[14][32] = 26'b00000000000000001010110100;
    W_ir[14][33] = 26'b00000000000001011011110101;
    W_ir[14][34] = 26'b11111111111111010001001101;
    W_ir[14][35] = 26'b11111111111111001001110111;
    W_ir[14][36] = 26'b00000000000000001100001111;
    W_ir[14][37] = 26'b00000000000000101010010111;
    W_ir[14][38] = 26'b00000000000010000000001100;
    W_ir[14][39] = 26'b11111111111111111110101010;
    W_ir[14][40] = 26'b00000000000001110001111000;
    W_ir[14][41] = 26'b11111111111111001010101010;
    W_ir[14][42] = 26'b00000000000001110110010111;
    W_ir[14][43] = 26'b11111111111111110011001010;
    W_ir[14][44] = 26'b00000000000000101100111111;
    W_ir[14][45] = 26'b00000000000000111111010011;
    W_ir[14][46] = 26'b00000000000000110001111000;
    W_ir[14][47] = 26'b00000000000000011001111101;
    W_ir[14][48] = 26'b00000000000000110011100010;
    W_ir[14][49] = 26'b00000000000000101011010101;
    W_ir[14][50] = 26'b11111111111110000101111111;
    W_ir[14][51] = 26'b00000000000001010111000001;
    W_ir[14][52] = 26'b00000000000001010001111110;
    W_ir[14][53] = 26'b00000000000000111001000101;
    W_ir[14][54] = 26'b11111111111100100101001000;
    W_ir[14][55] = 26'b00000000000001001011001000;
    W_ir[14][56] = 26'b00000000000000110010000111;
    W_ir[14][57] = 26'b11111111111101011100111010;
    W_ir[14][58] = 26'b11111111111110000111101110;
    W_ir[14][59] = 26'b11111111111110010110010101;
    W_ir[14][60] = 26'b00000000000010011001011000;
    W_ir[14][61] = 26'b00000000000001000110001101;
    W_ir[14][62] = 26'b00000000000010011111001000;
    W_ir[14][63] = 26'b00000000000100011010010100;
    W_ir[15][0] = 26'b11111111111111110111011110;
    W_ir[15][1] = 26'b00000000000011111101100001;
    W_ir[15][2] = 26'b00000000000000000000100000;
    W_ir[15][3] = 26'b00000000000011001010011110;
    W_ir[15][4] = 26'b11111111111101001000000010;
    W_ir[15][5] = 26'b00000000000000101001011000;
    W_ir[15][6] = 26'b00000000000000011110100000;
    W_ir[15][7] = 26'b11111111111110110011010110;
    W_ir[15][8] = 26'b11111111111111100011001101;
    W_ir[15][9] = 26'b00000000000010100110101101;
    W_ir[15][10] = 26'b11111111111110001001101000;
    W_ir[15][11] = 26'b11111111111111101001111110;
    W_ir[15][12] = 26'b11111111111101111110100110;
    W_ir[15][13] = 26'b11111111111111010100101010;
    W_ir[15][14] = 26'b11111111111111000111101011;
    W_ir[15][15] = 26'b11111111111111100011000101;
    W_ir[15][16] = 26'b00000000000000001001101100;
    W_ir[15][17] = 26'b00000000000000101010110110;
    W_ir[15][18] = 26'b11111111111110100111000111;
    W_ir[15][19] = 26'b00000000000010000001111100;
    W_ir[15][20] = 26'b11111111111111001100000011;
    W_ir[15][21] = 26'b00000000000000110011010100;
    W_ir[15][22] = 26'b00000000000001010100011010;
    W_ir[15][23] = 26'b00000000000000110110011111;
    W_ir[15][24] = 26'b00000000000011010100010011;
    W_ir[15][25] = 26'b00000000000000101110100101;
    W_ir[15][26] = 26'b11111111111111100010000100;
    W_ir[15][27] = 26'b11111111111110110010101011;
    W_ir[15][28] = 26'b00000000000000101101010001;
    W_ir[15][29] = 26'b00000000000000100110001010;
    W_ir[15][30] = 26'b11111111111101111000000011;
    W_ir[15][31] = 26'b00000000000100001000111101;
    W_ir[15][32] = 26'b00000000000010000111110010;
    W_ir[15][33] = 26'b11111111111101100010011101;
    W_ir[15][34] = 26'b00000000000001000000001100;
    W_ir[15][35] = 26'b00000000000000100100110100;
    W_ir[15][36] = 26'b00000000000000101110111111;
    W_ir[15][37] = 26'b11111111111100011111101010;
    W_ir[15][38] = 26'b00000000000001100010010000;
    W_ir[15][39] = 26'b00000000000000001110011010;
    W_ir[15][40] = 26'b11111111111111111011010001;
    W_ir[15][41] = 26'b00000000000010010101010100;
    W_ir[15][42] = 26'b11111111111101011000110011;
    W_ir[15][43] = 26'b00000000000000011000001110;
    W_ir[15][44] = 26'b11111111111110100111111100;
    W_ir[15][45] = 26'b11111111111110111000100101;
    W_ir[15][46] = 26'b00000000000011000101110111;
    W_ir[15][47] = 26'b11111111111110100011100010;
    W_ir[15][48] = 26'b11111111111111001010000110;
    W_ir[15][49] = 26'b11111111111111011001100010;
    W_ir[15][50] = 26'b11111111111110001111111010;
    W_ir[15][51] = 26'b11111111111110100000010011;
    W_ir[15][52] = 26'b11111111111110010111100111;
    W_ir[15][53] = 26'b11111111111110001011010010;
    W_ir[15][54] = 26'b11111111111110111101100001;
    W_ir[15][55] = 26'b11111111111100011000001000;
    W_ir[15][56] = 26'b11111111111110010011001000;
    W_ir[15][57] = 26'b00000000000001111100111001;
    W_ir[15][58] = 26'b11111111111101110011100010;
    W_ir[15][59] = 26'b11111111111110011100011110;
    W_ir[15][60] = 26'b11111111111110011111111101;
    W_ir[15][61] = 26'b11111111111110101101010110;
    W_ir[15][62] = 26'b11111111111101000001000110;
    W_ir[15][63] = 26'b11111111111110110000001010;

    // Initialize W_iz weights
    W_iz[0][0] = 26'b11111111111111110010000001;
    W_iz[0][1] = 26'b11111111111111001101101000;
    W_iz[0][2] = 26'b11111111111111011010110110;
    W_iz[0][3] = 26'b11111111111110011100111100;
    W_iz[0][4] = 26'b00000000000000000101000010;
    W_iz[0][5] = 26'b00000000000001011100011001;
    W_iz[0][6] = 26'b11111111111110001101011110;
    W_iz[0][7] = 26'b11111111111101011101000111;
    W_iz[0][8] = 26'b11111111111100010100000010;
    W_iz[0][9] = 26'b11111111111110100101100101;
    W_iz[0][10] = 26'b11111111111100101110000101;
    W_iz[0][11] = 26'b11111111111110111100001000;
    W_iz[0][12] = 26'b11111111111111011010011000;
    W_iz[0][13] = 26'b00000000000001011100001011;
    W_iz[0][14] = 26'b00000000000000011001001001;
    W_iz[0][15] = 26'b11111111111111011010010100;
    W_iz[0][16] = 26'b11111111111110000011001110;
    W_iz[0][17] = 26'b11111111111110100010010111;
    W_iz[0][18] = 26'b11111111111110000110011001;
    W_iz[0][19] = 26'b11111111111101101010011010;
    W_iz[0][20] = 26'b11111111111111011100100001;
    W_iz[0][21] = 26'b00000000000001101011001101;
    W_iz[0][22] = 26'b00000000000100001110110100;
    W_iz[0][23] = 26'b00000000000010010101111110;
    W_iz[0][24] = 26'b11111111111100100000100101;
    W_iz[0][25] = 26'b11111111111101001011010011;
    W_iz[0][26] = 26'b00000000000000001110100110;
    W_iz[0][27] = 26'b11111111111100100000010111;
    W_iz[0][28] = 26'b00000000000010111110010001;
    W_iz[0][29] = 26'b11111111111111110110101110;
    W_iz[0][30] = 26'b00000000000010110101110111;
    W_iz[0][31] = 26'b11111111111110000100100100;
    W_iz[0][32] = 26'b11111111111100101111111111;
    W_iz[0][33] = 26'b11111111111101001010101110;
    W_iz[0][34] = 26'b11111111111110000110001111;
    W_iz[0][35] = 26'b11111111111101111011100100;
    W_iz[0][36] = 26'b11111111111100110110011101;
    W_iz[0][37] = 26'b11111111111101010101011100;
    W_iz[0][38] = 26'b11111111111110010010000110;
    W_iz[0][39] = 26'b00000000000001000100110110;
    W_iz[0][40] = 26'b00000000000000101111111011;
    W_iz[0][41] = 26'b11111111111110001100011101;
    W_iz[0][42] = 26'b11111111111111101111100111;
    W_iz[0][43] = 26'b11111111111110100111101001;
    W_iz[0][44] = 26'b11111111111100001000111000;
    W_iz[0][45] = 26'b11111111111111010101111011;
    W_iz[0][46] = 26'b11111111111111010101001001;
    W_iz[0][47] = 26'b11111111111111100001011001;
    W_iz[0][48] = 26'b00000000000000000000100110;
    W_iz[0][49] = 26'b11111111111111001001110110;
    W_iz[0][50] = 26'b00000000000010100111001011;
    W_iz[0][51] = 26'b11111111111110011011111001;
    W_iz[0][52] = 26'b00000000000011101010001011;
    W_iz[0][53] = 26'b00000000000001110001010000;
    W_iz[0][54] = 26'b00000000000011110110001001;
    W_iz[0][55] = 26'b00000000000011001101011001;
    W_iz[0][56] = 26'b00000000000001010000010001;
    W_iz[0][57] = 26'b11111111111100100001110111;
    W_iz[0][58] = 26'b00000000000010000011010101;
    W_iz[0][59] = 26'b00000000000110111011010000;
    W_iz[0][60] = 26'b00000000000101001011001100;
    W_iz[0][61] = 26'b00000000000101011101011000;
    W_iz[0][62] = 26'b00000000000110011100100010;
    W_iz[0][63] = 26'b00000000000101110000001010;
    W_iz[1][0] = 26'b00000000000000101010000111;
    W_iz[1][1] = 26'b00000000000000101101010100;
    W_iz[1][2] = 26'b00000000000000110101100001;
    W_iz[1][3] = 26'b11111111111111100000111000;
    W_iz[1][4] = 26'b11111111111111011101011111;
    W_iz[1][5] = 26'b11111111111101101100001000;
    W_iz[1][6] = 26'b00000000000011000111010101;
    W_iz[1][7] = 26'b11111111111100010101001110;
    W_iz[1][8] = 26'b11111111111101001001110110;
    W_iz[1][9] = 26'b11111111111110111101100010;
    W_iz[1][10] = 26'b11111111111111111010100011;
    W_iz[1][11] = 26'b11111111111111011010011110;
    W_iz[1][12] = 26'b11111111111101110000101010;
    W_iz[1][13] = 26'b11111111111111010110000100;
    W_iz[1][14] = 26'b11111111111110000011110001;
    W_iz[1][15] = 26'b11111111111101111111011000;
    W_iz[1][16] = 26'b00000000000010010011111000;
    W_iz[1][17] = 26'b11111111111101011111000101;
    W_iz[1][18] = 26'b00000000000000011110111101;
    W_iz[1][19] = 26'b11111111111100110111101110;
    W_iz[1][20] = 26'b11111111111111011000000100;
    W_iz[1][21] = 26'b00000000000000000101011010;
    W_iz[1][22] = 26'b00000000000001010010011110;
    W_iz[1][23] = 26'b00000000000000110011011011;
    W_iz[1][24] = 26'b11111111111111101011111101;
    W_iz[1][25] = 26'b11111111111110011110011011;
    W_iz[1][26] = 26'b11111111111111101100111100;
    W_iz[1][27] = 26'b00000000000001011100110100;
    W_iz[1][28] = 26'b00000000000000010100000001;
    W_iz[1][29] = 26'b11111111111110001010000010;
    W_iz[1][30] = 26'b11111111111111000100001110;
    W_iz[1][31] = 26'b11111111111100100010000100;
    W_iz[1][32] = 26'b11111111111111110001011001;
    W_iz[1][33] = 26'b11111111111100000000010010;
    W_iz[1][34] = 26'b11111111111110111111011000;
    W_iz[1][35] = 26'b00000000000001111100100101;
    W_iz[1][36] = 26'b11111111111110000001111110;
    W_iz[1][37] = 26'b11111111111101000100011101;
    W_iz[1][38] = 26'b11111111111011101001010010;
    W_iz[1][39] = 26'b00000000000010100011011110;
    W_iz[1][40] = 26'b11111111111110101110101000;
    W_iz[1][41] = 26'b11111111111111011111111101;
    W_iz[1][42] = 26'b00000000000000001101101101;
    W_iz[1][43] = 26'b11111111111110100110001100;
    W_iz[1][44] = 26'b00000000000000100001000111;
    W_iz[1][45] = 26'b11111111111110101001111111;
    W_iz[1][46] = 26'b11111111111111011011001100;
    W_iz[1][47] = 26'b00000000000001111010001001;
    W_iz[1][48] = 26'b00000000000000111100110111;
    W_iz[1][49] = 26'b00000000000000110010000100;
    W_iz[1][50] = 26'b00000000000000101010101010;
    W_iz[1][51] = 26'b00000000000000101100011101;
    W_iz[1][52] = 26'b11111111111110111011001001;
    W_iz[1][53] = 26'b11111111111110101101110111;
    W_iz[1][54] = 26'b00000000000000111010100100;
    W_iz[1][55] = 26'b00000000000000000000101010;
    W_iz[1][56] = 26'b00000000000000101100001011;
    W_iz[1][57] = 26'b11111111111101101111011110;
    W_iz[1][58] = 26'b11111111111101111001100110;
    W_iz[1][59] = 26'b11111111111110110110001001;
    W_iz[1][60] = 26'b00000000000011101110101010;
    W_iz[1][61] = 26'b00000000000010100001110101;
    W_iz[1][62] = 26'b11111111111110110000001100;
    W_iz[1][63] = 26'b00000000000010010000110110;
    W_iz[2][0] = 26'b00000000000010111010101011;
    W_iz[2][1] = 26'b11111111111111001110101111;
    W_iz[2][2] = 26'b00000000000100101011010000;
    W_iz[2][3] = 26'b11111111111110110011011101;
    W_iz[2][4] = 26'b00000000000010100111110011;
    W_iz[2][5] = 26'b00000000000000100111010110;
    W_iz[2][6] = 26'b11111111111100101100000111;
    W_iz[2][7] = 26'b00000000000100101100001101;
    W_iz[2][8] = 26'b00000000000101011000111110;
    W_iz[2][9] = 26'b00000000000011001010011111;
    W_iz[2][10] = 26'b00000000000011110110101100;
    W_iz[2][11] = 26'b11111111111111111010000001;
    W_iz[2][12] = 26'b00000000000000000011010001;
    W_iz[2][13] = 26'b00000000000001001010011001;
    W_iz[2][14] = 26'b11111111111110110111110100;
    W_iz[2][15] = 26'b11111111111100101110000111;
    W_iz[2][16] = 26'b11111111111110101001000111;
    W_iz[2][17] = 26'b00000000000010011101100000;
    W_iz[2][18] = 26'b11111111111111111010010001;
    W_iz[2][19] = 26'b11111111111111110100101100;
    W_iz[2][20] = 26'b11111111111111010001011000;
    W_iz[2][21] = 26'b11111111111101010101011001;
    W_iz[2][22] = 26'b00000000000100010110000011;
    W_iz[2][23] = 26'b11111111111111110101110100;
    W_iz[2][24] = 26'b11111111111101011101001010;
    W_iz[2][25] = 26'b00000000000001010000101100;
    W_iz[2][26] = 26'b11111111111101001111000100;
    W_iz[2][27] = 26'b11111111111101111000000010;
    W_iz[2][28] = 26'b00000000000011000011010010;
    W_iz[2][29] = 26'b00000000000010101000111011;
    W_iz[2][30] = 26'b11111111111101011000001111;
    W_iz[2][31] = 26'b00000000000010011001111111;
    W_iz[2][32] = 26'b00000000000000001101011100;
    W_iz[2][33] = 26'b00000000000001010000110010;
    W_iz[2][34] = 26'b00000000000011010110101011;
    W_iz[2][35] = 26'b00000000000100000001010000;
    W_iz[2][36] = 26'b11111111111111101100010001;
    W_iz[2][37] = 26'b00000000000000111110101110;
    W_iz[2][38] = 26'b11111111111100000101101011;
    W_iz[2][39] = 26'b11111111111111100110101101;
    W_iz[2][40] = 26'b00000000000001111111101000;
    W_iz[2][41] = 26'b11111111111110011101111111;
    W_iz[2][42] = 26'b00000000000100011011110001;
    W_iz[2][43] = 26'b00000000000001000011110111;
    W_iz[2][44] = 26'b00000000000010001000010001;
    W_iz[2][45] = 26'b11111111111110001010001111;
    W_iz[2][46] = 26'b11111111111100101110011001;
    W_iz[2][47] = 26'b00000000000011111111110000;
    W_iz[2][48] = 26'b11111111111101000000100001;
    W_iz[2][49] = 26'b11111111111110001001000011;
    W_iz[2][50] = 26'b00000000000010000000110001;
    W_iz[2][51] = 26'b11111111111111101101011001;
    W_iz[2][52] = 26'b00000000000010001000001110;
    W_iz[2][53] = 26'b11111111111001001011110000;
    W_iz[2][54] = 26'b11111111111111000101010110;
    W_iz[2][55] = 26'b00000000000000100110010010;
    W_iz[2][56] = 26'b11111111111101100101010011;
    W_iz[2][57] = 26'b11111111111110111000010100;
    W_iz[2][58] = 26'b11111111111101011100000011;
    W_iz[2][59] = 26'b11111111111101000001111101;
    W_iz[2][60] = 26'b11111111111111000101011100;
    W_iz[2][61] = 26'b11111111111001110111111000;
    W_iz[2][62] = 26'b11111111111000100111111011;
    W_iz[2][63] = 26'b11111111111000001011111000;
    W_iz[3][0] = 26'b11111111111010100101000101;
    W_iz[3][1] = 26'b11111111111010011000010011;
    W_iz[3][2] = 26'b00000000000001100011101001;
    W_iz[3][3] = 26'b11111111111111001100010011;
    W_iz[3][4] = 26'b00000000000011000110100010;
    W_iz[3][5] = 26'b00000000000100001111001011;
    W_iz[3][6] = 26'b11111111111100100101011000;
    W_iz[3][7] = 26'b00000000000000110100001001;
    W_iz[3][8] = 26'b11111111111101011101100010;
    W_iz[3][9] = 26'b11111111111001110010100100;
    W_iz[3][10] = 26'b11111111111101110111010100;
    W_iz[3][11] = 26'b00000000000010011110010110;
    W_iz[3][12] = 26'b00000000000010111111000111;
    W_iz[3][13] = 26'b11111111111101001101010100;
    W_iz[3][14] = 26'b00000000000011000001110011;
    W_iz[3][15] = 26'b11111111111111111111011001;
    W_iz[3][16] = 26'b00000000000000100111100110;
    W_iz[3][17] = 26'b11111111111110011111111101;
    W_iz[3][18] = 26'b00000000000000100110111101;
    W_iz[3][19] = 26'b00000000000011101011001011;
    W_iz[3][20] = 26'b11111111111110001111101111;
    W_iz[3][21] = 26'b11111111111110100010011001;
    W_iz[3][22] = 26'b00000000000011111101010101;
    W_iz[3][23] = 26'b11111111111110010100110100;
    W_iz[3][24] = 26'b00000000000011100100001111;
    W_iz[3][25] = 26'b00000000000001101110001100;
    W_iz[3][26] = 26'b00000000000010001010100010;
    W_iz[3][27] = 26'b11111111111111000111000010;
    W_iz[3][28] = 26'b00000000000010110101010000;
    W_iz[3][29] = 26'b00000000000100010000111110;
    W_iz[3][30] = 26'b00000000000010110010010001;
    W_iz[3][31] = 26'b00000000000001011111110010;
    W_iz[3][32] = 26'b11111111111101011100110010;
    W_iz[3][33] = 26'b11111111111110011101100110;
    W_iz[3][34] = 26'b11111111111010001110110110;
    W_iz[3][35] = 26'b11111111111100110100101001;
    W_iz[3][36] = 26'b00000000000011110010010010;
    W_iz[3][37] = 26'b00000000000000000010001101;
    W_iz[3][38] = 26'b00000000000011001100111110;
    W_iz[3][39] = 26'b11111111111011101111101011;
    W_iz[3][40] = 26'b11111111111111110110110001;
    W_iz[3][41] = 26'b11111111111011110111111001;
    W_iz[3][42] = 26'b11111111111011100110100100;
    W_iz[3][43] = 26'b11111111111011011100000110;
    W_iz[3][44] = 26'b11111111111101101010000110;
    W_iz[3][45] = 26'b00000000000000100110011110;
    W_iz[3][46] = 26'b00000000001000110000011011;
    W_iz[3][47] = 26'b11111111111101101001010101;
    W_iz[3][48] = 26'b11111111111111100110110011;
    W_iz[3][49] = 26'b11111111111101011001110101;
    W_iz[3][50] = 26'b11111111111100001001111100;
    W_iz[3][51] = 26'b00000000000101110110001100;
    W_iz[3][52] = 26'b11111111111011101001101110;
    W_iz[3][53] = 26'b00000000000001011000101100;
    W_iz[3][54] = 26'b00000000000100011011111011;
    W_iz[3][55] = 26'b00000000000000101101000100;
    W_iz[3][56] = 26'b00000000001001000101101110;
    W_iz[3][57] = 26'b00000000000001001001101001;
    W_iz[3][58] = 26'b00000000001001010001010100;
    W_iz[3][59] = 26'b00000000000001011110100011;
    W_iz[3][60] = 26'b11111111111100001001110101;
    W_iz[3][61] = 26'b00000000000100011100000101;
    W_iz[3][62] = 26'b00000000000110000001100100;
    W_iz[3][63] = 26'b11111111111100001001111000;
    W_iz[4][0] = 26'b11111111111110001110100011;
    W_iz[4][1] = 26'b00000000000000111101111100;
    W_iz[4][2] = 26'b11111111111111001100010000;
    W_iz[4][3] = 26'b00000000000010001101110100;
    W_iz[4][4] = 26'b11111111111111011001001100;
    W_iz[4][5] = 26'b11111111111110111001011101;
    W_iz[4][6] = 26'b11111111111100100000000111;
    W_iz[4][7] = 26'b11111111111110000110100000;
    W_iz[4][8] = 26'b11111111111110111010010110;
    W_iz[4][9] = 26'b00000000000010010110010110;
    W_iz[4][10] = 26'b00000000000001000101101010;
    W_iz[4][11] = 26'b00000000000011011101110110;
    W_iz[4][12] = 26'b11111111111111000100010000;
    W_iz[4][13] = 26'b00000000000001110011000110;
    W_iz[4][14] = 26'b00000000000001110001111010;
    W_iz[4][15] = 26'b00000000000000110000101010;
    W_iz[4][16] = 26'b11111111111111010110011010;
    W_iz[4][17] = 26'b00000000000010101110101111;
    W_iz[4][18] = 26'b00000000000011111111000010;
    W_iz[4][19] = 26'b00000000000010001101110110;
    W_iz[4][20] = 26'b11111111111111100110101111;
    W_iz[4][21] = 26'b00000000000000101110110100;
    W_iz[4][22] = 26'b00000000000010110001101110;
    W_iz[4][23] = 26'b00000000000000101000000010;
    W_iz[4][24] = 26'b00000000000000001111011101;
    W_iz[4][25] = 26'b11111111111111010100011000;
    W_iz[4][26] = 26'b11111111111100010011001011;
    W_iz[4][27] = 26'b00000000000000110101111110;
    W_iz[4][28] = 26'b00000000000001111100110010;
    W_iz[4][29] = 26'b00000000000000001010111011;
    W_iz[4][30] = 26'b00000000000010011110011010;
    W_iz[4][31] = 26'b00000000000010000111010100;
    W_iz[4][32] = 26'b11111111111111011011000101;
    W_iz[4][33] = 26'b11111111111101101111100111;
    W_iz[4][34] = 26'b11111111111100111000000100;
    W_iz[4][35] = 26'b11111111111110011101101011;
    W_iz[4][36] = 26'b11111111111110010001001110;
    W_iz[4][37] = 26'b11111111111010110100100100;
    W_iz[4][38] = 26'b00000000000000111000111111;
    W_iz[4][39] = 26'b11111111111111101110010000;
    W_iz[4][40] = 26'b11111111111111010010111011;
    W_iz[4][41] = 26'b00000000000011011010111011;
    W_iz[4][42] = 26'b11111111111101010111001111;
    W_iz[4][43] = 26'b00000000000010001010111000;
    W_iz[4][44] = 26'b00000000000000000001011110;
    W_iz[4][45] = 26'b11111111111110000001111011;
    W_iz[4][46] = 26'b11111111111101101010011100;
    W_iz[4][47] = 26'b00000000000010101011101110;
    W_iz[4][48] = 26'b00000000000001000110010011;
    W_iz[4][49] = 26'b00000000000100101110100101;
    W_iz[4][50] = 26'b11111111111111111111000110;
    W_iz[4][51] = 26'b00000000000000111101101001;
    W_iz[4][52] = 26'b11111111111110110101000101;
    W_iz[4][53] = 26'b11111111111101000111100011;
    W_iz[4][54] = 26'b11111111111100101100100011;
    W_iz[4][55] = 26'b11111111111110010110111011;
    W_iz[4][56] = 26'b00000000000011101100000001;
    W_iz[4][57] = 26'b11111111111110110100110100;
    W_iz[4][58] = 26'b00000000000011110011100011;
    W_iz[4][59] = 26'b11111111111111001000010111;
    W_iz[4][60] = 26'b11111111111011101000101001;
    W_iz[4][61] = 26'b11111111111001000111111100;
    W_iz[4][62] = 26'b11111111111000000011011110;
    W_iz[4][63] = 26'b00000000000001101111011100;
    W_iz[5][0] = 26'b00000000000011001011001011;
    W_iz[5][1] = 26'b00000000000001000110010100;
    W_iz[5][2] = 26'b00000000000000101101100111;
    W_iz[5][3] = 26'b00000000000000000011001001;
    W_iz[5][4] = 26'b00000000000000011110111010;
    W_iz[5][5] = 26'b00000000000010011010001010;
    W_iz[5][6] = 26'b11111111111100110100011101;
    W_iz[5][7] = 26'b11111111111101011010001101;
    W_iz[5][8] = 26'b00000000000000000100111010;
    W_iz[5][9] = 26'b00000000000100000010001010;
    W_iz[5][10] = 26'b00000000000010000100111110;
    W_iz[5][11] = 26'b11111111111011110010010001;
    W_iz[5][12] = 26'b11111111111101011011110011;
    W_iz[5][13] = 26'b00000000000010101110000101;
    W_iz[5][14] = 26'b11111111111111001010110010;
    W_iz[5][15] = 26'b00000000000011001101001011;
    W_iz[5][16] = 26'b11111111111100001110001001;
    W_iz[5][17] = 26'b00000000000001110110101110;
    W_iz[5][18] = 26'b00000000000100100010000101;
    W_iz[5][19] = 26'b11111111111101010000110110;
    W_iz[5][20] = 26'b11111111111101100110010111;
    W_iz[5][21] = 26'b11111111111100010000011111;
    W_iz[5][22] = 26'b00000000000010001101100001;
    W_iz[5][23] = 26'b00000000000101001111010111;
    W_iz[5][24] = 26'b00000000000001111011111000;
    W_iz[5][25] = 26'b11111111111110000101010011;
    W_iz[5][26] = 26'b11111111111110011000000111;
    W_iz[5][27] = 26'b11111111111101111010111001;
    W_iz[5][28] = 26'b11111111111110101001110010;
    W_iz[5][29] = 26'b11111111111100110110000111;
    W_iz[5][30] = 26'b11111111111111000111010000;
    W_iz[5][31] = 26'b11111111111100110011011011;
    W_iz[5][32] = 26'b00000000000010011100111000;
    W_iz[5][33] = 26'b11111111111110111110010111;
    W_iz[5][34] = 26'b11111111111101111110001100;
    W_iz[5][35] = 26'b00000000000010100101101001;
    W_iz[5][36] = 26'b11111111111011011011011111;
    W_iz[5][37] = 26'b00000000000000101001110101;
    W_iz[5][38] = 26'b11111111111111111000110010;
    W_iz[5][39] = 26'b11111111111101111110000000;
    W_iz[5][40] = 26'b00000000000010110110011011;
    W_iz[5][41] = 26'b00000000000001011011111100;
    W_iz[5][42] = 26'b00000000000011101111110000;
    W_iz[5][43] = 26'b00000000000011001101101111;
    W_iz[5][44] = 26'b00000000000000001100010111;
    W_iz[5][45] = 26'b00000000000011101010100001;
    W_iz[5][46] = 26'b00000000000001000001010000;
    W_iz[5][47] = 26'b11111111111111001001011100;
    W_iz[5][48] = 26'b11111111111101000101000100;
    W_iz[5][49] = 26'b11111111111111011010111110;
    W_iz[5][50] = 26'b11111111111110010100101101;
    W_iz[5][51] = 26'b00000000000001110100100011;
    W_iz[5][52] = 26'b00000000000010101110000101;
    W_iz[5][53] = 26'b00000000000001100010000010;
    W_iz[5][54] = 26'b11111111111100001011111111;
    W_iz[5][55] = 26'b00000000000100110010111100;
    W_iz[5][56] = 26'b00000000000010011010001101;
    W_iz[5][57] = 26'b11111111111111000010100101;
    W_iz[5][58] = 26'b11111111111111101101111110;
    W_iz[5][59] = 26'b00000000000011011111000010;
    W_iz[5][60] = 26'b11111111111011101110001111;
    W_iz[5][61] = 26'b11111111111111110011001001;
    W_iz[5][62] = 26'b11111111111110010010000011;
    W_iz[5][63] = 26'b11111111111110100000000111;
    W_iz[6][0] = 26'b00000000000001011011101000;
    W_iz[6][1] = 26'b00000000000001111110011000;
    W_iz[6][2] = 26'b11111111111111010000100000;
    W_iz[6][3] = 26'b00000000000000110001101001;
    W_iz[6][4] = 26'b00000000000011001101001101;
    W_iz[6][5] = 26'b00000000000001011001000111;
    W_iz[6][6] = 26'b11111111111011011001111100;
    W_iz[6][7] = 26'b00000000000001011100100011;
    W_iz[6][8] = 26'b11111111111010000011000101;
    W_iz[6][9] = 26'b11111111111111001100110111;
    W_iz[6][10] = 26'b11111111111111111011010111;
    W_iz[6][11] = 26'b11111111111110001111010101;
    W_iz[6][12] = 26'b11111111111100100001110101;
    W_iz[6][13] = 26'b00000000000001100100110110;
    W_iz[6][14] = 26'b11111111111111110010000101;
    W_iz[6][15] = 26'b11111111111010100110100111;
    W_iz[6][16] = 26'b00000000000010000100010011;
    W_iz[6][17] = 26'b00000000000010010100011110;
    W_iz[6][18] = 26'b11111111111010000100000010;
    W_iz[6][19] = 26'b11111111111011110011011000;
    W_iz[6][20] = 26'b00000000000011010011010011;
    W_iz[6][21] = 26'b11111111111100110111101000;
    W_iz[6][22] = 26'b00000000000001010110100000;
    W_iz[6][23] = 26'b11111111111101000001100010;
    W_iz[6][24] = 26'b00000000000001100101010001;
    W_iz[6][25] = 26'b11111111111101010011011100;
    W_iz[6][26] = 26'b00000000000100101011101000;
    W_iz[6][27] = 26'b11111111111111001111100111;
    W_iz[6][28] = 26'b00000000000010110011111101;
    W_iz[6][29] = 26'b00000000000100011011101011;
    W_iz[6][30] = 26'b11111111111111011000010001;
    W_iz[6][31] = 26'b00000000000000000001001010;
    W_iz[6][32] = 26'b00000000000101011011111011;
    W_iz[6][33] = 26'b11111111111011111001110010;
    W_iz[6][34] = 26'b11111111111100001011101101;
    W_iz[6][35] = 26'b11111111111110001011000000;
    W_iz[6][36] = 26'b00000000000101000010111001;
    W_iz[6][37] = 26'b00000000000100001011011101;
    W_iz[6][38] = 26'b11111111111101011010000111;
    W_iz[6][39] = 26'b11111111111010101110101100;
    W_iz[6][40] = 26'b00000000000010001101110001;
    W_iz[6][41] = 26'b11111111111111101100110101;
    W_iz[6][42] = 26'b11111111111100001110011010;
    W_iz[6][43] = 26'b00000000000000101100100000;
    W_iz[6][44] = 26'b11111111111110101101101100;
    W_iz[6][45] = 26'b00000000000010011001111110;
    W_iz[6][46] = 26'b11111111111111000111001111;
    W_iz[6][47] = 26'b11111111111111000110001101;
    W_iz[6][48] = 26'b11111111111110011111100100;
    W_iz[6][49] = 26'b11111111111111111100010100;
    W_iz[6][50] = 26'b11111111111100001110000101;
    W_iz[6][51] = 26'b11111111111110011010011110;
    W_iz[6][52] = 26'b11111111111011111011111011;
    W_iz[6][53] = 26'b00000000000011011010011011;
    W_iz[6][54] = 26'b11111111111111011111111010;
    W_iz[6][55] = 26'b11111111111110001110001000;
    W_iz[6][56] = 26'b11111111111110010010100100;
    W_iz[6][57] = 26'b00000000000011100110100100;
    W_iz[6][58] = 26'b00000000000011110111001010;
    W_iz[6][59] = 26'b00000000000100110110011110;
    W_iz[6][60] = 26'b00000000000111100101011010;
    W_iz[6][61] = 26'b00000000000101000101101000;
    W_iz[6][62] = 26'b00000000001000101110110110;
    W_iz[6][63] = 26'b00000000000110011110011110;
    W_iz[7][0] = 26'b11111111111010011000111100;
    W_iz[7][1] = 26'b00000000000100000101101011;
    W_iz[7][2] = 26'b00000000000000010011010110;
    W_iz[7][3] = 26'b00000000000100011011110010;
    W_iz[7][4] = 26'b11111111111010111001000111;
    W_iz[7][5] = 26'b00000000000001000110101110;
    W_iz[7][6] = 26'b11111111111011100001000110;
    W_iz[7][7] = 26'b00000000000010011110011111;
    W_iz[7][8] = 26'b11111111111001000110111001;
    W_iz[7][9] = 26'b11111111111010011000001111;
    W_iz[7][10] = 26'b00000000000100101000010100;
    W_iz[7][11] = 26'b11111111111010011000101011;
    W_iz[7][12] = 26'b11111111111010100011011100;
    W_iz[7][13] = 26'b00000000000010010100100010;
    W_iz[7][14] = 26'b00000000000001111110100100;
    W_iz[7][15] = 26'b00000000000001111111010000;
    W_iz[7][16] = 26'b00000000000101010100010001;
    W_iz[7][17] = 26'b11111111111110111000110110;
    W_iz[7][18] = 26'b11111111111111111110100111;
    W_iz[7][19] = 26'b00000000000110010110001100;
    W_iz[7][20] = 26'b11111111111111000001111100;
    W_iz[7][21] = 26'b11111111111100001110001100;
    W_iz[7][22] = 26'b11111111111110100101010101;
    W_iz[7][23] = 26'b11111111111110001011010100;
    W_iz[7][24] = 26'b11111111111011000010110001;
    W_iz[7][25] = 26'b11111111111111000101100011;
    W_iz[7][26] = 26'b11111111111011111101100111;
    W_iz[7][27] = 26'b11111111111010111111100110;
    W_iz[7][28] = 26'b00000000000110100110110010;
    W_iz[7][29] = 26'b00000000000010001101101001;
    W_iz[7][30] = 26'b00000000000000011001101000;
    W_iz[7][31] = 26'b00000000000011101010100011;
    W_iz[7][32] = 26'b00000000000010001001111100;
    W_iz[7][33] = 26'b11111111111111000000100100;
    W_iz[7][34] = 26'b00000000000011100100111101;
    W_iz[7][35] = 26'b00000000000001110011010000;
    W_iz[7][36] = 26'b11111111111011101111001000;
    W_iz[7][37] = 26'b11111111111010110110110111;
    W_iz[7][38] = 26'b00000000000010001001011100;
    W_iz[7][39] = 26'b11111111111111110100110110;
    W_iz[7][40] = 26'b11111111111010000010010101;
    W_iz[7][41] = 26'b11111111111010110011000110;
    W_iz[7][42] = 26'b00000000000100000101011001;
    W_iz[7][43] = 26'b00000000000000010111101011;
    W_iz[7][44] = 26'b00000000000001011000101011;
    W_iz[7][45] = 26'b00000000000110001110001011;
    W_iz[7][46] = 26'b11111111111111011011111101;
    W_iz[7][47] = 26'b00000000000101000000101000;
    W_iz[7][48] = 26'b00000000000000100110000000;
    W_iz[7][49] = 26'b11111111111111011010110100;
    W_iz[7][50] = 26'b11111111111101010011011110;
    W_iz[7][51] = 26'b00000000000010110011000101;
    W_iz[7][52] = 26'b11111111111110110000100011;
    W_iz[7][53] = 26'b11111111111010111100011101;
    W_iz[7][54] = 26'b00000000000110001000111110;
    W_iz[7][55] = 26'b00000000000000111100101001;
    W_iz[7][56] = 26'b11111111111101000110100001;
    W_iz[7][57] = 26'b00000000000010110101111011;
    W_iz[7][58] = 26'b11111111111101100111011111;
    W_iz[7][59] = 26'b00000000000101100010100110;
    W_iz[7][60] = 26'b00000000000101011101001011;
    W_iz[7][61] = 26'b00000000000001010011010000;
    W_iz[7][62] = 26'b00000000000000011100100101;
    W_iz[7][63] = 26'b00000000000100101111011110;
    W_iz[8][0] = 26'b00000000000001010010011110;
    W_iz[8][1] = 26'b00000000000010011100011000;
    W_iz[8][2] = 26'b00000000000001110111001110;
    W_iz[8][3] = 26'b00000000000010001100110010;
    W_iz[8][4] = 26'b11111111111110110100110100;
    W_iz[8][5] = 26'b11111111111101010101000001;
    W_iz[8][6] = 26'b00000000000001110011010001;
    W_iz[8][7] = 26'b00000000000000111101101110;
    W_iz[8][8] = 26'b11111111111100100000101110;
    W_iz[8][9] = 26'b00000000000000010110011000;
    W_iz[8][10] = 26'b00000000000011111010111111;
    W_iz[8][11] = 26'b11111111111111111110101100;
    W_iz[8][12] = 26'b00000000000010011111111001;
    W_iz[8][13] = 26'b00000000000000101100000000;
    W_iz[8][14] = 26'b00000000000000100111011101;
    W_iz[8][15] = 26'b00000000000010111001011010;
    W_iz[8][16] = 26'b11111111111111100000000101;
    W_iz[8][17] = 26'b00000000000011011100110111;
    W_iz[8][18] = 26'b11111111111111100011001001;
    W_iz[8][19] = 26'b00000000000010010001001011;
    W_iz[8][20] = 26'b11111111111111100001111100;
    W_iz[8][21] = 26'b00000000000010000111001000;
    W_iz[8][22] = 26'b00000000000001100001111111;
    W_iz[8][23] = 26'b00000000000001100011100000;
    W_iz[8][24] = 26'b11111111111101011110111110;
    W_iz[8][25] = 26'b00000000000001111000001100;
    W_iz[8][26] = 26'b00000000000010001011100110;
    W_iz[8][27] = 26'b00000000000001011011010101;
    W_iz[8][28] = 26'b00000000000011100010100110;
    W_iz[8][29] = 26'b11111111111100101100001011;
    W_iz[8][30] = 26'b11111111111110110101100001;
    W_iz[8][31] = 26'b00000000000001100111000001;
    W_iz[8][32] = 26'b00000000000000110001101110;
    W_iz[8][33] = 26'b00000000000001111010001100;
    W_iz[8][34] = 26'b00000000000001111010011110;
    W_iz[8][35] = 26'b00000000000000011010111101;
    W_iz[8][36] = 26'b00000000000011111110101101;
    W_iz[8][37] = 26'b00000000000001010001000000;
    W_iz[8][38] = 26'b11111111111110111011001110;
    W_iz[8][39] = 26'b00000000000000111101100110;
    W_iz[8][40] = 26'b00000000000010010101101000;
    W_iz[8][41] = 26'b11111111111101000000111011;
    W_iz[8][42] = 26'b00000000000000111100111010;
    W_iz[8][43] = 26'b11111111111110100001001011;
    W_iz[8][44] = 26'b11111111111111111001001101;
    W_iz[8][45] = 26'b11111111111101110010100010;
    W_iz[8][46] = 26'b11111111111100111001111111;
    W_iz[8][47] = 26'b00000000000011011110110000;
    W_iz[8][48] = 26'b11111111111111000101001111;
    W_iz[8][49] = 26'b11111111111110011100100001;
    W_iz[8][50] = 26'b11111111111111100110010101;
    W_iz[8][51] = 26'b00000000000000000001001000;
    W_iz[8][52] = 26'b11111111111100011011000001;
    W_iz[8][53] = 26'b11111111111110101001001010;
    W_iz[8][54] = 26'b00000000000001000011001101;
    W_iz[8][55] = 26'b11111111111110011111000000;
    W_iz[8][56] = 26'b00000000000010011001010000;
    W_iz[8][57] = 26'b11111111111110010101100110;
    W_iz[8][58] = 26'b11111111111110101101100110;
    W_iz[8][59] = 26'b00000000000010000111111111;
    W_iz[8][60] = 26'b11111111111101010100000101;
    W_iz[8][61] = 26'b11111111111100110111101111;
    W_iz[8][62] = 26'b11111111111100110001111110;
    W_iz[8][63] = 26'b00000000000010000101110100;
    W_iz[9][0] = 26'b11111111111110001011100101;
    W_iz[9][1] = 26'b11111111111110011001011110;
    W_iz[9][2] = 26'b00000000000010111111010101;
    W_iz[9][3] = 26'b00000000000010010110010001;
    W_iz[9][4] = 26'b00000000000000010100010110;
    W_iz[9][5] = 26'b00000000000000111110001011;
    W_iz[9][6] = 26'b00000000000000110100100011;
    W_iz[9][7] = 26'b00000000000000100000111100;
    W_iz[9][8] = 26'b00000000000000101000000110;
    W_iz[9][9] = 26'b00000000000000100101000110;
    W_iz[9][10] = 26'b11111111111111100001110010;
    W_iz[9][11] = 26'b11111111111111111110110000;
    W_iz[9][12] = 26'b00000000000000101110101111;
    W_iz[9][13] = 26'b00000000000001110000000010;
    W_iz[9][14] = 26'b11111111111101010110100001;
    W_iz[9][15] = 26'b00000000000000100010000110;
    W_iz[9][16] = 26'b11111111111111111111010101;
    W_iz[9][17] = 26'b11111111111111111100011011;
    W_iz[9][18] = 26'b11111111111111110010001110;
    W_iz[9][19] = 26'b11111111111110101111110011;
    W_iz[9][20] = 26'b11111111111111110000001110;
    W_iz[9][21] = 26'b00000000000000101101101100;
    W_iz[9][22] = 26'b11111111111111000000000101;
    W_iz[9][23] = 26'b11111111111110100000000011;
    W_iz[9][24] = 26'b00000000000000000001010010;
    W_iz[9][25] = 26'b00000000000010111010010000;
    W_iz[9][26] = 26'b11111111111100110010100110;
    W_iz[9][27] = 26'b11111111111100111010100001;
    W_iz[9][28] = 26'b00000000000011010110011111;
    W_iz[9][29] = 26'b00000000000001000001001111;
    W_iz[9][30] = 26'b00000000000000001110100011;
    W_iz[9][31] = 26'b11111111111111111101101000;
    W_iz[9][32] = 26'b11111111111110000101001001;
    W_iz[9][33] = 26'b11111111111111110100011111;
    W_iz[9][34] = 26'b11111111111111101101010000;
    W_iz[9][35] = 26'b00000000000000001111000011;
    W_iz[9][36] = 26'b00000000000000111110110001;
    W_iz[9][37] = 26'b00000000000000100100010101;
    W_iz[9][38] = 26'b00000000000000110010010010;
    W_iz[9][39] = 26'b00000000000010000000010101;
    W_iz[9][40] = 26'b00000000000001001101001111;
    W_iz[9][41] = 26'b00000000000000000001100100;
    W_iz[9][42] = 26'b11111111111111110101010000;
    W_iz[9][43] = 26'b00000000000001000000110101;
    W_iz[9][44] = 26'b00000000000000011000101010;
    W_iz[9][45] = 26'b00000000000000110010011110;
    W_iz[9][46] = 26'b11111111111111110011101111;
    W_iz[9][47] = 26'b11111111111111011100010110;
    W_iz[9][48] = 26'b11111111111111011011011100;
    W_iz[9][49] = 26'b11111111111100101011101001;
    W_iz[9][50] = 26'b00000000000001111010010100;
    W_iz[9][51] = 26'b00000000000010101010101011;
    W_iz[9][52] = 26'b11111111111111001110000110;
    W_iz[9][53] = 26'b11111111111110011101101001;
    W_iz[9][54] = 26'b11111111111110100000000001;
    W_iz[9][55] = 26'b11111111111110010011011010;
    W_iz[9][56] = 26'b11111111111111000001100011;
    W_iz[9][57] = 26'b00000000000011001011011010;
    W_iz[9][58] = 26'b00000000000001110111010000;
    W_iz[9][59] = 26'b11111111111101111100010111;
    W_iz[9][60] = 26'b11111111111111011110011011;
    W_iz[9][61] = 26'b11111111111111001001101000;
    W_iz[9][62] = 26'b00000000000010101100001010;
    W_iz[9][63] = 26'b11111111111110011110111110;
    W_iz[10][0] = 26'b11111111111110100100011111;
    W_iz[10][1] = 26'b11111111111111000000011100;
    W_iz[10][2] = 26'b11111111111100100110000011;
    W_iz[10][3] = 26'b11111111111101111000110111;
    W_iz[10][4] = 26'b11111111111110110101100100;
    W_iz[10][5] = 26'b11111111111111011101011011;
    W_iz[10][6] = 26'b00000000000000010111100001;
    W_iz[10][7] = 26'b11111111111101011101100010;
    W_iz[10][8] = 26'b11111111111111010100001101;
    W_iz[10][9] = 26'b11111111111111010110000101;
    W_iz[10][10] = 26'b11111111111111010000011101;
    W_iz[10][11] = 26'b11111111111100010110011101;
    W_iz[10][12] = 26'b11111111111111011010111101;
    W_iz[10][13] = 26'b00000000000000110111100010;
    W_iz[10][14] = 26'b11111111111111010100001001;
    W_iz[10][15] = 26'b00000000000001010111110110;
    W_iz[10][16] = 26'b11111111111101011001111110;
    W_iz[10][17] = 26'b00000000000011100101011000;
    W_iz[10][18] = 26'b00000000000000001100000001;
    W_iz[10][19] = 26'b00000000000001001011110100;
    W_iz[10][20] = 26'b00000000000000110111101110;
    W_iz[10][21] = 26'b11111111111110110111111000;
    W_iz[10][22] = 26'b00000000000001110111110011;
    W_iz[10][23] = 26'b00000000000011010011111011;
    W_iz[10][24] = 26'b00000000000001101100000010;
    W_iz[10][25] = 26'b00000000000000100011010011;
    W_iz[10][26] = 26'b11111111111111110000001111;
    W_iz[10][27] = 26'b11111111111100101101101100;
    W_iz[10][28] = 26'b11111111111111000011110001;
    W_iz[10][29] = 26'b00000000000011110001010100;
    W_iz[10][30] = 26'b11111111111110011111111010;
    W_iz[10][31] = 26'b11111111111110100001000010;
    W_iz[10][32] = 26'b00000000000000001010110100;
    W_iz[10][33] = 26'b00000000000001011011110101;
    W_iz[10][34] = 26'b11111111111111010001001101;
    W_iz[10][35] = 26'b11111111111111001001110111;
    W_iz[10][36] = 26'b00000000000000001100001111;
    W_iz[10][37] = 26'b00000000000000101010010111;
    W_iz[10][38] = 26'b00000000000010000000001100;
    W_iz[10][39] = 26'b11111111111111111110101010;
    W_iz[10][40] = 26'b00000000000001110001111000;
    W_iz[10][41] = 26'b11111111111111001010101010;
    W_iz[10][42] = 26'b00000000000001110110010111;
    W_iz[10][43] = 26'b11111111111111110011001010;
    W_iz[10][44] = 26'b00000000000000101100111111;
    W_iz[10][45] = 26'b00000000000000111111010011;
    W_iz[10][46] = 26'b00000000000000110001111000;
    W_iz[10][47] = 26'b00000000000000011001111101;
    W_iz[10][48] = 26'b00000000000000110011100010;
    W_iz[10][49] = 26'b00000000000000101011010101;
    W_iz[10][50] = 26'b11111111111110000101111111;
    W_iz[10][51] = 26'b00000000000001010111000001;
    W_iz[10][52] = 26'b00000000000001010001111110;
    W_iz[10][53] = 26'b00000000000000111001000101;
    W_iz[10][54] = 26'b11111111111100100101001000;
    W_iz[10][55] = 26'b00000000000001001011001000;
    W_iz[10][56] = 26'b00000000000000110010000111;
    W_iz[10][57] = 26'b11111111111101011100111010;
    W_iz[10][58] = 26'b11111111111110000111101110;
    W_iz[10][59] = 26'b11111111111110010110010101;
    W_iz[10][60] = 26'b00000000000010011001011000;
    W_iz[10][61] = 26'b00000000000001000110001101;
    W_iz[10][62] = 26'b00000000000010011111001000;
    W_iz[10][63] = 26'b00000000000100011010010100;
    W_iz[11][0] = 26'b11111111111111110111011110;
    W_iz[11][1] = 26'b00000000000011111101100001;
    W_iz[11][2] = 26'b00000000000000000000100000;
    W_iz[11][3] = 26'b00000000000011001010011110;
    W_iz[11][4] = 26'b11111111111101001000000010;
    W_iz[11][5] = 26'b00000000000000101001011000;
    W_iz[11][6] = 26'b00000000000000011110100000;
    W_iz[11][7] = 26'b11111111111110110011010110;
    W_iz[11][8] = 26'b11111111111111100011001101;
    W_iz[11][9] = 26'b00000000000010100110101101;
    W_iz[11][10] = 26'b11111111111110001001101000;
    W_iz[11][11] = 26'b11111111111111101001111110;
    W_iz[11][12] = 26'b11111111111101111110100110;
    W_iz[11][13] = 26'b11111111111111010100101010;
    W_iz[11][14] = 26'b11111111111111000111101011;
    W_iz[11][15] = 26'b11111111111111100011000101;
    W_iz[11][16] = 26'b00000000000000001001101100;
    W_iz[11][17] = 26'b00000000000000101010110110;
    W_iz[11][18] = 26'b11111111111110100111000111;
    W_iz[11][19] = 26'b00000000000010000001111100;
    W_iz[11][20] = 26'b11111111111111001100000011;
    W_iz[11][21] = 26'b00000000000000110011010100;
    W_iz[11][22] = 26'b00000000000001010100011010;
    W_iz[11][23] = 26'b00000000000000110110011111;
    W_iz[11][24] = 26'b00000000000011010100010011;
    W_iz[11][25] = 26'b00000000000000101110100101;
    W_iz[11][26] = 26'b11111111111111100010000100;
    W_iz[11][27] = 26'b11111111111110110010101011;
    W_iz[11][28] = 26'b00000000000000101101010001;
    W_iz[11][29] = 26'b00000000000000100110001010;
    W_iz[11][30] = 26'b11111111111101111000000011;
    W_iz[11][31] = 26'b00000000000100001000111101;
    W_iz[11][32] = 26'b00000000000010000111110010;
    W_iz[11][33] = 26'b11111111111101100010011101;
    W_iz[11][34] = 26'b00000000000001000000001100;
    W_iz[11][35] = 26'b00000000000000100100110100;
    W_iz[11][36] = 26'b00000000000000101110111111;
    W_iz[11][37] = 26'b11111111111100011111101010;
    W_iz[11][38] = 26'b00000000000001100010010000;
    W_iz[11][39] = 26'b00000000000000001110011010;
    W_iz[11][40] = 26'b11111111111111111011010001;
    W_iz[11][41] = 26'b00000000000010010101010100;
    W_iz[11][42] = 26'b11111111111101011000110011;
    W_iz[11][43] = 26'b00000000000000011000001110;
    W_iz[11][44] = 26'b11111111111110100111111100;
    W_iz[11][45] = 26'b11111111111110111000100101;
    W_iz[11][46] = 26'b00000000000011000101110111;
    W_iz[11][47] = 26'b11111111111110100011100010;
    W_iz[11][48] = 26'b11111111111111001010000110;
    W_iz[11][49] = 26'b11111111111111011001100010;
    W_iz[11][50] = 26'b11111111111110001111111010;
    W_iz[11][51] = 26'b11111111111110100000010011;
    W_iz[11][52] = 26'b11111111111110010111100111;
    W_iz[11][53] = 26'b11111111111110001011010010;
    W_iz[11][54] = 26'b11111111111110111101100001;
    W_iz[11][55] = 26'b11111111111100011000001000;
    W_iz[11][56] = 26'b11111111111110010011001000;
    W_iz[11][57] = 26'b00000000000001111100111001;
    W_iz[11][58] = 26'b11111111111101110011100010;
    W_iz[11][59] = 26'b11111111111110011100011110;
    W_iz[11][60] = 26'b11111111111110011111111101;
    W_iz[11][61] = 26'b11111111111110101101010110;
    W_iz[11][62] = 26'b11111111111101000001000110;
    W_iz[11][63] = 26'b11111111111110110000001010;
    W_iz[12][0] = 26'b11111111111111110010000001;
    W_iz[12][1] = 26'b11111111111111001101101000;
    W_iz[12][2] = 26'b11111111111111011010110110;
    W_iz[12][3] = 26'b11111111111110011100111100;
    W_iz[12][4] = 26'b00000000000000000101000010;
    W_iz[12][5] = 26'b00000000000001011100011001;
    W_iz[12][6] = 26'b11111111111110001101011110;
    W_iz[12][7] = 26'b11111111111101011101000111;
    W_iz[12][8] = 26'b11111111111100010100000010;
    W_iz[12][9] = 26'b11111111111110100101100101;
    W_iz[12][10] = 26'b11111111111100101110000101;
    W_iz[12][11] = 26'b11111111111110111100001000;
    W_iz[12][12] = 26'b11111111111111011010011000;
    W_iz[12][13] = 26'b00000000000001011100001011;
    W_iz[12][14] = 26'b00000000000000011001001001;
    W_iz[12][15] = 26'b11111111111111011010010100;
    W_iz[12][16] = 26'b11111111111110000011001110;
    W_iz[12][17] = 26'b11111111111110100010010111;
    W_iz[12][18] = 26'b11111111111110000110011001;
    W_iz[12][19] = 26'b11111111111101101010011010;
    W_iz[12][20] = 26'b11111111111111011100100001;
    W_iz[12][21] = 26'b00000000000001101011001101;
    W_iz[12][22] = 26'b00000000000100001110110100;
    W_iz[12][23] = 26'b00000000000010010101111110;
    W_iz[12][24] = 26'b11111111111100100000100101;
    W_iz[12][25] = 26'b11111111111101001011010011;
    W_iz[12][26] = 26'b00000000000000001110100110;
    W_iz[12][27] = 26'b11111111111100100000010111;
    W_iz[12][28] = 26'b00000000000010111110010001;
    W_iz[12][29] = 26'b11111111111111110110101110;
    W_iz[12][30] = 26'b00000000000010110101110111;
    W_iz[12][31] = 26'b11111111111110000100100100;
    W_iz[12][32] = 26'b11111111111100101111111111;
    W_iz[12][33] = 26'b11111111111101001010101110;
    W_iz[12][34] = 26'b11111111111110000110001111;
    W_iz[12][35] = 26'b11111111111101111011100100;
    W_iz[12][36] = 26'b11111111111100110110011101;
    W_iz[12][37] = 26'b11111111111101010101011100;
    W_iz[12][38] = 26'b11111111111110010010000110;
    W_iz[12][39] = 26'b00000000000001000100110110;
    W_iz[12][40] = 26'b00000000000000101111111011;
    W_iz[12][41] = 26'b11111111111110001100011101;
    W_iz[12][42] = 26'b11111111111111101111100111;
    W_iz[12][43] = 26'b11111111111110100111101001;
    W_iz[12][44] = 26'b11111111111100001000111000;
    W_iz[12][45] = 26'b11111111111111010101111011;
    W_iz[12][46] = 26'b11111111111111010101001001;
    W_iz[12][47] = 26'b11111111111111100001011001;
    W_iz[12][48] = 26'b00000000000000000000100110;
    W_iz[12][49] = 26'b11111111111111001001110110;
    W_iz[12][50] = 26'b00000000000010100111001011;
    W_iz[12][51] = 26'b11111111111110011011111001;
    W_iz[12][52] = 26'b00000000000011101010001011;
    W_iz[12][53] = 26'b00000000000001110001010000;
    W_iz[12][54] = 26'b00000000000011110110001001;
    W_iz[12][55] = 26'b00000000000011001101011001;
    W_iz[12][56] = 26'b00000000000001010000010001;
    W_iz[12][57] = 26'b11111111111100100001110111;
    W_iz[12][58] = 26'b00000000000010000011010101;
    W_iz[12][59] = 26'b00000000000110111011010000;
    W_iz[12][60] = 26'b00000000000101001011001100;
    W_iz[12][61] = 26'b00000000000101011101011000;
    W_iz[12][62] = 26'b00000000000110011100100010;
    W_iz[12][63] = 26'b00000000000101110000001010;
    W_iz[13][0] = 26'b00000000000000101010000111;
    W_iz[13][1] = 26'b00000000000000101101010100;
    W_iz[13][2] = 26'b00000000000000110101100001;
    W_iz[13][3] = 26'b11111111111111100000111000;
    W_iz[13][4] = 26'b11111111111111011101011111;
    W_iz[13][5] = 26'b11111111111101101100001000;
    W_iz[13][6] = 26'b00000000000011000111010101;
    W_iz[13][7] = 26'b11111111111100010101001110;
    W_iz[13][8] = 26'b11111111111101001001110110;
    W_iz[13][9] = 26'b11111111111110111101100010;
    W_iz[13][10] = 26'b11111111111111111010100011;
    W_iz[13][11] = 26'b11111111111111011010011110;
    W_iz[13][12] = 26'b11111111111101110000101010;
    W_iz[13][13] = 26'b11111111111111010110000100;
    W_iz[13][14] = 26'b11111111111110000011110001;
    W_iz[13][15] = 26'b11111111111101111111011000;
    W_iz[13][16] = 26'b00000000000010010011111000;
    W_iz[13][17] = 26'b11111111111101011111000101;
    W_iz[13][18] = 26'b00000000000000011110111101;
    W_iz[13][19] = 26'b11111111111100110111101110;
    W_iz[13][20] = 26'b11111111111111011000000100;
    W_iz[13][21] = 26'b00000000000000000101011010;
    W_iz[13][22] = 26'b00000000000001010010011110;
    W_iz[13][23] = 26'b00000000000000110011011011;
    W_iz[13][24] = 26'b11111111111111101011111101;
    W_iz[13][25] = 26'b11111111111110011110011011;
    W_iz[13][26] = 26'b11111111111111101100111100;
    W_iz[13][27] = 26'b00000000000001011100110100;
    W_iz[13][28] = 26'b00000000000000010100000001;
    W_iz[13][29] = 26'b11111111111110001010000010;
    W_iz[13][30] = 26'b11111111111111000100001110;
    W_iz[13][31] = 26'b11111111111100100010000100;
    W_iz[13][32] = 26'b11111111111111110001011001;
    W_iz[13][33] = 26'b11111111111100000000010010;
    W_iz[13][34] = 26'b11111111111110111111011000;
    W_iz[13][35] = 26'b00000000000001111100100101;
    W_iz[13][36] = 26'b11111111111110000001111110;
    W_iz[13][37] = 26'b11111111111101000100011101;
    W_iz[13][38] = 26'b11111111111011101001010010;
    W_iz[13][39] = 26'b00000000000010100011011110;
    W_iz[13][40] = 26'b11111111111110101110101000;
    W_iz[13][41] = 26'b11111111111111011111111101;
    W_iz[13][42] = 26'b00000000000000001101101101;
    W_iz[13][43] = 26'b11111111111110100110001100;
    W_iz[13][44] = 26'b00000000000000100001000111;
    W_iz[13][45] = 26'b11111111111110101001111111;
    W_iz[13][46] = 26'b11111111111111011011001100;
    W_iz[13][47] = 26'b00000000000001111010001001;
    W_iz[13][48] = 26'b00000000000000111100110111;
    W_iz[13][49] = 26'b00000000000000110010000100;
    W_iz[13][50] = 26'b00000000000000101010101010;
    W_iz[13][51] = 26'b00000000000000101100011101;
    W_iz[13][52] = 26'b11111111111110111011001001;
    W_iz[13][53] = 26'b11111111111110101101110111;
    W_iz[13][54] = 26'b00000000000000111010100100;
    W_iz[13][55] = 26'b00000000000000000000101010;
    W_iz[13][56] = 26'b00000000000000101100001011;
    W_iz[13][57] = 26'b11111111111101101111011110;
    W_iz[13][58] = 26'b11111111111101111001100110;
    W_iz[13][59] = 26'b11111111111110110110001001;
    W_iz[13][60] = 26'b00000000000011101110101010;
    W_iz[13][61] = 26'b00000000000010100001110101;
    W_iz[13][62] = 26'b11111111111110110000001100;
    W_iz[13][63] = 26'b00000000000010010000110110;
    W_iz[14][0] = 26'b00000000000010111010101011;
    W_iz[14][1] = 26'b11111111111111001110101111;
    W_iz[14][2] = 26'b00000000000100101011010000;
    W_iz[14][3] = 26'b11111111111110110011011101;
    W_iz[14][4] = 26'b00000000000010100111110011;
    W_iz[14][5] = 26'b00000000000000100111010110;
    W_iz[14][6] = 26'b11111111111100101100000111;
    W_iz[14][7] = 26'b00000000000100101100001101;
    W_iz[14][8] = 26'b00000000000101011000111110;
    W_iz[14][9] = 26'b00000000000011001010011111;
    W_iz[14][10] = 26'b00000000000011110110101100;
    W_iz[14][11] = 26'b11111111111111111010000001;
    W_iz[14][12] = 26'b00000000000000000011010001;
    W_iz[14][13] = 26'b00000000000001001010011001;
    W_iz[14][14] = 26'b11111111111110110111110100;
    W_iz[14][15] = 26'b11111111111100101110000111;
    W_iz[14][16] = 26'b11111111111110101001000111;
    W_iz[14][17] = 26'b00000000000010011101100000;
    W_iz[14][18] = 26'b11111111111111111010010001;
    W_iz[14][19] = 26'b11111111111111110100101100;
    W_iz[14][20] = 26'b11111111111111010001011000;
    W_iz[14][21] = 26'b11111111111101010101011001;
    W_iz[14][22] = 26'b00000000000100010110000011;
    W_iz[14][23] = 26'b11111111111111110101110100;
    W_iz[14][24] = 26'b11111111111101011101001010;
    W_iz[14][25] = 26'b00000000000001010000101100;
    W_iz[14][26] = 26'b11111111111101001111000100;
    W_iz[14][27] = 26'b11111111111101111000000010;
    W_iz[14][28] = 26'b00000000000011000011010010;
    W_iz[14][29] = 26'b00000000000010101000111011;
    W_iz[14][30] = 26'b11111111111101011000001111;
    W_iz[14][31] = 26'b00000000000010011001111111;
    W_iz[14][32] = 26'b00000000000000001101011100;
    W_iz[14][33] = 26'b00000000000001010000110010;
    W_iz[14][34] = 26'b00000000000011010110101011;
    W_iz[14][35] = 26'b00000000000100000001010000;
    W_iz[14][36] = 26'b11111111111111101100010001;
    W_iz[14][37] = 26'b00000000000000111110101110;
    W_iz[14][38] = 26'b11111111111100000101101011;
    W_iz[14][39] = 26'b11111111111111100110101101;
    W_iz[14][40] = 26'b00000000000001111111101000;
    W_iz[14][41] = 26'b11111111111110011101111111;
    W_iz[14][42] = 26'b00000000000100011011110001;
    W_iz[14][43] = 26'b00000000000001000011110111;
    W_iz[14][44] = 26'b00000000000010001000010001;
    W_iz[14][45] = 26'b11111111111110001010001111;
    W_iz[14][46] = 26'b11111111111100101110011001;
    W_iz[14][47] = 26'b00000000000011111111110000;
    W_iz[14][48] = 26'b11111111111101000000100001;
    W_iz[14][49] = 26'b11111111111110001001000011;
    W_iz[14][50] = 26'b00000000000010000000110001;
    W_iz[14][51] = 26'b11111111111111101101011001;
    W_iz[14][52] = 26'b00000000000010001000001110;
    W_iz[14][53] = 26'b11111111111001001011110000;
    W_iz[14][54] = 26'b11111111111111000101010110;
    W_iz[14][55] = 26'b00000000000000100110010010;
    W_iz[14][56] = 26'b11111111111101100101010011;
    W_iz[14][57] = 26'b11111111111110111000010100;
    W_iz[14][58] = 26'b11111111111101011100000011;
    W_iz[14][59] = 26'b11111111111101000001111101;
    W_iz[14][60] = 26'b11111111111111000101011100;
    W_iz[14][61] = 26'b11111111111001110111111000;
    W_iz[14][62] = 26'b11111111111000100111111011;
    W_iz[14][63] = 26'b11111111111000001011111000;
    W_iz[15][0] = 26'b11111111111010100101000101;
    W_iz[15][1] = 26'b11111111111010011000010011;
    W_iz[15][2] = 26'b00000000000001100011101001;
    W_iz[15][3] = 26'b11111111111111001100010011;
    W_iz[15][4] = 26'b00000000000011000110100010;
    W_iz[15][5] = 26'b00000000000100001111001011;
    W_iz[15][6] = 26'b11111111111100100101011000;
    W_iz[15][7] = 26'b00000000000000110100001001;
    W_iz[15][8] = 26'b11111111111101011101100010;
    W_iz[15][9] = 26'b11111111111001110010100100;
    W_iz[15][10] = 26'b11111111111101110111010100;
    W_iz[15][11] = 26'b00000000000010011110010110;
    W_iz[15][12] = 26'b00000000000010111111000111;
    W_iz[15][13] = 26'b11111111111101001101010100;
    W_iz[15][14] = 26'b00000000000011000001110011;
    W_iz[15][15] = 26'b11111111111111111111011001;
    W_iz[15][16] = 26'b00000000000000100111100110;
    W_iz[15][17] = 26'b11111111111110011111111101;
    W_iz[15][18] = 26'b00000000000000100110111101;
    W_iz[15][19] = 26'b00000000000011101011001011;
    W_iz[15][20] = 26'b11111111111110001111101111;
    W_iz[15][21] = 26'b11111111111110100010011001;
    W_iz[15][22] = 26'b00000000000011111101010101;
    W_iz[15][23] = 26'b11111111111110010100110100;
    W_iz[15][24] = 26'b00000000000011100100001111;
    W_iz[15][25] = 26'b00000000000001101110001100;
    W_iz[15][26] = 26'b00000000000010001010100010;
    W_iz[15][27] = 26'b11111111111111000111000010;
    W_iz[15][28] = 26'b00000000000010110101010000;
    W_iz[15][29] = 26'b00000000000100010000111110;
    W_iz[15][30] = 26'b00000000000010110010010001;
    W_iz[15][31] = 26'b00000000000001011111110010;
    W_iz[15][32] = 26'b11111111111101011100110010;
    W_iz[15][33] = 26'b11111111111110011101100110;
    W_iz[15][34] = 26'b11111111111010001110110110;
    W_iz[15][35] = 26'b11111111111100110100101001;
    W_iz[15][36] = 26'b00000000000011110010010010;
    W_iz[15][37] = 26'b00000000000000000010001101;
    W_iz[15][38] = 26'b00000000000011001100111110;
    W_iz[15][39] = 26'b11111111111011101111101011;
    W_iz[15][40] = 26'b11111111111111110110110001;
    W_iz[15][41] = 26'b11111111111011110111111001;
    W_iz[15][42] = 26'b11111111111011100110100100;
    W_iz[15][43] = 26'b11111111111011011100000110;
    W_iz[15][44] = 26'b11111111111101101010000110;
    W_iz[15][45] = 26'b00000000000000100110011110;
    W_iz[15][46] = 26'b00000000001000110000011011;
    W_iz[15][47] = 26'b11111111111101101001010101;
    W_iz[15][48] = 26'b11111111111111100110110011;
    W_iz[15][49] = 26'b11111111111101011001110101;
    W_iz[15][50] = 26'b11111111111100001001111100;
    W_iz[15][51] = 26'b00000000000101110110001100;
    W_iz[15][52] = 26'b11111111111011101001101110;
    W_iz[15][53] = 26'b00000000000001011000101100;
    W_iz[15][54] = 26'b00000000000100011011111011;
    W_iz[15][55] = 26'b00000000000000101101000100;
    W_iz[15][56] = 26'b00000000001001000101101110;
    W_iz[15][57] = 26'b00000000000001001001101001;
    W_iz[15][58] = 26'b00000000001001010001010100;
    W_iz[15][59] = 26'b00000000000001011110100011;
    W_iz[15][60] = 26'b11111111111100001001110101;
    W_iz[15][61] = 26'b00000000000100011100000101;
    W_iz[15][62] = 26'b00000000000110000001100100;
    W_iz[15][63] = 26'b11111111111100001001111000;

    // Initialize W_in weights
    W_in[0][0] = 26'b11111111111110001110100011;
    W_in[0][1] = 26'b00000000000000111101111100;
    W_in[0][2] = 26'b11111111111111001100010000;
    W_in[0][3] = 26'b00000000000010001101110100;
    W_in[0][4] = 26'b11111111111111011001001100;
    W_in[0][5] = 26'b11111111111110111001011101;
    W_in[0][6] = 26'b11111111111100100000000111;
    W_in[0][7] = 26'b11111111111110000110100000;
    W_in[0][8] = 26'b11111111111110111010010110;
    W_in[0][9] = 26'b00000000000010010110010110;
    W_in[0][10] = 26'b00000000000001000101101010;
    W_in[0][11] = 26'b00000000000011011101110110;
    W_in[0][12] = 26'b11111111111111000100010000;
    W_in[0][13] = 26'b00000000000001110011000110;
    W_in[0][14] = 26'b00000000000001110001111010;
    W_in[0][15] = 26'b00000000000000110000101010;
    W_in[0][16] = 26'b11111111111111010110011010;
    W_in[0][17] = 26'b00000000000010101110101111;
    W_in[0][18] = 26'b00000000000011111111000010;
    W_in[0][19] = 26'b00000000000010001101110110;
    W_in[0][20] = 26'b11111111111111100110101111;
    W_in[0][21] = 26'b00000000000000101110110100;
    W_in[0][22] = 26'b00000000000010110001101110;
    W_in[0][23] = 26'b00000000000000101000000010;
    W_in[0][24] = 26'b00000000000000001111011101;
    W_in[0][25] = 26'b11111111111111010100011000;
    W_in[0][26] = 26'b11111111111100010011001011;
    W_in[0][27] = 26'b00000000000000110101111110;
    W_in[0][28] = 26'b00000000000001111100110010;
    W_in[0][29] = 26'b00000000000000001010111011;
    W_in[0][30] = 26'b00000000000010011110011010;
    W_in[0][31] = 26'b00000000000010000111010100;
    W_in[0][32] = 26'b11111111111111011011000101;
    W_in[0][33] = 26'b11111111111101101111100111;
    W_in[0][34] = 26'b11111111111100111000000100;
    W_in[0][35] = 26'b11111111111110011101101011;
    W_in[0][36] = 26'b11111111111110010001001110;
    W_in[0][37] = 26'b11111111111010110100100100;
    W_in[0][38] = 26'b00000000000000111000111111;
    W_in[0][39] = 26'b11111111111111101110010000;
    W_in[0][40] = 26'b11111111111111010010111011;
    W_in[0][41] = 26'b00000000000011011010111011;
    W_in[0][42] = 26'b11111111111101010111001111;
    W_in[0][43] = 26'b00000000000010001010111000;
    W_in[0][44] = 26'b00000000000000000001011110;
    W_in[0][45] = 26'b11111111111110000001111011;
    W_in[0][46] = 26'b11111111111101101010011100;
    W_in[0][47] = 26'b00000000000010101011101110;
    W_in[0][48] = 26'b00000000000001000110010011;
    W_in[0][49] = 26'b00000000000100101110100101;
    W_in[0][50] = 26'b11111111111111111111000110;
    W_in[0][51] = 26'b00000000000000111101101001;
    W_in[0][52] = 26'b11111111111110110101000101;
    W_in[0][53] = 26'b11111111111101000111100011;
    W_in[0][54] = 26'b11111111111100101100100011;
    W_in[0][55] = 26'b11111111111110010110111011;
    W_in[0][56] = 26'b00000000000011101100000001;
    W_in[0][57] = 26'b11111111111110110100110100;
    W_in[0][58] = 26'b00000000000011110011100011;
    W_in[0][59] = 26'b11111111111111001000010111;
    W_in[0][60] = 26'b11111111111011101000101001;
    W_in[0][61] = 26'b11111111111001000111111100;
    W_in[0][62] = 26'b11111111111000000011011110;
    W_in[0][63] = 26'b00000000000001101111011100;
    W_in[1][0] = 26'b00000000000011001011001011;
    W_in[1][1] = 26'b00000000000001000110010100;
    W_in[1][2] = 26'b00000000000000101101100111;
    W_in[1][3] = 26'b00000000000000000011001001;
    W_in[1][4] = 26'b00000000000000011110111010;
    W_in[1][5] = 26'b00000000000010011010001010;
    W_in[1][6] = 26'b11111111111100110100011101;
    W_in[1][7] = 26'b11111111111101011010001101;
    W_in[1][8] = 26'b00000000000000000100111010;
    W_in[1][9] = 26'b00000000000100000010001010;
    W_in[1][10] = 26'b00000000000010000100111110;
    W_in[1][11] = 26'b11111111111011110010010001;
    W_in[1][12] = 26'b11111111111101011011110011;
    W_in[1][13] = 26'b00000000000010101110000101;
    W_in[1][14] = 26'b11111111111111001010110010;
    W_in[1][15] = 26'b00000000000011001101001011;
    W_in[1][16] = 26'b11111111111100001110001001;
    W_in[1][17] = 26'b00000000000001110110101110;
    W_in[1][18] = 26'b00000000000100100010000101;
    W_in[1][19] = 26'b11111111111101010000110110;
    W_in[1][20] = 26'b11111111111101100110010111;
    W_in[1][21] = 26'b11111111111100010000011111;
    W_in[1][22] = 26'b00000000000010001101100001;
    W_in[1][23] = 26'b00000000000101001111010111;
    W_in[1][24] = 26'b00000000000001111011111000;
    W_in[1][25] = 26'b11111111111110000101010011;
    W_in[1][26] = 26'b11111111111110011000000111;
    W_in[1][27] = 26'b11111111111101111010111001;
    W_in[1][28] = 26'b11111111111110101001110010;
    W_in[1][29] = 26'b11111111111100110110000111;
    W_in[1][30] = 26'b11111111111111000111010000;
    W_in[1][31] = 26'b11111111111100110011011011;
    W_in[1][32] = 26'b00000000000010011100111000;
    W_in[1][33] = 26'b11111111111110111110010111;
    W_in[1][34] = 26'b11111111111101111110001100;
    W_in[1][35] = 26'b00000000000010100101101001;
    W_in[1][36] = 26'b11111111111011011011011111;
    W_in[1][37] = 26'b00000000000000101001110101;
    W_in[1][38] = 26'b11111111111111111000110010;
    W_in[1][39] = 26'b11111111111101111110000000;
    W_in[1][40] = 26'b00000000000010110110011011;
    W_in[1][41] = 26'b00000000000001011011111100;
    W_in[1][42] = 26'b00000000000011101111110000;
    W_in[1][43] = 26'b00000000000011001101101111;
    W_in[1][44] = 26'b00000000000000001100010111;
    W_in[1][45] = 26'b00000000000011101010100001;
    W_in[1][46] = 26'b00000000000001000001010000;
    W_in[1][47] = 26'b11111111111111001001011100;
    W_in[1][48] = 26'b11111111111101000101000100;
    W_in[1][49] = 26'b11111111111111011010111110;
    W_in[1][50] = 26'b11111111111110010100101101;
    W_in[1][51] = 26'b00000000000001110100100011;
    W_in[1][52] = 26'b00000000000010101110000101;
    W_in[1][53] = 26'b00000000000001100010000010;
    W_in[1][54] = 26'b11111111111100001011111111;
    W_in[1][55] = 26'b00000000000100110010111100;
    W_in[1][56] = 26'b00000000000010011010001101;
    W_in[1][57] = 26'b11111111111111000010100101;
    W_in[1][58] = 26'b11111111111111101101111110;
    W_in[1][59] = 26'b00000000000011011111000010;
    W_in[1][60] = 26'b11111111111011101110001111;
    W_in[1][61] = 26'b11111111111111110011001001;
    W_in[1][62] = 26'b11111111111110010010000011;
    W_in[1][63] = 26'b11111111111110100000000111;
    W_in[2][0] = 26'b00000000000001011011101000;
    W_in[2][1] = 26'b00000000000001111110011000;
    W_in[2][2] = 26'b11111111111111010000100000;
    W_in[2][3] = 26'b00000000000000110001101001;
    W_in[2][4] = 26'b00000000000011001101001101;
    W_in[2][5] = 26'b00000000000001011001000111;
    W_in[2][6] = 26'b11111111111011011001111100;
    W_in[2][7] = 26'b00000000000001011100100011;
    W_in[2][8] = 26'b11111111111010000011000101;
    W_in[2][9] = 26'b11111111111111001100110111;
    W_in[2][10] = 26'b11111111111111111011010111;
    W_in[2][11] = 26'b11111111111110001111010101;
    W_in[2][12] = 26'b11111111111100100001110101;
    W_in[2][13] = 26'b00000000000001100100110110;
    W_in[2][14] = 26'b11111111111111110010000101;
    W_in[2][15] = 26'b11111111111010100110100111;
    W_in[2][16] = 26'b00000000000010000100010011;
    W_in[2][17] = 26'b00000000000010010100011110;
    W_in[2][18] = 26'b11111111111010000100000010;
    W_in[2][19] = 26'b11111111111011110011011000;
    W_in[2][20] = 26'b00000000000011010011010011;
    W_in[2][21] = 26'b11111111111100110111101000;
    W_in[2][22] = 26'b00000000000001010110100000;
    W_in[2][23] = 26'b11111111111101000001100010;
    W_in[2][24] = 26'b00000000000001100101010001;
    W_in[2][25] = 26'b11111111111101010011011100;
    W_in[2][26] = 26'b00000000000100101011101000;
    W_in[2][27] = 26'b11111111111111001111100111;
    W_in[2][28] = 26'b00000000000010110011111101;
    W_in[2][29] = 26'b00000000000100011011101011;
    W_in[2][30] = 26'b11111111111111011000010001;
    W_in[2][31] = 26'b00000000000000000001001010;
    W_in[2][32] = 26'b00000000000101011011111011;
    W_in[2][33] = 26'b11111111111011111001110010;
    W_in[2][34] = 26'b11111111111100001011101101;
    W_in[2][35] = 26'b11111111111110001011000000;
    W_in[2][36] = 26'b00000000000101000010111001;
    W_in[2][37] = 26'b00000000000100001011011101;
    W_in[2][38] = 26'b11111111111101011010000111;
    W_in[2][39] = 26'b11111111111010101110101100;
    W_in[2][40] = 26'b00000000000010001101110001;
    W_in[2][41] = 26'b11111111111111101100110101;
    W_in[2][42] = 26'b11111111111100001110011010;
    W_in[2][43] = 26'b00000000000000101100100000;
    W_in[2][44] = 26'b11111111111110101101101100;
    W_in[2][45] = 26'b00000000000010011001111110;
    W_in[2][46] = 26'b11111111111111000111001111;
    W_in[2][47] = 26'b11111111111111000110001101;
    W_in[2][48] = 26'b11111111111110011111100100;
    W_in[2][49] = 26'b11111111111111111100010100;
    W_in[2][50] = 26'b11111111111100001110000101;
    W_in[2][51] = 26'b11111111111110011010011110;
    W_in[2][52] = 26'b11111111111011111011111011;
    W_in[2][53] = 26'b00000000000011011010011011;
    W_in[2][54] = 26'b11111111111111011111111010;
    W_in[2][55] = 26'b11111111111110001110001000;
    W_in[2][56] = 26'b11111111111110010010100100;
    W_in[2][57] = 26'b00000000000011100110100100;
    W_in[2][58] = 26'b00000000000011110111001010;
    W_in[2][59] = 26'b00000000000100110110011110;
    W_in[2][60] = 26'b00000000000111100101011010;
    W_in[2][61] = 26'b00000000000101000101101000;
    W_in[2][62] = 26'b00000000001000101110110110;
    W_in[2][63] = 26'b00000000000110011110011110;
    W_in[3][0] = 26'b11111111111010011000111100;
    W_in[3][1] = 26'b00000000000100000101101011;
    W_in[3][2] = 26'b00000000000000010011010110;
    W_in[3][3] = 26'b00000000000100011011110010;
    W_in[3][4] = 26'b11111111111010111001000111;
    W_in[3][5] = 26'b00000000000001000110101110;
    W_in[3][6] = 26'b11111111111011100001000110;
    W_in[3][7] = 26'b00000000000010011110011111;
    W_in[3][8] = 26'b11111111111001000110111001;
    W_in[3][9] = 26'b11111111111010011000001111;
    W_in[3][10] = 26'b00000000000100101000010100;
    W_in[3][11] = 26'b11111111111010011000101011;
    W_in[3][12] = 26'b11111111111010100011011100;
    W_in[3][13] = 26'b00000000000010010100100010;
    W_in[3][14] = 26'b00000000000001111110100100;
    W_in[3][15] = 26'b00000000000001111111010000;
    W_in[3][16] = 26'b00000000000101010100010001;
    W_in[3][17] = 26'b11111111111110111000110110;
    W_in[3][18] = 26'b11111111111111111110100111;
    W_in[3][19] = 26'b00000000000110010110001100;
    W_in[3][20] = 26'b11111111111111000001111100;
    W_in[3][21] = 26'b11111111111100001110001100;
    W_in[3][22] = 26'b11111111111110100101010101;
    W_in[3][23] = 26'b11111111111110001011010100;
    W_in[3][24] = 26'b11111111111011000010110001;
    W_in[3][25] = 26'b11111111111111000101100011;
    W_in[3][26] = 26'b11111111111011111101100111;
    W_in[3][27] = 26'b11111111111010111111100110;
    W_in[3][28] = 26'b00000000000110100110110010;
    W_in[3][29] = 26'b00000000000010001101101001;
    W_in[3][30] = 26'b00000000000000011001101000;
    W_in[3][31] = 26'b00000000000011101010100011;
    W_in[3][32] = 26'b00000000000010001001111100;
    W_in[3][33] = 26'b11111111111111000000100100;
    W_in[3][34] = 26'b00000000000011100100111101;
    W_in[3][35] = 26'b00000000000001110011010000;
    W_in[3][36] = 26'b11111111111011101111001000;
    W_in[3][37] = 26'b11111111111010110110110111;
    W_in[3][38] = 26'b00000000000010001001011100;
    W_in[3][39] = 26'b11111111111111110100110110;
    W_in[3][40] = 26'b11111111111010000010010101;
    W_in[3][41] = 26'b11111111111010110011000110;
    W_in[3][42] = 26'b00000000000100000101011001;
    W_in[3][43] = 26'b00000000000000010111101011;
    W_in[3][44] = 26'b00000000000001011000101011;
    W_in[3][45] = 26'b00000000000110001110001011;
    W_in[3][46] = 26'b11111111111111011011111101;
    W_in[3][47] = 26'b00000000000101000000101000;
    W_in[3][48] = 26'b00000000000000100110000000;
    W_in[3][49] = 26'b11111111111111011010110100;
    W_in[3][50] = 26'b11111111111101010011011110;
    W_in[3][51] = 26'b00000000000010110011000101;
    W_in[3][52] = 26'b11111111111110110000100011;
    W_in[3][53] = 26'b11111111111010111100011101;
    W_in[3][54] = 26'b00000000000110001000111110;
    W_in[3][55] = 26'b00000000000000111100101001;
    W_in[3][56] = 26'b11111111111101000110100001;
    W_in[3][57] = 26'b00000000000010110101111011;
    W_in[3][58] = 26'b11111111111101100111011111;
    W_in[3][59] = 26'b00000000000101100010100110;
    W_in[3][60] = 26'b00000000000101011101001011;
    W_in[3][61] = 26'b00000000000001010011010000;
    W_in[3][62] = 26'b00000000000000011100100101;
    W_in[3][63] = 26'b00000000000100101111011110;
    W_in[4][0] = 26'b00000000000001010010011110;
    W_in[4][1] = 26'b00000000000010011100011000;
    W_in[4][2] = 26'b00000000000001110111001110;
    W_in[4][3] = 26'b00000000000010001100110010;
    W_in[4][4] = 26'b11111111111110110100110100;
    W_in[4][5] = 26'b11111111111101010101000001;
    W_in[4][6] = 26'b00000000000001110011010001;
    W_in[4][7] = 26'b00000000000000111101101110;
    W_in[4][8] = 26'b11111111111100100000101110;
    W_in[4][9] = 26'b00000000000000010110011000;
    W_in[4][10] = 26'b00000000000011111010111111;
    W_in[4][11] = 26'b11111111111111111110101100;
    W_in[4][12] = 26'b00000000000010011111111001;
    W_in[4][13] = 26'b00000000000000101100000000;
    W_in[4][14] = 26'b00000000000000100111011101;
    W_in[4][15] = 26'b00000000000010111001011010;
    W_in[4][16] = 26'b11111111111111100000000101;
    W_in[4][17] = 26'b00000000000011011100110111;
    W_in[4][18] = 26'b11111111111111100011001001;
    W_in[4][19] = 26'b00000000000010010001001011;
    W_in[4][20] = 26'b11111111111111100001111100;
    W_in[4][21] = 26'b00000000000010000111001000;
    W_in[4][22] = 26'b00000000000001100001111111;
    W_in[4][23] = 26'b00000000000001100011100000;
    W_in[4][24] = 26'b11111111111101011110111110;
    W_in[4][25] = 26'b00000000000001111000001100;
    W_in[4][26] = 26'b00000000000010001011100110;
    W_in[4][27] = 26'b00000000000001011011010101;
    W_in[4][28] = 26'b00000000000011100010100110;
    W_in[4][29] = 26'b11111111111100101100001011;
    W_in[4][30] = 26'b11111111111110110101100001;
    W_in[4][31] = 26'b00000000000001100111000001;
    W_in[4][32] = 26'b00000000000000110001101110;
    W_in[4][33] = 26'b00000000000001111010001100;
    W_in[4][34] = 26'b00000000000001111010011110;
    W_in[4][35] = 26'b00000000000000011010111101;
    W_in[4][36] = 26'b00000000000011111110101101;
    W_in[4][37] = 26'b00000000000001010001000000;
    W_in[4][38] = 26'b11111111111110111011001110;
    W_in[4][39] = 26'b00000000000000111101100110;
    W_in[4][40] = 26'b00000000000010010101101000;
    W_in[4][41] = 26'b11111111111101000000111011;
    W_in[4][42] = 26'b00000000000000111100111010;
    W_in[4][43] = 26'b11111111111110100001001011;
    W_in[4][44] = 26'b11111111111111111001001101;
    W_in[4][45] = 26'b11111111111101110010100010;
    W_in[4][46] = 26'b11111111111100111001111111;
    W_in[4][47] = 26'b00000000000011011110110000;
    W_in[4][48] = 26'b11111111111111000101001111;
    W_in[4][49] = 26'b11111111111110011100100001;
    W_in[4][50] = 26'b11111111111111100110010101;
    W_in[4][51] = 26'b00000000000000000001001000;
    W_in[4][52] = 26'b11111111111100011011000001;
    W_in[4][53] = 26'b11111111111110101001001010;
    W_in[4][54] = 26'b00000000000001000011001101;
    W_in[4][55] = 26'b11111111111110011111000000;
    W_in[4][56] = 26'b00000000000010011001010000;
    W_in[4][57] = 26'b11111111111110010101100110;
    W_in[4][58] = 26'b11111111111110101101100110;
    W_in[4][59] = 26'b00000000000010000111111111;
    W_in[4][60] = 26'b11111111111101010100000101;
    W_in[4][61] = 26'b11111111111100110111101111;
    W_in[4][62] = 26'b11111111111100110001111110;
    W_in[4][63] = 26'b00000000000010000101110100;
    W_in[5][0] = 26'b11111111111110001011100101;
    W_in[5][1] = 26'b11111111111110011001011110;
    W_in[5][2] = 26'b00000000000010111111010101;
    W_in[5][3] = 26'b00000000000010010110010001;
    W_in[5][4] = 26'b00000000000000010100010110;
    W_in[5][5] = 26'b00000000000000111110001011;
    W_in[5][6] = 26'b00000000000000110100100011;
    W_in[5][7] = 26'b00000000000000100000111100;
    W_in[5][8] = 26'b00000000000000101000000110;
    W_in[5][9] = 26'b00000000000000100101000110;
    W_in[5][10] = 26'b11111111111111100001110010;
    W_in[5][11] = 26'b11111111111111111110110000;
    W_in[5][12] = 26'b00000000000000101110101111;
    W_in[5][13] = 26'b00000000000001110000000010;
    W_in[5][14] = 26'b11111111111101010110100001;
    W_in[5][15] = 26'b00000000000000100010000110;
    W_in[5][16] = 26'b11111111111111111111010101;
    W_in[5][17] = 26'b11111111111111111100011011;
    W_in[5][18] = 26'b11111111111111110010001110;
    W_in[5][19] = 26'b11111111111110101111110011;
    W_in[5][20] = 26'b11111111111111110000001110;
    W_in[5][21] = 26'b00000000000000101101101100;
    W_in[5][22] = 26'b11111111111111000000000101;
    W_in[5][23] = 26'b11111111111110100000000011;
    W_in[5][24] = 26'b00000000000000000001010010;
    W_in[5][25] = 26'b00000000000010111010010000;
    W_in[5][26] = 26'b11111111111100110010100110;
    W_in[5][27] = 26'b11111111111100111010100001;
    W_in[5][28] = 26'b00000000000011010110011111;
    W_in[5][29] = 26'b00000000000001000001001111;
    W_in[5][30] = 26'b00000000000000001110100011;
    W_in[5][31] = 26'b11111111111111111101101000;
    W_in[5][32] = 26'b11111111111110000101001001;
    W_in[5][33] = 26'b11111111111111110100011111;
    W_in[5][34] = 26'b11111111111111101101010000;
    W_in[5][35] = 26'b00000000000000001111000011;
    W_in[5][36] = 26'b00000000000000111110110001;
    W_in[5][37] = 26'b00000000000000100100010101;
    W_in[5][38] = 26'b00000000000000110010010010;
    W_in[5][39] = 26'b00000000000010000000010101;
    W_in[5][40] = 26'b00000000000001001101001111;
    W_in[5][41] = 26'b00000000000000000001100100;
    W_in[5][42] = 26'b11111111111111110101010000;
    W_in[5][43] = 26'b00000000000001000000110101;
    W_in[5][44] = 26'b00000000000000011000101010;
    W_in[5][45] = 26'b00000000000000110010011110;
    W_in[5][46] = 26'b11111111111111110011101111;
    W_in[5][47] = 26'b11111111111111011100010110;
    W_in[5][48] = 26'b11111111111111011011011100;
    W_in[5][49] = 26'b11111111111100101011101001;
    W_in[5][50] = 26'b00000000000001111010010100;
    W_in[5][51] = 26'b00000000000010101010101011;
    W_in[5][52] = 26'b11111111111111001110000110;
    W_in[5][53] = 26'b11111111111110011101101001;
    W_in[5][54] = 26'b11111111111110100000000001;
    W_in[5][55] = 26'b11111111111110010011011010;
    W_in[5][56] = 26'b11111111111111000001100011;
    W_in[5][57] = 26'b00000000000011001011011010;
    W_in[5][58] = 26'b00000000000001110111010000;
    W_in[5][59] = 26'b11111111111101111100010111;
    W_in[5][60] = 26'b11111111111111011110011011;
    W_in[5][61] = 26'b11111111111111001001101000;
    W_in[5][62] = 26'b00000000000010101100001010;
    W_in[5][63] = 26'b11111111111110011110111110;
    W_in[6][0] = 26'b11111111111110100100011111;
    W_in[6][1] = 26'b11111111111111000000011100;
    W_in[6][2] = 26'b11111111111100100110000011;
    W_in[6][3] = 26'b11111111111101111000110111;
    W_in[6][4] = 26'b11111111111110110101100100;
    W_in[6][5] = 26'b11111111111111011101011011;
    W_in[6][6] = 26'b00000000000000010111100001;
    W_in[6][7] = 26'b11111111111101011101100010;
    W_in[6][8] = 26'b11111111111111010100001101;
    W_in[6][9] = 26'b11111111111111010110000101;
    W_in[6][10] = 26'b11111111111111010000011101;
    W_in[6][11] = 26'b11111111111100010110011101;
    W_in[6][12] = 26'b11111111111111011010111101;
    W_in[6][13] = 26'b00000000000000110111100010;
    W_in[6][14] = 26'b11111111111111010100001001;
    W_in[6][15] = 26'b00000000000001010111110110;
    W_in[6][16] = 26'b11111111111101011001111110;
    W_in[6][17] = 26'b00000000000011100101011000;
    W_in[6][18] = 26'b00000000000000001100000001;
    W_in[6][19] = 26'b00000000000001001011110100;
    W_in[6][20] = 26'b00000000000000110111101110;
    W_in[6][21] = 26'b11111111111110110111111000;
    W_in[6][22] = 26'b00000000000001110111110011;
    W_in[6][23] = 26'b00000000000011010011111011;
    W_in[6][24] = 26'b00000000000001101100000010;
    W_in[6][25] = 26'b00000000000000100011010011;
    W_in[6][26] = 26'b11111111111111110000001111;
    W_in[6][27] = 26'b11111111111100101101101100;
    W_in[6][28] = 26'b11111111111111000011110001;
    W_in[6][29] = 26'b00000000000011110001010100;
    W_in[6][30] = 26'b11111111111110011111111010;
    W_in[6][31] = 26'b11111111111110100001000010;
    W_in[6][32] = 26'b00000000000000001010110100;
    W_in[6][33] = 26'b00000000000001011011110101;
    W_in[6][34] = 26'b11111111111111010001001101;
    W_in[6][35] = 26'b11111111111111001001110111;
    W_in[6][36] = 26'b00000000000000001100001111;
    W_in[6][37] = 26'b00000000000000101010010111;
    W_in[6][38] = 26'b00000000000010000000001100;
    W_in[6][39] = 26'b11111111111111111110101010;
    W_in[6][40] = 26'b00000000000001110001111000;
    W_in[6][41] = 26'b11111111111111001010101010;
    W_in[6][42] = 26'b00000000000001110110010111;
    W_in[6][43] = 26'b11111111111111110011001010;
    W_in[6][44] = 26'b00000000000000101100111111;
    W_in[6][45] = 26'b00000000000000111111010011;
    W_in[6][46] = 26'b00000000000000110001111000;
    W_in[6][47] = 26'b00000000000000011001111101;
    W_in[6][48] = 26'b00000000000000110011100010;
    W_in[6][49] = 26'b00000000000000101011010101;
    W_in[6][50] = 26'b11111111111110000101111111;
    W_in[6][51] = 26'b00000000000001010111000001;
    W_in[6][52] = 26'b00000000000001010001111110;
    W_in[6][53] = 26'b00000000000000111001000101;
    W_in[6][54] = 26'b11111111111100100101001000;
    W_in[6][55] = 26'b00000000000001001011001000;
    W_in[6][56] = 26'b00000000000000110010000111;
    W_in[6][57] = 26'b11111111111101011100111010;
    W_in[6][58] = 26'b11111111111110000111101110;
    W_in[6][59] = 26'b11111111111110010110010101;
    W_in[6][60] = 26'b00000000000010011001011000;
    W_in[6][61] = 26'b00000000000001000110001101;
    W_in[6][62] = 26'b00000000000010011111001000;
    W_in[6][63] = 26'b00000000000100011010010100;
    W_in[7][0] = 26'b11111111111111110111011110;
    W_in[7][1] = 26'b00000000000011111101100001;
    W_in[7][2] = 26'b00000000000000000000100000;
    W_in[7][3] = 26'b00000000000011001010011110;
    W_in[7][4] = 26'b11111111111101001000000010;
    W_in[7][5] = 26'b00000000000000101001011000;
    W_in[7][6] = 26'b00000000000000011110100000;
    W_in[7][7] = 26'b11111111111110110011010110;
    W_in[7][8] = 26'b11111111111111100011001101;
    W_in[7][9] = 26'b00000000000010100110101101;
    W_in[7][10] = 26'b11111111111110001001101000;
    W_in[7][11] = 26'b11111111111111101001111110;
    W_in[7][12] = 26'b11111111111101111110100110;
    W_in[7][13] = 26'b11111111111111010100101010;
    W_in[7][14] = 26'b11111111111111000111101011;
    W_in[7][15] = 26'b11111111111111100011000101;
    W_in[7][16] = 26'b00000000000000001001101100;
    W_in[7][17] = 26'b00000000000000101010110110;
    W_in[7][18] = 26'b11111111111110100111000111;
    W_in[7][19] = 26'b00000000000010000001111100;
    W_in[7][20] = 26'b11111111111111001100000011;
    W_in[7][21] = 26'b00000000000000110011010100;
    W_in[7][22] = 26'b00000000000001010100011010;
    W_in[7][23] = 26'b00000000000000110110011111;
    W_in[7][24] = 26'b00000000000011010100010011;
    W_in[7][25] = 26'b00000000000000101110100101;
    W_in[7][26] = 26'b11111111111111100010000100;
    W_in[7][27] = 26'b11111111111110110010101011;
    W_in[7][28] = 26'b00000000000000101101010001;
    W_in[7][29] = 26'b00000000000000100110001010;
    W_in[7][30] = 26'b11111111111101111000000011;
    W_in[7][31] = 26'b00000000000100001000111101;
    W_in[7][32] = 26'b00000000000010000111110010;
    W_in[7][33] = 26'b11111111111101100010011101;
    W_in[7][34] = 26'b00000000000001000000001100;
    W_in[7][35] = 26'b00000000000000100100110100;
    W_in[7][36] = 26'b00000000000000101110111111;
    W_in[7][37] = 26'b11111111111100011111101010;
    W_in[7][38] = 26'b00000000000001100010010000;
    W_in[7][39] = 26'b00000000000000001110011010;
    W_in[7][40] = 26'b11111111111111111011010001;
    W_in[7][41] = 26'b00000000000010010101010100;
    W_in[7][42] = 26'b11111111111101011000110011;
    W_in[7][43] = 26'b00000000000000011000001110;
    W_in[7][44] = 26'b11111111111110100111111100;
    W_in[7][45] = 26'b11111111111110111000100101;
    W_in[7][46] = 26'b00000000000011000101110111;
    W_in[7][47] = 26'b11111111111110100011100010;
    W_in[7][48] = 26'b11111111111111001010000110;
    W_in[7][49] = 26'b11111111111111011001100010;
    W_in[7][50] = 26'b11111111111110001111111010;
    W_in[7][51] = 26'b11111111111110100000010011;
    W_in[7][52] = 26'b11111111111110010111100111;
    W_in[7][53] = 26'b11111111111110001011010010;
    W_in[7][54] = 26'b11111111111110111101100001;
    W_in[7][55] = 26'b11111111111100011000001000;
    W_in[7][56] = 26'b11111111111110010011001000;
    W_in[7][57] = 26'b00000000000001111100111001;
    W_in[7][58] = 26'b11111111111101110011100010;
    W_in[7][59] = 26'b11111111111110011100011110;
    W_in[7][60] = 26'b11111111111110011111111101;
    W_in[7][61] = 26'b11111111111110101101010110;
    W_in[7][62] = 26'b11111111111101000001000110;
    W_in[7][63] = 26'b11111111111110110000001010;
    W_in[8][0] = 26'b11111111111111110010000001;
    W_in[8][1] = 26'b11111111111111001101101000;
    W_in[8][2] = 26'b11111111111111011010110110;
    W_in[8][3] = 26'b11111111111110011100111100;
    W_in[8][4] = 26'b00000000000000000101000010;
    W_in[8][5] = 26'b00000000000001011100011001;
    W_in[8][6] = 26'b11111111111110001101011110;
    W_in[8][7] = 26'b11111111111101011101000111;
    W_in[8][8] = 26'b11111111111100010100000010;
    W_in[8][9] = 26'b11111111111110100101100101;
    W_in[8][10] = 26'b11111111111100101110000101;
    W_in[8][11] = 26'b11111111111110111100001000;
    W_in[8][12] = 26'b11111111111111011010011000;
    W_in[8][13] = 26'b00000000000001011100001011;
    W_in[8][14] = 26'b00000000000000011001001001;
    W_in[8][15] = 26'b11111111111111011010010100;
    W_in[8][16] = 26'b11111111111110000011001110;
    W_in[8][17] = 26'b11111111111110100010010111;
    W_in[8][18] = 26'b11111111111110000110011001;
    W_in[8][19] = 26'b11111111111101101010011010;
    W_in[8][20] = 26'b11111111111111011100100001;
    W_in[8][21] = 26'b00000000000001101011001101;
    W_in[8][22] = 26'b00000000000100001110110100;
    W_in[8][23] = 26'b00000000000010010101111110;
    W_in[8][24] = 26'b11111111111100100000100101;
    W_in[8][25] = 26'b11111111111101001011010011;
    W_in[8][26] = 26'b00000000000000001110100110;
    W_in[8][27] = 26'b11111111111100100000010111;
    W_in[8][28] = 26'b00000000000010111110010001;
    W_in[8][29] = 26'b11111111111111110110101110;
    W_in[8][30] = 26'b00000000000010110101110111;
    W_in[8][31] = 26'b11111111111110000100100100;
    W_in[8][32] = 26'b11111111111100101111111111;
    W_in[8][33] = 26'b11111111111101001010101110;
    W_in[8][34] = 26'b11111111111110000110001111;
    W_in[8][35] = 26'b11111111111101111011100100;
    W_in[8][36] = 26'b11111111111100110110011101;
    W_in[8][37] = 26'b11111111111101010101011100;
    W_in[8][38] = 26'b11111111111110010010000110;
    W_in[8][39] = 26'b00000000000001000100110110;
    W_in[8][40] = 26'b00000000000000101111111011;
    W_in[8][41] = 26'b11111111111110001100011101;
    W_in[8][42] = 26'b11111111111111101111100111;
    W_in[8][43] = 26'b11111111111110100111101001;
    W_in[8][44] = 26'b11111111111100001000111000;
    W_in[8][45] = 26'b11111111111111010101111011;
    W_in[8][46] = 26'b11111111111111010101001001;
    W_in[8][47] = 26'b11111111111111100001011001;
    W_in[8][48] = 26'b00000000000000000000100110;
    W_in[8][49] = 26'b11111111111111001001110110;
    W_in[8][50] = 26'b00000000000010100111001011;
    W_in[8][51] = 26'b11111111111110011011111001;
    W_in[8][52] = 26'b00000000000011101010001011;
    W_in[8][53] = 26'b00000000000001110001010000;
    W_in[8][54] = 26'b00000000000011110110001001;
    W_in[8][55] = 26'b00000000000011001101011001;
    W_in[8][56] = 26'b00000000000001010000010001;
    W_in[8][57] = 26'b11111111111100100001110111;
    W_in[8][58] = 26'b00000000000010000011010101;
    W_in[8][59] = 26'b00000000000110111011010000;
    W_in[8][60] = 26'b00000000000101001011001100;
    W_in[8][61] = 26'b00000000000101011101011000;
    W_in[8][62] = 26'b00000000000110011100100010;
    W_in[8][63] = 26'b00000000000101110000001010;
    W_in[9][0] = 26'b00000000000000101010000111;
    W_in[9][1] = 26'b00000000000000101101010100;
    W_in[9][2] = 26'b00000000000000110101100001;
    W_in[9][3] = 26'b11111111111111100000111000;
    W_in[9][4] = 26'b11111111111111011101011111;
    W_in[9][5] = 26'b11111111111101101100001000;
    W_in[9][6] = 26'b00000000000011000111010101;
    W_in[9][7] = 26'b11111111111100010101001110;
    W_in[9][8] = 26'b11111111111101001001110110;
    W_in[9][9] = 26'b11111111111110111101100010;
    W_in[9][10] = 26'b11111111111111111010100011;
    W_in[9][11] = 26'b11111111111111011010011110;
    W_in[9][12] = 26'b11111111111101110000101010;
    W_in[9][13] = 26'b11111111111111010110000100;
    W_in[9][14] = 26'b11111111111110000011110001;
    W_in[9][15] = 26'b11111111111101111111011000;
    W_in[9][16] = 26'b00000000000010010011111000;
    W_in[9][17] = 26'b11111111111101011111000101;
    W_in[9][18] = 26'b00000000000000011110111101;
    W_in[9][19] = 26'b11111111111100110111101110;
    W_in[9][20] = 26'b11111111111111011000000100;
    W_in[9][21] = 26'b00000000000000000101011010;
    W_in[9][22] = 26'b00000000000001010010011110;
    W_in[9][23] = 26'b00000000000000110011011011;
    W_in[9][24] = 26'b11111111111111101011111101;
    W_in[9][25] = 26'b11111111111110011110011011;
    W_in[9][26] = 26'b11111111111111101100111100;
    W_in[9][27] = 26'b00000000000001011100110100;
    W_in[9][28] = 26'b00000000000000010100000001;
    W_in[9][29] = 26'b11111111111110001010000010;
    W_in[9][30] = 26'b11111111111111000100001110;
    W_in[9][31] = 26'b11111111111100100010000100;
    W_in[9][32] = 26'b11111111111111110001011001;
    W_in[9][33] = 26'b11111111111100000000010010;
    W_in[9][34] = 26'b11111111111110111111011000;
    W_in[9][35] = 26'b00000000000001111100100101;
    W_in[9][36] = 26'b11111111111110000001111110;
    W_in[9][37] = 26'b11111111111101000100011101;
    W_in[9][38] = 26'b11111111111011101001010010;
    W_in[9][39] = 26'b00000000000010100011011110;
    W_in[9][40] = 26'b11111111111110101110101000;
    W_in[9][41] = 26'b11111111111111011111111101;
    W_in[9][42] = 26'b00000000000000001101101101;
    W_in[9][43] = 26'b11111111111110100110001100;
    W_in[9][44] = 26'b00000000000000100001000111;
    W_in[9][45] = 26'b11111111111110101001111111;
    W_in[9][46] = 26'b11111111111111011011001100;
    W_in[9][47] = 26'b00000000000001111010001001;
    W_in[9][48] = 26'b00000000000000111100110111;
    W_in[9][49] = 26'b00000000000000110010000100;
    W_in[9][50] = 26'b00000000000000101010101010;
    W_in[9][51] = 26'b00000000000000101100011101;
    W_in[9][52] = 26'b11111111111110111011001001;
    W_in[9][53] = 26'b11111111111110101101110111;
    W_in[9][54] = 26'b00000000000000111010100100;
    W_in[9][55] = 26'b00000000000000000000101010;
    W_in[9][56] = 26'b00000000000000101100001011;
    W_in[9][57] = 26'b11111111111101101111011110;
    W_in[9][58] = 26'b11111111111101111001100110;
    W_in[9][59] = 26'b11111111111110110110001001;
    W_in[9][60] = 26'b00000000000011101110101010;
    W_in[9][61] = 26'b00000000000010100001110101;
    W_in[9][62] = 26'b11111111111110110000001100;
    W_in[9][63] = 26'b00000000000010010000110110;
    W_in[10][0] = 26'b00000000000010111010101011;
    W_in[10][1] = 26'b11111111111111001110101111;
    W_in[10][2] = 26'b00000000000100101011010000;
    W_in[10][3] = 26'b11111111111110110011011101;
    W_in[10][4] = 26'b00000000000010100111110011;
    W_in[10][5] = 26'b00000000000000100111010110;
    W_in[10][6] = 26'b11111111111100101100000111;
    W_in[10][7] = 26'b00000000000100101100001101;
    W_in[10][8] = 26'b00000000000101011000111110;
    W_in[10][9] = 26'b00000000000011001010011111;
    W_in[10][10] = 26'b00000000000011110110101100;
    W_in[10][11] = 26'b11111111111111111010000001;
    W_in[10][12] = 26'b00000000000000000011010001;
    W_in[10][13] = 26'b00000000000001001010011001;
    W_in[10][14] = 26'b11111111111110110111110100;
    W_in[10][15] = 26'b11111111111100101110000111;
    W_in[10][16] = 26'b11111111111110101001000111;
    W_in[10][17] = 26'b00000000000010011101100000;
    W_in[10][18] = 26'b11111111111111111010010001;
    W_in[10][19] = 26'b11111111111111110100101100;
    W_in[10][20] = 26'b11111111111111010001011000;
    W_in[10][21] = 26'b11111111111101010101011001;
    W_in[10][22] = 26'b00000000000100010110000011;
    W_in[10][23] = 26'b11111111111111110101110100;
    W_in[10][24] = 26'b11111111111101011101001010;
    W_in[10][25] = 26'b00000000000001010000101100;
    W_in[10][26] = 26'b11111111111101001111000100;
    W_in[10][27] = 26'b11111111111101111000000010;
    W_in[10][28] = 26'b00000000000011000011010010;
    W_in[10][29] = 26'b00000000000010101000111011;
    W_in[10][30] = 26'b11111111111101011000001111;
    W_in[10][31] = 26'b00000000000010011001111111;
    W_in[10][32] = 26'b00000000000000001101011100;
    W_in[10][33] = 26'b00000000000001010000110010;
    W_in[10][34] = 26'b00000000000011010110101011;
    W_in[10][35] = 26'b00000000000100000001010000;
    W_in[10][36] = 26'b11111111111111101100010001;
    W_in[10][37] = 26'b00000000000000111110101110;
    W_in[10][38] = 26'b11111111111100000101101011;
    W_in[10][39] = 26'b11111111111111100110101101;
    W_in[10][40] = 26'b00000000000001111111101000;
    W_in[10][41] = 26'b11111111111110011101111111;
    W_in[10][42] = 26'b00000000000100011011110001;
    W_in[10][43] = 26'b00000000000001000011110111;
    W_in[10][44] = 26'b00000000000010001000010001;
    W_in[10][45] = 26'b11111111111110001010001111;
    W_in[10][46] = 26'b11111111111100101110011001;
    W_in[10][47] = 26'b00000000000011111111110000;
    W_in[10][48] = 26'b11111111111101000000100001;
    W_in[10][49] = 26'b11111111111110001001000011;
    W_in[10][50] = 26'b00000000000010000000110001;
    W_in[10][51] = 26'b11111111111111101101011001;
    W_in[10][52] = 26'b00000000000010001000001110;
    W_in[10][53] = 26'b11111111111001001011110000;
    W_in[10][54] = 26'b11111111111111000101010110;
    W_in[10][55] = 26'b00000000000000100110010010;
    W_in[10][56] = 26'b11111111111101100101010011;
    W_in[10][57] = 26'b11111111111110111000010100;
    W_in[10][58] = 26'b11111111111101011100000011;
    W_in[10][59] = 26'b11111111111101000001111101;
    W_in[10][60] = 26'b11111111111111000101011100;
    W_in[10][61] = 26'b11111111111001110111111000;
    W_in[10][62] = 26'b11111111111000100111111011;
    W_in[10][63] = 26'b11111111111000001011111000;
    W_in[11][0] = 26'b11111111111010100101000101;
    W_in[11][1] = 26'b11111111111010011000010011;
    W_in[11][2] = 26'b00000000000001100011101001;
    W_in[11][3] = 26'b11111111111111001100010011;
    W_in[11][4] = 26'b00000000000011000110100010;
    W_in[11][5] = 26'b00000000000100001111001011;
    W_in[11][6] = 26'b11111111111100100101011000;
    W_in[11][7] = 26'b00000000000000110100001001;
    W_in[11][8] = 26'b11111111111101011101100010;
    W_in[11][9] = 26'b11111111111001110010100100;
    W_in[11][10] = 26'b11111111111101110111010100;
    W_in[11][11] = 26'b00000000000010011110010110;
    W_in[11][12] = 26'b00000000000010111111000111;
    W_in[11][13] = 26'b11111111111101001101010100;
    W_in[11][14] = 26'b00000000000011000001110011;
    W_in[11][15] = 26'b11111111111111111111011001;
    W_in[11][16] = 26'b00000000000000100111100110;
    W_in[11][17] = 26'b11111111111110011111111101;
    W_in[11][18] = 26'b00000000000000100110111101;
    W_in[11][19] = 26'b00000000000011101011001011;
    W_in[11][20] = 26'b11111111111110001111101111;
    W_in[11][21] = 26'b11111111111110100010011001;
    W_in[11][22] = 26'b00000000000011111101010101;
    W_in[11][23] = 26'b11111111111110010100110100;
    W_in[11][24] = 26'b00000000000011100100001111;
    W_in[11][25] = 26'b00000000000001101110001100;
    W_in[11][26] = 26'b00000000000010001010100010;
    W_in[11][27] = 26'b11111111111111000111000010;
    W_in[11][28] = 26'b00000000000010110101010000;
    W_in[11][29] = 26'b00000000000100010000111110;
    W_in[11][30] = 26'b00000000000010110010010001;
    W_in[11][31] = 26'b00000000000001011111110010;
    W_in[11][32] = 26'b11111111111101011100110010;
    W_in[11][33] = 26'b11111111111110011101100110;
    W_in[11][34] = 26'b11111111111010001110110110;
    W_in[11][35] = 26'b11111111111100110100101001;
    W_in[11][36] = 26'b00000000000011110010010010;
    W_in[11][37] = 26'b00000000000000000010001101;
    W_in[11][38] = 26'b00000000000011001100111110;
    W_in[11][39] = 26'b11111111111011101111101011;
    W_in[11][40] = 26'b11111111111111110110110001;
    W_in[11][41] = 26'b11111111111011110111111001;
    W_in[11][42] = 26'b11111111111011100110100100;
    W_in[11][43] = 26'b11111111111011011100000110;
    W_in[11][44] = 26'b11111111111101101010000110;
    W_in[11][45] = 26'b00000000000000100110011110;
    W_in[11][46] = 26'b00000000001000110000011011;
    W_in[11][47] = 26'b11111111111101101001010101;
    W_in[11][48] = 26'b11111111111111100110110011;
    W_in[11][49] = 26'b11111111111101011001110101;
    W_in[11][50] = 26'b11111111111100001001111100;
    W_in[11][51] = 26'b00000000000101110110001100;
    W_in[11][52] = 26'b11111111111011101001101110;
    W_in[11][53] = 26'b00000000000001011000101100;
    W_in[11][54] = 26'b00000000000100011011111011;
    W_in[11][55] = 26'b00000000000000101101000100;
    W_in[11][56] = 26'b00000000001001000101101110;
    W_in[11][57] = 26'b00000000000001001001101001;
    W_in[11][58] = 26'b00000000001001010001010100;
    W_in[11][59] = 26'b00000000000001011110100011;
    W_in[11][60] = 26'b11111111111100001001110101;
    W_in[11][61] = 26'b00000000000100011100000101;
    W_in[11][62] = 26'b00000000000110000001100100;
    W_in[11][63] = 26'b11111111111100001001111000;
    W_in[12][0] = 26'b11111111111110001110100011;
    W_in[12][1] = 26'b00000000000000111101111100;
    W_in[12][2] = 26'b11111111111111001100010000;
    W_in[12][3] = 26'b00000000000010001101110100;
    W_in[12][4] = 26'b11111111111111011001001100;
    W_in[12][5] = 26'b11111111111110111001011101;
    W_in[12][6] = 26'b11111111111100100000000111;
    W_in[12][7] = 26'b11111111111110000110100000;
    W_in[12][8] = 26'b11111111111110111010010110;
    W_in[12][9] = 26'b00000000000010010110010110;
    W_in[12][10] = 26'b00000000000001000101101010;
    W_in[12][11] = 26'b00000000000011011101110110;
    W_in[12][12] = 26'b11111111111111000100010000;
    W_in[12][13] = 26'b00000000000001110011000110;
    W_in[12][14] = 26'b00000000000001110001111010;
    W_in[12][15] = 26'b00000000000000110000101010;
    W_in[12][16] = 26'b11111111111111010110011010;
    W_in[12][17] = 26'b00000000000010101110101111;
    W_in[12][18] = 26'b00000000000011111111000010;
    W_in[12][19] = 26'b00000000000010001101110110;
    W_in[12][20] = 26'b11111111111111100110101111;
    W_in[12][21] = 26'b00000000000000101110110100;
    W_in[12][22] = 26'b00000000000010110001101110;
    W_in[12][23] = 26'b00000000000000101000000010;
    W_in[12][24] = 26'b00000000000000001111011101;
    W_in[12][25] = 26'b11111111111111010100011000;
    W_in[12][26] = 26'b11111111111100010011001011;
    W_in[12][27] = 26'b00000000000000110101111110;
    W_in[12][28] = 26'b00000000000001111100110010;
    W_in[12][29] = 26'b00000000000000001010111011;
    W_in[12][30] = 26'b00000000000010011110011010;
    W_in[12][31] = 26'b00000000000010000111010100;
    W_in[12][32] = 26'b11111111111111011011000101;
    W_in[12][33] = 26'b11111111111101101111100111;
    W_in[12][34] = 26'b11111111111100111000000100;
    W_in[12][35] = 26'b11111111111110011101101011;
    W_in[12][36] = 26'b11111111111110010001001110;
    W_in[12][37] = 26'b11111111111010110100100100;
    W_in[12][38] = 26'b00000000000000111000111111;
    W_in[12][39] = 26'b11111111111111101110010000;
    W_in[12][40] = 26'b11111111111111010010111011;
    W_in[12][41] = 26'b00000000000011011010111011;
    W_in[12][42] = 26'b11111111111101010111001111;
    W_in[12][43] = 26'b00000000000010001010111000;
    W_in[12][44] = 26'b00000000000000000001011110;
    W_in[12][45] = 26'b11111111111110000001111011;
    W_in[12][46] = 26'b11111111111101101010011100;
    W_in[12][47] = 26'b00000000000010101011101110;
    W_in[12][48] = 26'b00000000000001000110010011;
    W_in[12][49] = 26'b00000000000100101110100101;
    W_in[12][50] = 26'b11111111111111111111000110;
    W_in[12][51] = 26'b00000000000000111101101001;
    W_in[12][52] = 26'b11111111111110110101000101;
    W_in[12][53] = 26'b11111111111101000111100011;
    W_in[12][54] = 26'b11111111111100101100100011;
    W_in[12][55] = 26'b11111111111110010110111011;
    W_in[12][56] = 26'b00000000000011101100000001;
    W_in[12][57] = 26'b11111111111110110100110100;
    W_in[12][58] = 26'b00000000000011110011100011;
    W_in[12][59] = 26'b11111111111111001000010111;
    W_in[12][60] = 26'b11111111111011101000101001;
    W_in[12][61] = 26'b11111111111001000111111100;
    W_in[12][62] = 26'b11111111111000000011011110;
    W_in[12][63] = 26'b00000000000001101111011100;
    W_in[13][0] = 26'b00000000000011001011001011;
    W_in[13][1] = 26'b00000000000001000110010100;
    W_in[13][2] = 26'b00000000000000101101100111;
    W_in[13][3] = 26'b00000000000000000011001001;
    W_in[13][4] = 26'b00000000000000011110111010;
    W_in[13][5] = 26'b00000000000010011010001010;
    W_in[13][6] = 26'b11111111111100110100011101;
    W_in[13][7] = 26'b11111111111101011010001101;
    W_in[13][8] = 26'b00000000000000000100111010;
    W_in[13][9] = 26'b00000000000100000010001010;
    W_in[13][10] = 26'b00000000000010000100111110;
    W_in[13][11] = 26'b11111111111011110010010001;
    W_in[13][12] = 26'b11111111111101011011110011;
    W_in[13][13] = 26'b00000000000010101110000101;
    W_in[13][14] = 26'b11111111111111001010110010;
    W_in[13][15] = 26'b00000000000011001101001011;
    W_in[13][16] = 26'b11111111111100001110001001;
    W_in[13][17] = 26'b00000000000001110110101110;
    W_in[13][18] = 26'b00000000000100100010000101;
    W_in[13][19] = 26'b11111111111101010000110110;
    W_in[13][20] = 26'b11111111111101100110010111;
    W_in[13][21] = 26'b11111111111100010000011111;
    W_in[13][22] = 26'b00000000000010001101100001;
    W_in[13][23] = 26'b00000000000101001111010111;
    W_in[13][24] = 26'b00000000000001111011111000;
    W_in[13][25] = 26'b11111111111110000101010011;
    W_in[13][26] = 26'b11111111111110011000000111;
    W_in[13][27] = 26'b11111111111101111010111001;
    W_in[13][28] = 26'b11111111111110101001110010;
    W_in[13][29] = 26'b11111111111100110110000111;
    W_in[13][30] = 26'b11111111111111000111010000;
    W_in[13][31] = 26'b11111111111100110011011011;
    W_in[13][32] = 26'b00000000000010011100111000;
    W_in[13][33] = 26'b11111111111110111110010111;
    W_in[13][34] = 26'b11111111111101111110001100;
    W_in[13][35] = 26'b00000000000010100101101001;
    W_in[13][36] = 26'b11111111111011011011011111;
    W_in[13][37] = 26'b00000000000000101001110101;
    W_in[13][38] = 26'b11111111111111111000110010;
    W_in[13][39] = 26'b11111111111101111110000000;
    W_in[13][40] = 26'b00000000000010110110011011;
    W_in[13][41] = 26'b00000000000001011011111100;
    W_in[13][42] = 26'b00000000000011101111110000;
    W_in[13][43] = 26'b00000000000011001101101111;
    W_in[13][44] = 26'b00000000000000001100010111;
    W_in[13][45] = 26'b00000000000011101010100001;
    W_in[13][46] = 26'b00000000000001000001010000;
    W_in[13][47] = 26'b11111111111111001001011100;
    W_in[13][48] = 26'b11111111111101000101000100;
    W_in[13][49] = 26'b11111111111111011010111110;
    W_in[13][50] = 26'b11111111111110010100101101;
    W_in[13][51] = 26'b00000000000001110100100011;
    W_in[13][52] = 26'b00000000000010101110000101;
    W_in[13][53] = 26'b00000000000001100010000010;
    W_in[13][54] = 26'b11111111111100001011111111;
    W_in[13][55] = 26'b00000000000100110010111100;
    W_in[13][56] = 26'b00000000000010011010001101;
    W_in[13][57] = 26'b11111111111111000010100101;
    W_in[13][58] = 26'b11111111111111101101111110;
    W_in[13][59] = 26'b00000000000011011111000010;
    W_in[13][60] = 26'b11111111111011101110001111;
    W_in[13][61] = 26'b11111111111111110011001001;
    W_in[13][62] = 26'b11111111111110010010000011;
    W_in[13][63] = 26'b11111111111110100000000111;
    W_in[14][0] = 26'b00000000000001011011101000;
    W_in[14][1] = 26'b00000000000001111110011000;
    W_in[14][2] = 26'b11111111111111010000100000;
    W_in[14][3] = 26'b00000000000000110001101001;
    W_in[14][4] = 26'b00000000000011001101001101;
    W_in[14][5] = 26'b00000000000001011001000111;
    W_in[14][6] = 26'b11111111111011011001111100;
    W_in[14][7] = 26'b00000000000001011100100011;
    W_in[14][8] = 26'b11111111111010000011000101;
    W_in[14][9] = 26'b11111111111111001100110111;
    W_in[14][10] = 26'b11111111111111111011010111;
    W_in[14][11] = 26'b11111111111110001111010101;
    W_in[14][12] = 26'b11111111111100100001110101;
    W_in[14][13] = 26'b00000000000001100100110110;
    W_in[14][14] = 26'b11111111111111110010000101;
    W_in[14][15] = 26'b11111111111010100110100111;
    W_in[14][16] = 26'b00000000000010000100010011;
    W_in[14][17] = 26'b00000000000010010100011110;
    W_in[14][18] = 26'b11111111111010000100000010;
    W_in[14][19] = 26'b11111111111011110011011000;
    W_in[14][20] = 26'b00000000000011010011010011;
    W_in[14][21] = 26'b11111111111100110111101000;
    W_in[14][22] = 26'b00000000000001010110100000;
    W_in[14][23] = 26'b11111111111101000001100010;
    W_in[14][24] = 26'b00000000000001100101010001;
    W_in[14][25] = 26'b11111111111101010011011100;
    W_in[14][26] = 26'b00000000000100101011101000;
    W_in[14][27] = 26'b11111111111111001111100111;
    W_in[14][28] = 26'b00000000000010110011111101;
    W_in[14][29] = 26'b00000000000100011011101011;
    W_in[14][30] = 26'b11111111111111011000010001;
    W_in[14][31] = 26'b00000000000000000001001010;
    W_in[14][32] = 26'b00000000000101011011111011;
    W_in[14][33] = 26'b11111111111011111001110010;
    W_in[14][34] = 26'b11111111111100001011101101;
    W_in[14][35] = 26'b11111111111110001011000000;
    W_in[14][36] = 26'b00000000000101000010111001;
    W_in[14][37] = 26'b00000000000100001011011101;
    W_in[14][38] = 26'b11111111111101011010000111;
    W_in[14][39] = 26'b11111111111010101110101100;
    W_in[14][40] = 26'b00000000000010001101110001;
    W_in[14][41] = 26'b11111111111111101100110101;
    W_in[14][42] = 26'b11111111111100001110011010;
    W_in[14][43] = 26'b00000000000000101100100000;
    W_in[14][44] = 26'b11111111111110101101101100;
    W_in[14][45] = 26'b00000000000010011001111110;
    W_in[14][46] = 26'b11111111111111000111001111;
    W_in[14][47] = 26'b11111111111111000110001101;
    W_in[14][48] = 26'b11111111111110011111100100;
    W_in[14][49] = 26'b11111111111111111100010100;
    W_in[14][50] = 26'b11111111111100001110000101;
    W_in[14][51] = 26'b11111111111110011010011110;
    W_in[14][52] = 26'b11111111111011111011111011;
    W_in[14][53] = 26'b00000000000011011010011011;
    W_in[14][54] = 26'b11111111111111011111111010;
    W_in[14][55] = 26'b11111111111110001110001000;
    W_in[14][56] = 26'b11111111111110010010100100;
    W_in[14][57] = 26'b00000000000011100110100100;
    W_in[14][58] = 26'b00000000000011110111001010;
    W_in[14][59] = 26'b00000000000100110110011110;
    W_in[14][60] = 26'b00000000000111100101011010;
    W_in[14][61] = 26'b00000000000101000101101000;
    W_in[14][62] = 26'b00000000001000101110110110;
    W_in[14][63] = 26'b00000000000110011110011110;
    W_in[15][0] = 26'b11111111111010011000111100;
    W_in[15][1] = 26'b00000000000100000101101011;
    W_in[15][2] = 26'b00000000000000010011010110;
    W_in[15][3] = 26'b00000000000100011011110010;
    W_in[15][4] = 26'b11111111111010111001000111;
    W_in[15][5] = 26'b00000000000001000110101110;
    W_in[15][6] = 26'b11111111111011100001000110;
    W_in[15][7] = 26'b00000000000010011110011111;
    W_in[15][8] = 26'b11111111111001000110111001;
    W_in[15][9] = 26'b11111111111010011000001111;
    W_in[15][10] = 26'b00000000000100101000010100;
    W_in[15][11] = 26'b11111111111010011000101011;
    W_in[15][12] = 26'b11111111111010100011011100;
    W_in[15][13] = 26'b00000000000010010100100010;
    W_in[15][14] = 26'b00000000000001111110100100;
    W_in[15][15] = 26'b00000000000001111111010000;
    W_in[15][16] = 26'b00000000000101010100010001;
    W_in[15][17] = 26'b11111111111110111000110110;
    W_in[15][18] = 26'b11111111111111111110100111;
    W_in[15][19] = 26'b00000000000110010110001100;
    W_in[15][20] = 26'b11111111111111000001111100;
    W_in[15][21] = 26'b11111111111100001110001100;
    W_in[15][22] = 26'b11111111111110100101010101;
    W_in[15][23] = 26'b11111111111110001011010100;
    W_in[15][24] = 26'b11111111111011000010110001;
    W_in[15][25] = 26'b11111111111111000101100011;
    W_in[15][26] = 26'b11111111111011111101100111;
    W_in[15][27] = 26'b11111111111010111111100110;
    W_in[15][28] = 26'b00000000000110100110110010;
    W_in[15][29] = 26'b00000000000010001101101001;
    W_in[15][30] = 26'b00000000000000011001101000;
    W_in[15][31] = 26'b00000000000011101010100011;
    W_in[15][32] = 26'b00000000000010001001111100;
    W_in[15][33] = 26'b11111111111111000000100100;
    W_in[15][34] = 26'b00000000000011100100111101;
    W_in[15][35] = 26'b00000000000001110011010000;
    W_in[15][36] = 26'b11111111111011101111001000;
    W_in[15][37] = 26'b11111111111010110110110111;
    W_in[15][38] = 26'b00000000000010001001011100;
    W_in[15][39] = 26'b11111111111111110100110110;
    W_in[15][40] = 26'b11111111111010000010010101;
    W_in[15][41] = 26'b11111111111010110011000110;
    W_in[15][42] = 26'b00000000000100000101011001;
    W_in[15][43] = 26'b00000000000000010111101011;
    W_in[15][44] = 26'b00000000000001011000101011;
    W_in[15][45] = 26'b00000000000110001110001011;
    W_in[15][46] = 26'b11111111111111011011111101;
    W_in[15][47] = 26'b00000000000101000000101000;
    W_in[15][48] = 26'b00000000000000100110000000;
    W_in[15][49] = 26'b11111111111111011010110100;
    W_in[15][50] = 26'b11111111111101010011011110;
    W_in[15][51] = 26'b00000000000010110011000101;
    W_in[15][52] = 26'b11111111111110110000100011;
    W_in[15][53] = 26'b11111111111010111100011101;
    W_in[15][54] = 26'b00000000000110001000111110;
    W_in[15][55] = 26'b00000000000000111100101001;
    W_in[15][56] = 26'b11111111111101000110100001;
    W_in[15][57] = 26'b00000000000010110101111011;
    W_in[15][58] = 26'b11111111111101100111011111;
    W_in[15][59] = 26'b00000000000101100010100110;
    W_in[15][60] = 26'b00000000000101011101001011;
    W_in[15][61] = 26'b00000000000001010011010000;
    W_in[15][62] = 26'b00000000000000011100100101;
    W_in[15][63] = 26'b00000000000100101111011110;

    // Initialize W_hr weights
    W_hr[0][0] = 26'b00000000000000001110001111;
    W_hr[0][1] = 26'b00000000000000100110100111;
    W_hr[0][2] = 26'b00000000000000111110011110;
    W_hr[0][3] = 26'b11111111111101011100011110;
    W_hr[0][4] = 26'b00000000000100011000010001;
    W_hr[0][5] = 26'b00000000000100101101011110;
    W_hr[0][6] = 26'b00000000000100101010111010;
    W_hr[0][7] = 26'b11111111111011011000011110;
    W_hr[0][8] = 26'b00000000000011111110000011;
    W_hr[0][9] = 26'b00000000000100011111101001;
    W_hr[0][10] = 26'b11111111111101111101110000;
    W_hr[0][11] = 26'b11111111111101100011011100;
    W_hr[0][12] = 26'b00000000000001111101000010;
    W_hr[0][13] = 26'b00000000000010011111110110;
    W_hr[0][14] = 26'b00000000000101101000010000;
    W_hr[0][15] = 26'b11111111111100001101000111;
    W_hr[1][0] = 26'b00000000000011011011110111;
    W_hr[1][1] = 26'b00000000000001110010011111;
    W_hr[1][2] = 26'b11111111111110101100001111;
    W_hr[1][3] = 26'b00000000000010000010011101;
    W_hr[1][4] = 26'b00000000000110100001001011;
    W_hr[1][5] = 26'b11111111111001111001000010;
    W_hr[1][6] = 26'b00000000000000000110101010;
    W_hr[1][7] = 26'b00000000000100011110110101;
    W_hr[1][8] = 26'b00000000000011011001011001;
    W_hr[1][9] = 26'b00000000000000000101010101;
    W_hr[1][10] = 26'b11111111111000001010001111;
    W_hr[1][11] = 26'b00000000000111000111011000;
    W_hr[1][12] = 26'b00000000000101111110111000;
    W_hr[1][13] = 26'b00000000000010001011011110;
    W_hr[1][14] = 26'b11111111111011010011000011;
    W_hr[1][15] = 26'b00000000001010010111010110;
    W_hr[2][0] = 26'b11111111111111010111010000;
    W_hr[2][1] = 26'b11111111111110110011000110;
    W_hr[2][2] = 26'b00000000000010010001100001;
    W_hr[2][3] = 26'b11111111111100110001010111;
    W_hr[2][4] = 26'b11111111111101001011010001;
    W_hr[2][5] = 26'b11111111111111100111010101;
    W_hr[2][6] = 26'b00000000001011101110000101;
    W_hr[2][7] = 26'b11111111111010001000010011;
    W_hr[2][8] = 26'b11111111111111010111001001;
    W_hr[2][9] = 26'b00000000000110110011100000;
    W_hr[2][10] = 26'b00000000001001111100011011;
    W_hr[2][11] = 26'b11111111111001000001001111;
    W_hr[2][12] = 26'b11111111111101011001011001;
    W_hr[2][13] = 26'b11111111111011001100011001;
    W_hr[2][14] = 26'b11111111111100101110000101;
    W_hr[2][15] = 26'b00000000000100111010101011;
    W_hr[3][0] = 26'b00000000000000001110001111;
    W_hr[3][1] = 26'b00000000000000100110100111;
    W_hr[3][2] = 26'b00000000000000111110011110;
    W_hr[3][3] = 26'b11111111111101011100011110;
    W_hr[3][4] = 26'b00000000000100011000010001;
    W_hr[3][5] = 26'b00000000000100101101011110;
    W_hr[3][6] = 26'b00000000000100101010111010;
    W_hr[3][7] = 26'b11111111111011011000011110;
    W_hr[3][8] = 26'b00000000000011111110000011;
    W_hr[3][9] = 26'b00000000000100011111101001;
    W_hr[3][10] = 26'b11111111111101111101110000;
    W_hr[3][11] = 26'b11111111111101100011011100;
    W_hr[3][12] = 26'b00000000000001111101000010;
    W_hr[3][13] = 26'b00000000000010011111110110;
    W_hr[3][14] = 26'b00000000000101101000010000;
    W_hr[3][15] = 26'b11111111111100001101000111;
    W_hr[4][0] = 26'b00000000000011011011110111;
    W_hr[4][1] = 26'b00000000000001110010011111;
    W_hr[4][2] = 26'b11111111111110101100001111;
    W_hr[4][3] = 26'b00000000000010000010011101;
    W_hr[4][4] = 26'b00000000000110100001001011;
    W_hr[4][5] = 26'b11111111111001111001000010;
    W_hr[4][6] = 26'b00000000000000000110101010;
    W_hr[4][7] = 26'b00000000000100011110110101;
    W_hr[4][8] = 26'b00000000000011011001011001;
    W_hr[4][9] = 26'b00000000000000000101010101;
    W_hr[4][10] = 26'b11111111111000001010001111;
    W_hr[4][11] = 26'b00000000000111000111011000;
    W_hr[4][12] = 26'b00000000000101111110111000;
    W_hr[4][13] = 26'b00000000000010001011011110;
    W_hr[4][14] = 26'b11111111111011010011000011;
    W_hr[4][15] = 26'b00000000001010010111010110;
    W_hr[5][0] = 26'b11111111111111010111010000;
    W_hr[5][1] = 26'b11111111111110110011000110;
    W_hr[5][2] = 26'b00000000000010010001100001;
    W_hr[5][3] = 26'b11111111111100110001010111;
    W_hr[5][4] = 26'b11111111111101001011010001;
    W_hr[5][5] = 26'b11111111111111100111010101;
    W_hr[5][6] = 26'b00000000001011101110000101;
    W_hr[5][7] = 26'b11111111111010001000010011;
    W_hr[5][8] = 26'b11111111111111010111001001;
    W_hr[5][9] = 26'b00000000000110110011100000;
    W_hr[5][10] = 26'b00000000001001111100011011;
    W_hr[5][11] = 26'b11111111111001000001001111;
    W_hr[5][12] = 26'b11111111111101011001011001;
    W_hr[5][13] = 26'b11111111111011001100011001;
    W_hr[5][14] = 26'b11111111111100101110000101;
    W_hr[5][15] = 26'b00000000000100111010101011;
    W_hr[6][0] = 26'b00000000000000001110001111;
    W_hr[6][1] = 26'b00000000000000100110100111;
    W_hr[6][2] = 26'b00000000000000111110011110;
    W_hr[6][3] = 26'b11111111111101011100011110;
    W_hr[6][4] = 26'b00000000000100011000010001;
    W_hr[6][5] = 26'b00000000000100101101011110;
    W_hr[6][6] = 26'b00000000000100101010111010;
    W_hr[6][7] = 26'b11111111111011011000011110;
    W_hr[6][8] = 26'b00000000000011111110000011;
    W_hr[6][9] = 26'b00000000000100011111101001;
    W_hr[6][10] = 26'b11111111111101111101110000;
    W_hr[6][11] = 26'b11111111111101100011011100;
    W_hr[6][12] = 26'b00000000000001111101000010;
    W_hr[6][13] = 26'b00000000000010011111110110;
    W_hr[6][14] = 26'b00000000000101101000010000;
    W_hr[6][15] = 26'b11111111111100001101000111;
    W_hr[7][0] = 26'b00000000000011011011110111;
    W_hr[7][1] = 26'b00000000000001110010011111;
    W_hr[7][2] = 26'b11111111111110101100001111;
    W_hr[7][3] = 26'b00000000000010000010011101;
    W_hr[7][4] = 26'b00000000000110100001001011;
    W_hr[7][5] = 26'b11111111111001111001000010;
    W_hr[7][6] = 26'b00000000000000000110101010;
    W_hr[7][7] = 26'b00000000000100011110110101;
    W_hr[7][8] = 26'b00000000000011011001011001;
    W_hr[7][9] = 26'b00000000000000000101010101;
    W_hr[7][10] = 26'b11111111111000001010001111;
    W_hr[7][11] = 26'b00000000000111000111011000;
    W_hr[7][12] = 26'b00000000000101111110111000;
    W_hr[7][13] = 26'b00000000000010001011011110;
    W_hr[7][14] = 26'b11111111111011010011000011;
    W_hr[7][15] = 26'b00000000001010010111010110;
    W_hr[8][0] = 26'b11111111111111010111010000;
    W_hr[8][1] = 26'b11111111111110110011000110;
    W_hr[8][2] = 26'b00000000000010010001100001;
    W_hr[8][3] = 26'b11111111111100110001010111;
    W_hr[8][4] = 26'b11111111111101001011010001;
    W_hr[8][5] = 26'b11111111111111100111010101;
    W_hr[8][6] = 26'b00000000001011101110000101;
    W_hr[8][7] = 26'b11111111111010001000010011;
    W_hr[8][8] = 26'b11111111111111010111001001;
    W_hr[8][9] = 26'b00000000000110110011100000;
    W_hr[8][10] = 26'b00000000001001111100011011;
    W_hr[8][11] = 26'b11111111111001000001001111;
    W_hr[8][12] = 26'b11111111111101011001011001;
    W_hr[8][13] = 26'b11111111111011001100011001;
    W_hr[8][14] = 26'b11111111111100101110000101;
    W_hr[8][15] = 26'b00000000000100111010101011;
    W_hr[9][0] = 26'b00000000000000001110001111;
    W_hr[9][1] = 26'b00000000000000100110100111;
    W_hr[9][2] = 26'b00000000000000111110011110;
    W_hr[9][3] = 26'b11111111111101011100011110;
    W_hr[9][4] = 26'b00000000000100011000010001;
    W_hr[9][5] = 26'b00000000000100101101011110;
    W_hr[9][6] = 26'b00000000000100101010111010;
    W_hr[9][7] = 26'b11111111111011011000011110;
    W_hr[9][8] = 26'b00000000000011111110000011;
    W_hr[9][9] = 26'b00000000000100011111101001;
    W_hr[9][10] = 26'b11111111111101111101110000;
    W_hr[9][11] = 26'b11111111111101100011011100;
    W_hr[9][12] = 26'b00000000000001111101000010;
    W_hr[9][13] = 26'b00000000000010011111110110;
    W_hr[9][14] = 26'b00000000000101101000010000;
    W_hr[9][15] = 26'b11111111111100001101000111;
    W_hr[10][0] = 26'b00000000000011011011110111;
    W_hr[10][1] = 26'b00000000000001110010011111;
    W_hr[10][2] = 26'b11111111111110101100001111;
    W_hr[10][3] = 26'b00000000000010000010011101;
    W_hr[10][4] = 26'b00000000000110100001001011;
    W_hr[10][5] = 26'b11111111111001111001000010;
    W_hr[10][6] = 26'b00000000000000000110101010;
    W_hr[10][7] = 26'b00000000000100011110110101;
    W_hr[10][8] = 26'b00000000000011011001011001;
    W_hr[10][9] = 26'b00000000000000000101010101;
    W_hr[10][10] = 26'b11111111111000001010001111;
    W_hr[10][11] = 26'b00000000000111000111011000;
    W_hr[10][12] = 26'b00000000000101111110111000;
    W_hr[10][13] = 26'b00000000000010001011011110;
    W_hr[10][14] = 26'b11111111111011010011000011;
    W_hr[10][15] = 26'b00000000001010010111010110;
    W_hr[11][0] = 26'b11111111111111010111010000;
    W_hr[11][1] = 26'b11111111111110110011000110;
    W_hr[11][2] = 26'b00000000000010010001100001;
    W_hr[11][3] = 26'b11111111111100110001010111;
    W_hr[11][4] = 26'b11111111111101001011010001;
    W_hr[11][5] = 26'b11111111111111100111010101;
    W_hr[11][6] = 26'b00000000001011101110000101;
    W_hr[11][7] = 26'b11111111111010001000010011;
    W_hr[11][8] = 26'b11111111111111010111001001;
    W_hr[11][9] = 26'b00000000000110110011100000;
    W_hr[11][10] = 26'b00000000001001111100011011;
    W_hr[11][11] = 26'b11111111111001000001001111;
    W_hr[11][12] = 26'b11111111111101011001011001;
    W_hr[11][13] = 26'b11111111111011001100011001;
    W_hr[11][14] = 26'b11111111111100101110000101;
    W_hr[11][15] = 26'b00000000000100111010101011;
    W_hr[12][0] = 26'b00000000000000001110001111;
    W_hr[12][1] = 26'b00000000000000100110100111;
    W_hr[12][2] = 26'b00000000000000111110011110;
    W_hr[12][3] = 26'b11111111111101011100011110;
    W_hr[12][4] = 26'b00000000000100011000010001;
    W_hr[12][5] = 26'b00000000000100101101011110;
    W_hr[12][6] = 26'b00000000000100101010111010;
    W_hr[12][7] = 26'b11111111111011011000011110;
    W_hr[12][8] = 26'b00000000000011111110000011;
    W_hr[12][9] = 26'b00000000000100011111101001;
    W_hr[12][10] = 26'b11111111111101111101110000;
    W_hr[12][11] = 26'b11111111111101100011011100;
    W_hr[12][12] = 26'b00000000000001111101000010;
    W_hr[12][13] = 26'b00000000000010011111110110;
    W_hr[12][14] = 26'b00000000000101101000010000;
    W_hr[12][15] = 26'b11111111111100001101000111;
    W_hr[13][0] = 26'b00000000000011011011110111;
    W_hr[13][1] = 26'b00000000000001110010011111;
    W_hr[13][2] = 26'b11111111111110101100001111;
    W_hr[13][3] = 26'b00000000000010000010011101;
    W_hr[13][4] = 26'b00000000000110100001001011;
    W_hr[13][5] = 26'b11111111111001111001000010;
    W_hr[13][6] = 26'b00000000000000000110101010;
    W_hr[13][7] = 26'b00000000000100011110110101;
    W_hr[13][8] = 26'b00000000000011011001011001;
    W_hr[13][9] = 26'b00000000000000000101010101;
    W_hr[13][10] = 26'b11111111111000001010001111;
    W_hr[13][11] = 26'b00000000000111000111011000;
    W_hr[13][12] = 26'b00000000000101111110111000;
    W_hr[13][13] = 26'b00000000000010001011011110;
    W_hr[13][14] = 26'b11111111111011010011000011;
    W_hr[13][15] = 26'b00000000001010010111010110;
    W_hr[14][0] = 26'b11111111111111010111010000;
    W_hr[14][1] = 26'b11111111111110110011000110;
    W_hr[14][2] = 26'b00000000000010010001100001;
    W_hr[14][3] = 26'b11111111111100110001010111;
    W_hr[14][4] = 26'b11111111111101001011010001;
    W_hr[14][5] = 26'b11111111111111100111010101;
    W_hr[14][6] = 26'b00000000001011101110000101;
    W_hr[14][7] = 26'b11111111111010001000010011;
    W_hr[14][8] = 26'b11111111111111010111001001;
    W_hr[14][9] = 26'b00000000000110110011100000;
    W_hr[14][10] = 26'b00000000001001111100011011;
    W_hr[14][11] = 26'b11111111111001000001001111;
    W_hr[14][12] = 26'b11111111111101011001011001;
    W_hr[14][13] = 26'b11111111111011001100011001;
    W_hr[14][14] = 26'b11111111111100101110000101;
    W_hr[14][15] = 26'b00000000000100111010101011;
    W_hr[15][0] = 26'b00000000000000001110001111;
    W_hr[15][1] = 26'b00000000000000100110100111;
    W_hr[15][2] = 26'b00000000000000111110011110;
    W_hr[15][3] = 26'b11111111111101011100011110;
    W_hr[15][4] = 26'b00000000000100011000010001;
    W_hr[15][5] = 26'b00000000000100101101011110;
    W_hr[15][6] = 26'b00000000000100101010111010;
    W_hr[15][7] = 26'b11111111111011011000011110;
    W_hr[15][8] = 26'b00000000000011111110000011;
    W_hr[15][9] = 26'b00000000000100011111101001;
    W_hr[15][10] = 26'b11111111111101111101110000;
    W_hr[15][11] = 26'b11111111111101100011011100;
    W_hr[15][12] = 26'b00000000000001111101000010;
    W_hr[15][13] = 26'b00000000000010011111110110;
    W_hr[15][14] = 26'b00000000000101101000010000;
    W_hr[15][15] = 26'b11111111111100001101000111;

    // Initialize W_hz weights
    W_hz[0][0] = 26'b00000000000011011011110111;
    W_hz[0][1] = 26'b00000000000001110010011111;
    W_hz[0][2] = 26'b11111111111110101100001111;
    W_hz[0][3] = 26'b00000000000010000010011101;
    W_hz[0][4] = 26'b00000000000110100001001011;
    W_hz[0][5] = 26'b11111111111001111001000010;
    W_hz[0][6] = 26'b00000000000000000110101010;
    W_hz[0][7] = 26'b00000000000100011110110101;
    W_hz[0][8] = 26'b00000000000011011001011001;
    W_hz[0][9] = 26'b00000000000000000101010101;
    W_hz[0][10] = 26'b11111111111000001010001111;
    W_hz[0][11] = 26'b00000000000111000111011000;
    W_hz[0][12] = 26'b00000000000101111110111000;
    W_hz[0][13] = 26'b00000000000010001011011110;
    W_hz[0][14] = 26'b11111111111011010011000011;
    W_hz[0][15] = 26'b00000000001010010111010110;
    W_hz[1][0] = 26'b11111111111111010111010000;
    W_hz[1][1] = 26'b11111111111110110011000110;
    W_hz[1][2] = 26'b00000000000010010001100001;
    W_hz[1][3] = 26'b11111111111100110001010111;
    W_hz[1][4] = 26'b11111111111101001011010001;
    W_hz[1][5] = 26'b11111111111111100111010101;
    W_hz[1][6] = 26'b00000000001011101110000101;
    W_hz[1][7] = 26'b11111111111010001000010011;
    W_hz[1][8] = 26'b11111111111111010111001001;
    W_hz[1][9] = 26'b00000000000110110011100000;
    W_hz[1][10] = 26'b00000000001001111100011011;
    W_hz[1][11] = 26'b11111111111001000001001111;
    W_hz[1][12] = 26'b11111111111101011001011001;
    W_hz[1][13] = 26'b11111111111011001100011001;
    W_hz[1][14] = 26'b11111111111100101110000101;
    W_hz[1][15] = 26'b00000000000100111010101011;
    W_hz[2][0] = 26'b00000000000000001110001111;
    W_hz[2][1] = 26'b00000000000000100110100111;
    W_hz[2][2] = 26'b00000000000000111110011110;
    W_hz[2][3] = 26'b11111111111101011100011110;
    W_hz[2][4] = 26'b00000000000100011000010001;
    W_hz[2][5] = 26'b00000000000100101101011110;
    W_hz[2][6] = 26'b00000000000100101010111010;
    W_hz[2][7] = 26'b11111111111011011000011110;
    W_hz[2][8] = 26'b00000000000011111110000011;
    W_hz[2][9] = 26'b00000000000100011111101001;
    W_hz[2][10] = 26'b11111111111101111101110000;
    W_hz[2][11] = 26'b11111111111101100011011100;
    W_hz[2][12] = 26'b00000000000001111101000010;
    W_hz[2][13] = 26'b00000000000010011111110110;
    W_hz[2][14] = 26'b00000000000101101000010000;
    W_hz[2][15] = 26'b11111111111100001101000111;
    W_hz[3][0] = 26'b00000000000011011011110111;
    W_hz[3][1] = 26'b00000000000001110010011111;
    W_hz[3][2] = 26'b11111111111110101100001111;
    W_hz[3][3] = 26'b00000000000010000010011101;
    W_hz[3][4] = 26'b00000000000110100001001011;
    W_hz[3][5] = 26'b11111111111001111001000010;
    W_hz[3][6] = 26'b00000000000000000110101010;
    W_hz[3][7] = 26'b00000000000100011110110101;
    W_hz[3][8] = 26'b00000000000011011001011001;
    W_hz[3][9] = 26'b00000000000000000101010101;
    W_hz[3][10] = 26'b11111111111000001010001111;
    W_hz[3][11] = 26'b00000000000111000111011000;
    W_hz[3][12] = 26'b00000000000101111110111000;
    W_hz[3][13] = 26'b00000000000010001011011110;
    W_hz[3][14] = 26'b11111111111011010011000011;
    W_hz[3][15] = 26'b00000000001010010111010110;
    W_hz[4][0] = 26'b11111111111111010111010000;
    W_hz[4][1] = 26'b11111111111110110011000110;
    W_hz[4][2] = 26'b00000000000010010001100001;
    W_hz[4][3] = 26'b11111111111100110001010111;
    W_hz[4][4] = 26'b11111111111101001011010001;
    W_hz[4][5] = 26'b11111111111111100111010101;
    W_hz[4][6] = 26'b00000000001011101110000101;
    W_hz[4][7] = 26'b11111111111010001000010011;
    W_hz[4][8] = 26'b11111111111111010111001001;
    W_hz[4][9] = 26'b00000000000110110011100000;
    W_hz[4][10] = 26'b00000000001001111100011011;
    W_hz[4][11] = 26'b11111111111001000001001111;
    W_hz[4][12] = 26'b11111111111101011001011001;
    W_hz[4][13] = 26'b11111111111011001100011001;
    W_hz[4][14] = 26'b11111111111100101110000101;
    W_hz[4][15] = 26'b00000000000100111010101011;
    W_hz[5][0] = 26'b00000000000000001110001111;
    W_hz[5][1] = 26'b00000000000000100110100111;
    W_hz[5][2] = 26'b00000000000000111110011110;
    W_hz[5][3] = 26'b11111111111101011100011110;
    W_hz[5][4] = 26'b00000000000100011000010001;
    W_hz[5][5] = 26'b00000000000100101101011110;
    W_hz[5][6] = 26'b00000000000100101010111010;
    W_hz[5][7] = 26'b11111111111011011000011110;
    W_hz[5][8] = 26'b00000000000011111110000011;
    W_hz[5][9] = 26'b00000000000100011111101001;
    W_hz[5][10] = 26'b11111111111101111101110000;
    W_hz[5][11] = 26'b11111111111101100011011100;
    W_hz[5][12] = 26'b00000000000001111101000010;
    W_hz[5][13] = 26'b00000000000010011111110110;
    W_hz[5][14] = 26'b00000000000101101000010000;
    W_hz[5][15] = 26'b11111111111100001101000111;
    W_hz[6][0] = 26'b00000000000011011011110111;
    W_hz[6][1] = 26'b00000000000001110010011111;
    W_hz[6][2] = 26'b11111111111110101100001111;
    W_hz[6][3] = 26'b00000000000010000010011101;
    W_hz[6][4] = 26'b00000000000110100001001011;
    W_hz[6][5] = 26'b11111111111001111001000010;
    W_hz[6][6] = 26'b00000000000000000110101010;
    W_hz[6][7] = 26'b00000000000100011110110101;
    W_hz[6][8] = 26'b00000000000011011001011001;
    W_hz[6][9] = 26'b00000000000000000101010101;
    W_hz[6][10] = 26'b11111111111000001010001111;
    W_hz[6][11] = 26'b00000000000111000111011000;
    W_hz[6][12] = 26'b00000000000101111110111000;
    W_hz[6][13] = 26'b00000000000010001011011110;
    W_hz[6][14] = 26'b11111111111011010011000011;
    W_hz[6][15] = 26'b00000000001010010111010110;
    W_hz[7][0] = 26'b11111111111111010111010000;
    W_hz[7][1] = 26'b11111111111110110011000110;
    W_hz[7][2] = 26'b00000000000010010001100001;
    W_hz[7][3] = 26'b11111111111100110001010111;
    W_hz[7][4] = 26'b11111111111101001011010001;
    W_hz[7][5] = 26'b11111111111111100111010101;
    W_hz[7][6] = 26'b00000000001011101110000101;
    W_hz[7][7] = 26'b11111111111010001000010011;
    W_hz[7][8] = 26'b11111111111111010111001001;
    W_hz[7][9] = 26'b00000000000110110011100000;
    W_hz[7][10] = 26'b00000000001001111100011011;
    W_hz[7][11] = 26'b11111111111001000001001111;
    W_hz[7][12] = 26'b11111111111101011001011001;
    W_hz[7][13] = 26'b11111111111011001100011001;
    W_hz[7][14] = 26'b11111111111100101110000101;
    W_hz[7][15] = 26'b00000000000100111010101011;
    W_hz[8][0] = 26'b00000000000000001110001111;
    W_hz[8][1] = 26'b00000000000000100110100111;
    W_hz[8][2] = 26'b00000000000000111110011110;
    W_hz[8][3] = 26'b11111111111101011100011110;
    W_hz[8][4] = 26'b00000000000100011000010001;
    W_hz[8][5] = 26'b00000000000100101101011110;
    W_hz[8][6] = 26'b00000000000100101010111010;
    W_hz[8][7] = 26'b11111111111011011000011110;
    W_hz[8][8] = 26'b00000000000011111110000011;
    W_hz[8][9] = 26'b00000000000100011111101001;
    W_hz[8][10] = 26'b11111111111101111101110000;
    W_hz[8][11] = 26'b11111111111101100011011100;
    W_hz[8][12] = 26'b00000000000001111101000010;
    W_hz[8][13] = 26'b00000000000010011111110110;
    W_hz[8][14] = 26'b00000000000101101000010000;
    W_hz[8][15] = 26'b11111111111100001101000111;
    W_hz[9][0] = 26'b00000000000011011011110111;
    W_hz[9][1] = 26'b00000000000001110010011111;
    W_hz[9][2] = 26'b11111111111110101100001111;
    W_hz[9][3] = 26'b00000000000010000010011101;
    W_hz[9][4] = 26'b00000000000110100001001011;
    W_hz[9][5] = 26'b11111111111001111001000010;
    W_hz[9][6] = 26'b00000000000000000110101010;
    W_hz[9][7] = 26'b00000000000100011110110101;
    W_hz[9][8] = 26'b00000000000011011001011001;
    W_hz[9][9] = 26'b00000000000000000101010101;
    W_hz[9][10] = 26'b11111111111000001010001111;
    W_hz[9][11] = 26'b00000000000111000111011000;
    W_hz[9][12] = 26'b00000000000101111110111000;
    W_hz[9][13] = 26'b00000000000010001011011110;
    W_hz[9][14] = 26'b11111111111011010011000011;
    W_hz[9][15] = 26'b00000000001010010111010110;
    W_hz[10][0] = 26'b11111111111111010111010000;
    W_hz[10][1] = 26'b11111111111110110011000110;
    W_hz[10][2] = 26'b00000000000010010001100001;
    W_hz[10][3] = 26'b11111111111100110001010111;
    W_hz[10][4] = 26'b11111111111101001011010001;
    W_hz[10][5] = 26'b11111111111111100111010101;
    W_hz[10][6] = 26'b00000000001011101110000101;
    W_hz[10][7] = 26'b11111111111010001000010011;
    W_hz[10][8] = 26'b11111111111111010111001001;
    W_hz[10][9] = 26'b00000000000110110011100000;
    W_hz[10][10] = 26'b00000000001001111100011011;
    W_hz[10][11] = 26'b11111111111001000001001111;
    W_hz[10][12] = 26'b11111111111101011001011001;
    W_hz[10][13] = 26'b11111111111011001100011001;
    W_hz[10][14] = 26'b11111111111100101110000101;
    W_hz[10][15] = 26'b00000000000100111010101011;
    W_hz[11][0] = 26'b00000000000000001110001111;
    W_hz[11][1] = 26'b00000000000000100110100111;
    W_hz[11][2] = 26'b00000000000000111110011110;
    W_hz[11][3] = 26'b11111111111101011100011110;
    W_hz[11][4] = 26'b00000000000100011000010001;
    W_hz[11][5] = 26'b00000000000100101101011110;
    W_hz[11][6] = 26'b00000000000100101010111010;
    W_hz[11][7] = 26'b11111111111011011000011110;
    W_hz[11][8] = 26'b00000000000011111110000011;
    W_hz[11][9] = 26'b00000000000100011111101001;
    W_hz[11][10] = 26'b11111111111101111101110000;
    W_hz[11][11] = 26'b11111111111101100011011100;
    W_hz[11][12] = 26'b00000000000001111101000010;
    W_hz[11][13] = 26'b00000000000010011111110110;
    W_hz[11][14] = 26'b00000000000101101000010000;
    W_hz[11][15] = 26'b11111111111100001101000111;
    W_hz[12][0] = 26'b00000000000011011011110111;
    W_hz[12][1] = 26'b00000000000001110010011111;
    W_hz[12][2] = 26'b11111111111110101100001111;
    W_hz[12][3] = 26'b00000000000010000010011101;
    W_hz[12][4] = 26'b00000000000110100001001011;
    W_hz[12][5] = 26'b11111111111001111001000010;
    W_hz[12][6] = 26'b00000000000000000110101010;
    W_hz[12][7] = 26'b00000000000100011110110101;
    W_hz[12][8] = 26'b00000000000011011001011001;
    W_hz[12][9] = 26'b00000000000000000101010101;
    W_hz[12][10] = 26'b11111111111000001010001111;
    W_hz[12][11] = 26'b00000000000111000111011000;
    W_hz[12][12] = 26'b00000000000101111110111000;
    W_hz[12][13] = 26'b00000000000010001011011110;
    W_hz[12][14] = 26'b11111111111011010011000011;
    W_hz[12][15] = 26'b00000000001010010111010110;
    W_hz[13][0] = 26'b11111111111111010111010000;
    W_hz[13][1] = 26'b11111111111110110011000110;
    W_hz[13][2] = 26'b00000000000010010001100001;
    W_hz[13][3] = 26'b11111111111100110001010111;
    W_hz[13][4] = 26'b11111111111101001011010001;
    W_hz[13][5] = 26'b11111111111111100111010101;
    W_hz[13][6] = 26'b00000000001011101110000101;
    W_hz[13][7] = 26'b11111111111010001000010011;
    W_hz[13][8] = 26'b11111111111111010111001001;
    W_hz[13][9] = 26'b00000000000110110011100000;
    W_hz[13][10] = 26'b00000000001001111100011011;
    W_hz[13][11] = 26'b11111111111001000001001111;
    W_hz[13][12] = 26'b11111111111101011001011001;
    W_hz[13][13] = 26'b11111111111011001100011001;
    W_hz[13][14] = 26'b11111111111100101110000101;
    W_hz[13][15] = 26'b00000000000100111010101011;
    W_hz[14][0] = 26'b00000000000000001110001111;
    W_hz[14][1] = 26'b00000000000000100110100111;
    W_hz[14][2] = 26'b00000000000000111110011110;
    W_hz[14][3] = 26'b11111111111101011100011110;
    W_hz[14][4] = 26'b00000000000100011000010001;
    W_hz[14][5] = 26'b00000000000100101101011110;
    W_hz[14][6] = 26'b00000000000100101010111010;
    W_hz[14][7] = 26'b11111111111011011000011110;
    W_hz[14][8] = 26'b00000000000011111110000011;
    W_hz[14][9] = 26'b00000000000100011111101001;
    W_hz[14][10] = 26'b11111111111101111101110000;
    W_hz[14][11] = 26'b11111111111101100011011100;
    W_hz[14][12] = 26'b00000000000001111101000010;
    W_hz[14][13] = 26'b00000000000010011111110110;
    W_hz[14][14] = 26'b00000000000101101000010000;
    W_hz[14][15] = 26'b11111111111100001101000111;
    W_hz[15][0] = 26'b00000000000011011011110111;
    W_hz[15][1] = 26'b00000000000001110010011111;
    W_hz[15][2] = 26'b11111111111110101100001111;
    W_hz[15][3] = 26'b00000000000010000010011101;
    W_hz[15][4] = 26'b00000000000110100001001011;
    W_hz[15][5] = 26'b11111111111001111001000010;
    W_hz[15][6] = 26'b00000000000000000110101010;
    W_hz[15][7] = 26'b00000000000100011110110101;
    W_hz[15][8] = 26'b00000000000011011001011001;
    W_hz[15][9] = 26'b00000000000000000101010101;
    W_hz[15][10] = 26'b11111111111000001010001111;
    W_hz[15][11] = 26'b00000000000111000111011000;
    W_hz[15][12] = 26'b00000000000101111110111000;
    W_hz[15][13] = 26'b00000000000010001011011110;
    W_hz[15][14] = 26'b11111111111011010011000011;
    W_hz[15][15] = 26'b00000000001010010111010110;

    // Initialize W_hn weights
    W_hn[0][0] = 26'b11111111111111010111010000;
    W_hn[0][1] = 26'b11111111111110110011000110;
    W_hn[0][2] = 26'b00000000000010010001100001;
    W_hn[0][3] = 26'b11111111111100110001010111;
    W_hn[0][4] = 26'b11111111111101001011010001;
    W_hn[0][5] = 26'b11111111111111100111010101;
    W_hn[0][6] = 26'b00000000001011101110000101;
    W_hn[0][7] = 26'b11111111111010001000010011;
    W_hn[0][8] = 26'b11111111111111010111001001;
    W_hn[0][9] = 26'b00000000000110110011100000;
    W_hn[0][10] = 26'b00000000001001111100011011;
    W_hn[0][11] = 26'b11111111111001000001001111;
    W_hn[0][12] = 26'b11111111111101011001011001;
    W_hn[0][13] = 26'b11111111111011001100011001;
    W_hn[0][14] = 26'b11111111111100101110000101;
    W_hn[0][15] = 26'b00000000000100111010101011;
    W_hn[1][0] = 26'b00000000000000001110001111;
    W_hn[1][1] = 26'b00000000000000100110100111;
    W_hn[1][2] = 26'b00000000000000111110011110;
    W_hn[1][3] = 26'b11111111111101011100011110;
    W_hn[1][4] = 26'b00000000000100011000010001;
    W_hn[1][5] = 26'b00000000000100101101011110;
    W_hn[1][6] = 26'b00000000000100101010111010;
    W_hn[1][7] = 26'b11111111111011011000011110;
    W_hn[1][8] = 26'b00000000000011111110000011;
    W_hn[1][9] = 26'b00000000000100011111101001;
    W_hn[1][10] = 26'b11111111111101111101110000;
    W_hn[1][11] = 26'b11111111111101100011011100;
    W_hn[1][12] = 26'b00000000000001111101000010;
    W_hn[1][13] = 26'b00000000000010011111110110;
    W_hn[1][14] = 26'b00000000000101101000010000;
    W_hn[1][15] = 26'b11111111111100001101000111;
    W_hn[2][0] = 26'b00000000000011011011110111;
    W_hn[2][1] = 26'b00000000000001110010011111;
    W_hn[2][2] = 26'b11111111111110101100001111;
    W_hn[2][3] = 26'b00000000000010000010011101;
    W_hn[2][4] = 26'b00000000000110100001001011;
    W_hn[2][5] = 26'b11111111111001111001000010;
    W_hn[2][6] = 26'b00000000000000000110101010;
    W_hn[2][7] = 26'b00000000000100011110110101;
    W_hn[2][8] = 26'b00000000000011011001011001;
    W_hn[2][9] = 26'b00000000000000000101010101;
    W_hn[2][10] = 26'b11111111111000001010001111;
    W_hn[2][11] = 26'b00000000000111000111011000;
    W_hn[2][12] = 26'b00000000000101111110111000;
    W_hn[2][13] = 26'b00000000000010001011011110;
    W_hn[2][14] = 26'b11111111111011010011000011;
    W_hn[2][15] = 26'b00000000001010010111010110;
    W_hn[3][0] = 26'b11111111111111010111010000;
    W_hn[3][1] = 26'b11111111111110110011000110;
    W_hn[3][2] = 26'b00000000000010010001100001;
    W_hn[3][3] = 26'b11111111111100110001010111;
    W_hn[3][4] = 26'b11111111111101001011010001;
    W_hn[3][5] = 26'b11111111111111100111010101;
    W_hn[3][6] = 26'b00000000001011101110000101;
    W_hn[3][7] = 26'b11111111111010001000010011;
    W_hn[3][8] = 26'b11111111111111010111001001;
    W_hn[3][9] = 26'b00000000000110110011100000;
    W_hn[3][10] = 26'b00000000001001111100011011;
    W_hn[3][11] = 26'b11111111111001000001001111;
    W_hn[3][12] = 26'b11111111111101011001011001;
    W_hn[3][13] = 26'b11111111111011001100011001;
    W_hn[3][14] = 26'b11111111111100101110000101;
    W_hn[3][15] = 26'b00000000000100111010101011;
    W_hn[4][0] = 26'b00000000000000001110001111;
    W_hn[4][1] = 26'b00000000000000100110100111;
    W_hn[4][2] = 26'b00000000000000111110011110;
    W_hn[4][3] = 26'b11111111111101011100011110;
    W_hn[4][4] = 26'b00000000000100011000010001;
    W_hn[4][5] = 26'b00000000000100101101011110;
    W_hn[4][6] = 26'b00000000000100101010111010;
    W_hn[4][7] = 26'b11111111111011011000011110;
    W_hn[4][8] = 26'b00000000000011111110000011;
    W_hn[4][9] = 26'b00000000000100011111101001;
    W_hn[4][10] = 26'b11111111111101111101110000;
    W_hn[4][11] = 26'b11111111111101100011011100;
    W_hn[4][12] = 26'b00000000000001111101000010;
    W_hn[4][13] = 26'b00000000000010011111110110;
    W_hn[4][14] = 26'b00000000000101101000010000;
    W_hn[4][15] = 26'b11111111111100001101000111;
    W_hn[5][0] = 26'b00000000000011011011110111;
    W_hn[5][1] = 26'b00000000000001110010011111;
    W_hn[5][2] = 26'b11111111111110101100001111;
    W_hn[5][3] = 26'b00000000000010000010011101;
    W_hn[5][4] = 26'b00000000000110100001001011;
    W_hn[5][5] = 26'b11111111111001111001000010;
    W_hn[5][6] = 26'b00000000000000000110101010;
    W_hn[5][7] = 26'b00000000000100011110110101;
    W_hn[5][8] = 26'b00000000000011011001011001;
    W_hn[5][9] = 26'b00000000000000000101010101;
    W_hn[5][10] = 26'b11111111111000001010001111;
    W_hn[5][11] = 26'b00000000000111000111011000;
    W_hn[5][12] = 26'b00000000000101111110111000;
    W_hn[5][13] = 26'b00000000000010001011011110;
    W_hn[5][14] = 26'b11111111111011010011000011;
    W_hn[5][15] = 26'b00000000001010010111010110;
    W_hn[6][0] = 26'b11111111111111010111010000;
    W_hn[6][1] = 26'b11111111111110110011000110;
    W_hn[6][2] = 26'b00000000000010010001100001;
    W_hn[6][3] = 26'b11111111111100110001010111;
    W_hn[6][4] = 26'b11111111111101001011010001;
    W_hn[6][5] = 26'b11111111111111100111010101;
    W_hn[6][6] = 26'b00000000001011101110000101;
    W_hn[6][7] = 26'b11111111111010001000010011;
    W_hn[6][8] = 26'b11111111111111010111001001;
    W_hn[6][9] = 26'b00000000000110110011100000;
    W_hn[6][10] = 26'b00000000001001111100011011;
    W_hn[6][11] = 26'b11111111111001000001001111;
    W_hn[6][12] = 26'b11111111111101011001011001;
    W_hn[6][13] = 26'b11111111111011001100011001;
    W_hn[6][14] = 26'b11111111111100101110000101;
    W_hn[6][15] = 26'b00000000000100111010101011;
    W_hn[7][0] = 26'b00000000000000001110001111;
    W_hn[7][1] = 26'b00000000000000100110100111;
    W_hn[7][2] = 26'b00000000000000111110011110;
    W_hn[7][3] = 26'b11111111111101011100011110;
    W_hn[7][4] = 26'b00000000000100011000010001;
    W_hn[7][5] = 26'b00000000000100101101011110;
    W_hn[7][6] = 26'b00000000000100101010111010;
    W_hn[7][7] = 26'b11111111111011011000011110;
    W_hn[7][8] = 26'b00000000000011111110000011;
    W_hn[7][9] = 26'b00000000000100011111101001;
    W_hn[7][10] = 26'b11111111111101111101110000;
    W_hn[7][11] = 26'b11111111111101100011011100;
    W_hn[7][12] = 26'b00000000000001111101000010;
    W_hn[7][13] = 26'b00000000000010011111110110;
    W_hn[7][14] = 26'b00000000000101101000010000;
    W_hn[7][15] = 26'b11111111111100001101000111;
    W_hn[8][0] = 26'b00000000000011011011110111;
    W_hn[8][1] = 26'b00000000000001110010011111;
    W_hn[8][2] = 26'b11111111111110101100001111;
    W_hn[8][3] = 26'b00000000000010000010011101;
    W_hn[8][4] = 26'b00000000000110100001001011;
    W_hn[8][5] = 26'b11111111111001111001000010;
    W_hn[8][6] = 26'b00000000000000000110101010;
    W_hn[8][7] = 26'b00000000000100011110110101;
    W_hn[8][8] = 26'b00000000000011011001011001;
    W_hn[8][9] = 26'b00000000000000000101010101;
    W_hn[8][10] = 26'b11111111111000001010001111;
    W_hn[8][11] = 26'b00000000000111000111011000;
    W_hn[8][12] = 26'b00000000000101111110111000;
    W_hn[8][13] = 26'b00000000000010001011011110;
    W_hn[8][14] = 26'b11111111111011010011000011;
    W_hn[8][15] = 26'b00000000001010010111010110;
    W_hn[9][0] = 26'b11111111111111010111010000;
    W_hn[9][1] = 26'b11111111111110110011000110;
    W_hn[9][2] = 26'b00000000000010010001100001;
    W_hn[9][3] = 26'b11111111111100110001010111;
    W_hn[9][4] = 26'b11111111111101001011010001;
    W_hn[9][5] = 26'b11111111111111100111010101;
    W_hn[9][6] = 26'b00000000001011101110000101;
    W_hn[9][7] = 26'b11111111111010001000010011;
    W_hn[9][8] = 26'b11111111111111010111001001;
    W_hn[9][9] = 26'b00000000000110110011100000;
    W_hn[9][10] = 26'b00000000001001111100011011;
    W_hn[9][11] = 26'b11111111111001000001001111;
    W_hn[9][12] = 26'b11111111111101011001011001;
    W_hn[9][13] = 26'b11111111111011001100011001;
    W_hn[9][14] = 26'b11111111111100101110000101;
    W_hn[9][15] = 26'b00000000000100111010101011;
    W_hn[10][0] = 26'b00000000000000001110001111;
    W_hn[10][1] = 26'b00000000000000100110100111;
    W_hn[10][2] = 26'b00000000000000111110011110;
    W_hn[10][3] = 26'b11111111111101011100011110;
    W_hn[10][4] = 26'b00000000000100011000010001;
    W_hn[10][5] = 26'b00000000000100101101011110;
    W_hn[10][6] = 26'b00000000000100101010111010;
    W_hn[10][7] = 26'b11111111111011011000011110;
    W_hn[10][8] = 26'b00000000000011111110000011;
    W_hn[10][9] = 26'b00000000000100011111101001;
    W_hn[10][10] = 26'b11111111111101111101110000;
    W_hn[10][11] = 26'b11111111111101100011011100;
    W_hn[10][12] = 26'b00000000000001111101000010;
    W_hn[10][13] = 26'b00000000000010011111110110;
    W_hn[10][14] = 26'b00000000000101101000010000;
    W_hn[10][15] = 26'b11111111111100001101000111;
    W_hn[11][0] = 26'b00000000000011011011110111;
    W_hn[11][1] = 26'b00000000000001110010011111;
    W_hn[11][2] = 26'b11111111111110101100001111;
    W_hn[11][3] = 26'b00000000000010000010011101;
    W_hn[11][4] = 26'b00000000000110100001001011;
    W_hn[11][5] = 26'b11111111111001111001000010;
    W_hn[11][6] = 26'b00000000000000000110101010;
    W_hn[11][7] = 26'b00000000000100011110110101;
    W_hn[11][8] = 26'b00000000000011011001011001;
    W_hn[11][9] = 26'b00000000000000000101010101;
    W_hn[11][10] = 26'b11111111111000001010001111;
    W_hn[11][11] = 26'b00000000000111000111011000;
    W_hn[11][12] = 26'b00000000000101111110111000;
    W_hn[11][13] = 26'b00000000000010001011011110;
    W_hn[11][14] = 26'b11111111111011010011000011;
    W_hn[11][15] = 26'b00000000001010010111010110;
    W_hn[12][0] = 26'b11111111111111010111010000;
    W_hn[12][1] = 26'b11111111111110110011000110;
    W_hn[12][2] = 26'b00000000000010010001100001;
    W_hn[12][3] = 26'b11111111111100110001010111;
    W_hn[12][4] = 26'b11111111111101001011010001;
    W_hn[12][5] = 26'b11111111111111100111010101;
    W_hn[12][6] = 26'b00000000001011101110000101;
    W_hn[12][7] = 26'b11111111111010001000010011;
    W_hn[12][8] = 26'b11111111111111010111001001;
    W_hn[12][9] = 26'b00000000000110110011100000;
    W_hn[12][10] = 26'b00000000001001111100011011;
    W_hn[12][11] = 26'b11111111111001000001001111;
    W_hn[12][12] = 26'b11111111111101011001011001;
    W_hn[12][13] = 26'b11111111111011001100011001;
    W_hn[12][14] = 26'b11111111111100101110000101;
    W_hn[12][15] = 26'b00000000000100111010101011;
    W_hn[13][0] = 26'b00000000000000001110001111;
    W_hn[13][1] = 26'b00000000000000100110100111;
    W_hn[13][2] = 26'b00000000000000111110011110;
    W_hn[13][3] = 26'b11111111111101011100011110;
    W_hn[13][4] = 26'b00000000000100011000010001;
    W_hn[13][5] = 26'b00000000000100101101011110;
    W_hn[13][6] = 26'b00000000000100101010111010;
    W_hn[13][7] = 26'b11111111111011011000011110;
    W_hn[13][8] = 26'b00000000000011111110000011;
    W_hn[13][9] = 26'b00000000000100011111101001;
    W_hn[13][10] = 26'b11111111111101111101110000;
    W_hn[13][11] = 26'b11111111111101100011011100;
    W_hn[13][12] = 26'b00000000000001111101000010;
    W_hn[13][13] = 26'b00000000000010011111110110;
    W_hn[13][14] = 26'b00000000000101101000010000;
    W_hn[13][15] = 26'b11111111111100001101000111;
    W_hn[14][0] = 26'b00000000000011011011110111;
    W_hn[14][1] = 26'b00000000000001110010011111;
    W_hn[14][2] = 26'b11111111111110101100001111;
    W_hn[14][3] = 26'b00000000000010000010011101;
    W_hn[14][4] = 26'b00000000000110100001001011;
    W_hn[14][5] = 26'b11111111111001111001000010;
    W_hn[14][6] = 26'b00000000000000000110101010;
    W_hn[14][7] = 26'b00000000000100011110110101;
    W_hn[14][8] = 26'b00000000000011011001011001;
    W_hn[14][9] = 26'b00000000000000000101010101;
    W_hn[14][10] = 26'b11111111111000001010001111;
    W_hn[14][11] = 26'b00000000000111000111011000;
    W_hn[14][12] = 26'b00000000000101111110111000;
    W_hn[14][13] = 26'b00000000000010001011011110;
    W_hn[14][14] = 26'b11111111111011010011000011;
    W_hn[14][15] = 26'b00000000001010010111010110;
    W_hn[15][0] = 26'b11111111111111010111010000;
    W_hn[15][1] = 26'b11111111111110110011000110;
    W_hn[15][2] = 26'b00000000000010010001100001;
    W_hn[15][3] = 26'b11111111111100110001010111;
    W_hn[15][4] = 26'b11111111111101001011010001;
    W_hn[15][5] = 26'b11111111111111100111010101;
    W_hn[15][6] = 26'b00000000001011101110000101;
    W_hn[15][7] = 26'b11111111111010001000010011;
    W_hn[15][8] = 26'b11111111111111010111001001;
    W_hn[15][9] = 26'b00000000000110110011100000;
    W_hn[15][10] = 26'b00000000001001111100011011;
    W_hn[15][11] = 26'b11111111111001000001001111;
    W_hn[15][12] = 26'b11111111111101011001011001;
    W_hn[15][13] = 26'b11111111111011001100011001;
    W_hn[15][14] = 26'b11111111111100101110000101;
    W_hn[15][15] = 26'b00000000000100111010101011;

    // Initialize biases

    // Initialize b_ir biases
    b_ir[0] = 26'b00000000000000010111000011;
    b_ir[1] = 26'b00000000000100001010110000;
    b_ir[2] = 26'b00000000000111011011000010;
    b_ir[3] = 26'b00000000000010100011010101;
    b_ir[4] = 26'b00000000000011000010010111;
    b_ir[5] = 26'b00000000000010001001011011;
    b_ir[6] = 26'b00000000000111111000100010;
    b_ir[7] = 26'b11111111111111110100000001;
    b_ir[8] = 26'b00000000000101010100001011;
    b_ir[9] = 26'b00000000000000111010000100;
    b_ir[10] = 26'b00000000000111000010000011;
    b_ir[11] = 26'b00000000000001001100001100;
    b_ir[12] = 26'b00000000000001001001001110;
    b_ir[13] = 26'b00000000000100111000110101;
    b_ir[14] = 26'b00000000000011011100000100;
    b_ir[15] = 26'b00000000000110100011001110;

    // Initialize b_iz biases
    b_iz[0] = 26'b00000000000011010001000110;
    b_iz[1] = 26'b00000000000100100100110001;
    b_iz[2] = 26'b00000000000010011111101001;
    b_iz[3] = 26'b00000000001100111011001100;
    b_iz[4] = 26'b00000000000001100001001011;
    b_iz[5] = 26'b00000000001001011111100011;
    b_iz[6] = 26'b00000000000011101001111111;
    b_iz[7] = 26'b11111111111000010000100110;
    b_iz[8] = 26'b00000000000000010111000011;
    b_iz[9] = 26'b00000000000100001010110000;
    b_iz[10] = 26'b00000000000111011011000010;
    b_iz[11] = 26'b00000000000010100011010101;
    b_iz[12] = 26'b00000000000011000010010111;
    b_iz[13] = 26'b00000000000010001001011011;
    b_iz[14] = 26'b00000000000111111000100010;
    b_iz[15] = 26'b11111111111111110100000001;

    // Initialize b_in biases
    b_in[0] = 26'b00000000000101010100001011;
    b_in[1] = 26'b00000000000000111010000100;
    b_in[2] = 26'b00000000000111000010000011;
    b_in[3] = 26'b00000000000001001100001100;
    b_in[4] = 26'b00000000000001001001001110;
    b_in[5] = 26'b00000000000100111000110101;
    b_in[6] = 26'b00000000000011011100000100;
    b_in[7] = 26'b00000000000110100011001110;
    b_in[8] = 26'b00000000000011010001000110;
    b_in[9] = 26'b00000000000100100100110001;
    b_in[10] = 26'b00000000000010011111101001;
    b_in[11] = 26'b00000000001100111011001100;
    b_in[12] = 26'b00000000000001100001001011;
    b_in[13] = 26'b00000000001001011111100011;
    b_in[14] = 26'b00000000000011101001111111;
    b_in[15] = 26'b11111111111000010000100110;

    // Initialize b_hr biases
    b_hr[0] = 26'b00000000000000010111000011;
    b_hr[1] = 26'b00000000000100001010110000;
    b_hr[2] = 26'b00000000000111011011000010;
    b_hr[3] = 26'b00000000000010100011010101;
    b_hr[4] = 26'b00000000000011000010010111;
    b_hr[5] = 26'b00000000000010001001011011;
    b_hr[6] = 26'b00000000000111111000100010;
    b_hr[7] = 26'b11111111111111110100000001;
    b_hr[8] = 26'b00000000000101010100001011;
    b_hr[9] = 26'b00000000000000111010000100;
    b_hr[10] = 26'b00000000000111000010000011;
    b_hr[11] = 26'b00000000000001001100001100;
    b_hr[12] = 26'b00000000000001001001001110;
    b_hr[13] = 26'b00000000000100111000110101;
    b_hr[14] = 26'b00000000000011011100000100;
    b_hr[15] = 26'b00000000000110100011001110;

    // Initialize b_hz biases
    b_hz[0] = 26'b00000000000011010001000110;
    b_hz[1] = 26'b00000000000100100100110001;
    b_hz[2] = 26'b00000000000010011111101001;
    b_hz[3] = 26'b00000000001100111011001100;
    b_hz[4] = 26'b00000000000001100001001011;
    b_hz[5] = 26'b00000000001001011111100011;
    b_hz[6] = 26'b00000000000011101001111111;
    b_hz[7] = 26'b11111111111000010000100110;
    b_hz[8] = 26'b00000000000000010111000011;
    b_hz[9] = 26'b00000000000100001010110000;
    b_hz[10] = 26'b00000000000111011011000010;
    b_hz[11] = 26'b00000000000010100011010101;
    b_hz[12] = 26'b00000000000011000010010111;
    b_hz[13] = 26'b00000000000010001001011011;
    b_hz[14] = 26'b00000000000111111000100010;
    b_hz[15] = 26'b11111111111111110100000001;

    // Initialize b_hn biases
    b_hn[0] = 26'b00000000000101010100001011;
    b_hn[1] = 26'b00000000000000111010000100;
    b_hn[2] = 26'b00000000000111000010000011;
    b_hn[3] = 26'b00000000000001001100001100;
    b_hn[4] = 26'b00000000000001001001001110;
    b_hn[5] = 26'b00000000000100111000110101;
    b_hn[6] = 26'b00000000000011011100000100;
    b_hn[7] = 26'b00000000000110100011001110;
    b_hn[8] = 26'b00000000000011010001000110;
    b_hn[9] = 26'b00000000000100100100110001;
    b_hn[10] = 26'b00000000000010011111101001;
    b_hn[11] = 26'b00000000001100111011001100;
    b_hn[12] = 26'b00000000000001100001001011;
    b_hn[13] = 26'b00000000001001011111100011;
    b_hn[14] = 26'b00000000000011101001111111;
    b_hn[15] = 26'b11111111111000010000100110;

    // Reset sequence
    rst_n = 0;
    start = 0;
    test_start_cycle = 0;
    test_cycles = 0;
    total_cycles = 0;
    test_timeout = 0;
    repeat(10) @(posedge clk);
    rst_n = 1;
    repeat(5) @(posedge clk);

    // Test Vector 1
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000010010001001001110;
        x_t[1] = 26'b00000000011011011000100100;
        x_t[2] = 26'b00000000100000100100110110;
        x_t[3] = 26'b00000000100100011001110110;
        x_t[4] = 26'b00000000011101010011011111;
        x_t[5] = 26'b00000000011010111000010001;
        x_t[6] = 26'b00000000010011101000101111;
        x_t[7] = 26'b00000000010010011111000010;
        x_t[8] = 26'b00000000011110000101000011;
        x_t[9] = 26'b00000000100100001000011111;
        x_t[10] = 26'b00000000100101101001011010;
        x_t[11] = 26'b00000000100100100100101101;
        x_t[12] = 26'b00000000100011101100000011;
        x_t[13] = 26'b00000000010110010001101000;
        x_t[14] = 26'b00000000011101010111011101;
        x_t[15] = 26'b00000000100011001000001010;
        x_t[16] = 26'b00000000100100111101001010;
        x_t[17] = 26'b00000000100110011111001111;
        x_t[18] = 26'b00000000100111101101100110;
        x_t[19] = 26'b00000000100110110001000110;
        x_t[20] = 26'b00000000011011011111000010;
        x_t[21] = 26'b00000000001000010001110100;
        x_t[22] = 26'b00000000001001111010110111;
        x_t[23] = 26'b00000000001011101110010101;
        x_t[24] = 26'b00000000000101110100111101;
        x_t[25] = 26'b00000000000111001100111111;
        x_t[26] = 26'b00000000010100010010101110;
        x_t[27] = 26'b00000000001101110110110111;
        x_t[28] = 26'b00000000001110111110101111;
        x_t[29] = 26'b00000000000101110001000100;
        x_t[30] = 26'b00000000001011110100010001;
        x_t[31] = 26'b00000000011000111010001000;
        x_t[32] = 26'b00000000011110110100110100;
        x_t[33] = 26'b00000000011111000001100111;
        x_t[34] = 26'b00000000011011111001001110;
        x_t[35] = 26'b00000000010111101000001001;
        x_t[36] = 26'b00000000010011110010101101;
        x_t[37] = 26'b00000000001010001111110101;
        x_t[38] = 26'b00000000001011100111100100;
        x_t[39] = 26'b00000000010001110011011011;
        x_t[40] = 26'b00000000010101001111101101;
        x_t[41] = 26'b00000000011010001100110111;
        x_t[42] = 26'b00000000010000001101000011;
        x_t[43] = 26'b00000000001101011111110010;
        x_t[44] = 26'b00000000011000010101001100;
        x_t[45] = 26'b00000000001011100101000010;
        x_t[46] = 26'b00000000011101010000110001;
        x_t[47] = 26'b00000000100001010111110000;
        x_t[48] = 26'b00000000011111101111011101;
        x_t[49] = 26'b00000000100010110001000111;
        x_t[50] = 26'b00000000101000100101100111;
        x_t[51] = 26'b00000000101010101101001100;
        x_t[52] = 26'b00000000101000011011100111;
        x_t[53] = 26'b00000000100011000010110101;
        x_t[54] = 26'b00000000011011010010000110;
        x_t[55] = 26'b00000000011011010101111111;
        x_t[56] = 26'b00000000100001010111111000;
        x_t[57] = 26'b00000000100011000010000100;
        x_t[58] = 26'b00000000100100011111010011;
        x_t[59] = 26'b00000000010111011000111101;
        x_t[60] = 26'b00000000010111111010000011;
        x_t[61] = 26'b00000000011001100100010100;
        x_t[62] = 26'b00000000010010101100000010;
        x_t[63] = 26'b00000000010111111100100001;
        
        h_t_prev[0] = 26'b00000000010010001001001110;
        h_t_prev[1] = 26'b00000000011011011000100100;
        h_t_prev[2] = 26'b00000000100000100100110110;
        h_t_prev[3] = 26'b00000000100100011001110110;
        h_t_prev[4] = 26'b00000000011101010011011111;
        h_t_prev[5] = 26'b00000000011010111000010001;
        h_t_prev[6] = 26'b00000000010011101000101111;
        h_t_prev[7] = 26'b00000000010010011111000010;
        h_t_prev[8] = 26'b00000000011110000101000011;
        h_t_prev[9] = 26'b00000000100100001000011111;
        h_t_prev[10] = 26'b00000000100101101001011010;
        h_t_prev[11] = 26'b00000000100100100100101101;
        h_t_prev[12] = 26'b00000000100011101100000011;
        h_t_prev[13] = 26'b00000000010110010001101000;
        h_t_prev[14] = 26'b00000000011101010111011101;
        h_t_prev[15] = 26'b00000000100011001000001010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 1 timeout!");
                $fdisplay(fd_cycles, "Test Vector   1: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   1: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 1");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 2
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000010111000100111011;
        x_t[1] = 26'b00000000100100100011111001;
        x_t[2] = 26'b00000000101000110001010001;
        x_t[3] = 26'b00000000101010101111111010;
        x_t[4] = 26'b00000000100111101110010111;
        x_t[5] = 26'b00000000100101111110010010;
        x_t[6] = 26'b00000000011111101100011101;
        x_t[7] = 26'b00000000011011011001000101;
        x_t[8] = 26'b00000000101000101101110011;
        x_t[9] = 26'b00000000101100111001101111;
        x_t[10] = 26'b00000000101101010010101010;
        x_t[11] = 26'b00000000101111011001110000;
        x_t[12] = 26'b00000000101101001100110010;
        x_t[13] = 26'b00000000100000000100100010;
        x_t[14] = 26'b00000000100110100110000110;
        x_t[15] = 26'b00000000101011011001000010;
        x_t[16] = 26'b00000000101100000101001011;
        x_t[17] = 26'b00000000101110100000011110;
        x_t[18] = 26'b00000000101110111101011100;
        x_t[19] = 26'b00000000101110010100011000;
        x_t[20] = 26'b00000000100001101111011110;
        x_t[21] = 26'b00000000001001010100000111;
        x_t[22] = 26'b00000000001001111010110111;
        x_t[23] = 26'b00000000001011001011100010;
        x_t[24] = 26'b00000000001100000110110111;
        x_t[25] = 26'b00000000001100110101100000;
        x_t[26] = 26'b00000000010110011001111001;
        x_t[27] = 26'b00000000010000100011110011;
        x_t[28] = 26'b00000000001101001101011000;
        x_t[29] = 26'b00000000010001011101110010;
        x_t[30] = 26'b00000000010100110101110111;
        x_t[31] = 26'b00000000011100001111000010;
        x_t[32] = 26'b00000000100001000110001100;
        x_t[33] = 26'b00000000011111111001001000;
        x_t[34] = 26'b00000000011100110010011000;
        x_t[35] = 26'b00000000011010011001110010;
        x_t[36] = 26'b00000000010100101110010110;
        x_t[37] = 26'b00000000001100100010100110;
        x_t[38] = 26'b00000000011010011011100011;
        x_t[39] = 26'b00000000001010111010011111;
        x_t[40] = 26'b00000000100001001000100100;
        x_t[41] = 26'b11111111111110011000100000;
        x_t[42] = 26'b00000000011101001011001000;
        x_t[43] = 26'b00000000010010010010111111;
        x_t[44] = 26'b00000000100011110110100001;
        x_t[45] = 26'b00000000000010011000111101;
        x_t[46] = 26'b00000000100100011000101010;
        x_t[47] = 26'b00000000100100011110101100;
        x_t[48] = 26'b00000000100000000010100001;
        x_t[49] = 26'b00000000100000011100110110;
        x_t[50] = 26'b00000000100110110011100101;
        x_t[51] = 26'b00000000101000111001010010;
        x_t[52] = 26'b00000000100100100110000100;
        x_t[53] = 26'b00000000011101110100110010;
        x_t[54] = 26'b00000000010100111010100101;
        x_t[55] = 26'b00000000011010010000111011;
        x_t[56] = 26'b00000000011110111101001101;
        x_t[57] = 26'b00000000011111000010010010;
        x_t[58] = 26'b00000000100001001101111100;
        x_t[59] = 26'b00000000010100011011011111;
        x_t[60] = 26'b00000000010111001100000011;
        x_t[61] = 26'b00000000011001110100111000;
        x_t[62] = 26'b00000000010011001001101000;
        x_t[63] = 26'b00000000010110100100100001;
        
        h_t_prev[0] = 26'b00000000010111000100111011;
        h_t_prev[1] = 26'b00000000100100100011111001;
        h_t_prev[2] = 26'b00000000101000110001010001;
        h_t_prev[3] = 26'b00000000101010101111111010;
        h_t_prev[4] = 26'b00000000100111101110010111;
        h_t_prev[5] = 26'b00000000100101111110010010;
        h_t_prev[6] = 26'b00000000011111101100011101;
        h_t_prev[7] = 26'b00000000011011011001000101;
        h_t_prev[8] = 26'b00000000101000101101110011;
        h_t_prev[9] = 26'b00000000101100111001101111;
        h_t_prev[10] = 26'b00000000101101010010101010;
        h_t_prev[11] = 26'b00000000101111011001110000;
        h_t_prev[12] = 26'b00000000101101001100110010;
        h_t_prev[13] = 26'b00000000100000000100100010;
        h_t_prev[14] = 26'b00000000100110100110000110;
        h_t_prev[15] = 26'b00000000101011011001000010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 2 timeout!");
                $fdisplay(fd_cycles, "Test Vector   2: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   2: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 2");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 3
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000011111101101011000;
        x_t[1] = 26'b00000000100001100000000111;
        x_t[2] = 26'b00000000100000010001011011;
        x_t[3] = 26'b00000000011111110111110100;
        x_t[4] = 26'b00000000011011011010001111;
        x_t[5] = 26'b00000000010110010111110100;
        x_t[6] = 26'b00000000001110111110000001;
        x_t[7] = 26'b00000000011000110110001101;
        x_t[8] = 26'b00000000100000111110101101;
        x_t[9] = 26'b00000000100000101100000000;
        x_t[10] = 26'b00000000100000001001001010;
        x_t[11] = 26'b00000000100001101101010000;
        x_t[12] = 26'b00000000011010001011010100;
        x_t[13] = 26'b00000000000110111100010111;
        x_t[14] = 26'b00000000100000010101010011;
        x_t[15] = 26'b00000000100001001110000111;
        x_t[16] = 26'b00000000100000010011101111;
        x_t[17] = 26'b00000000100001100011011001;
        x_t[18] = 26'b00000000100000011101110000;
        x_t[19] = 26'b00000000011101110101111101;
        x_t[20] = 26'b00000000001110100101000111;
        x_t[21] = 26'b00000000010000100100010000;
        x_t[22] = 26'b00000000001100111001010000;
        x_t[23] = 26'b00000000001011101110010101;
        x_t[24] = 26'b00000000010110000000001100;
        x_t[25] = 26'b00000000010110100011000110;
        x_t[26] = 26'b00000000010001111010101001;
        x_t[27] = 26'b00000000001101110110110111;
        x_t[28] = 26'b00000000001011110101001110;
        x_t[29] = 26'b00000000011101101011110001;
        x_t[30] = 26'b00000000010101100100101101;
        x_t[31] = 26'b00000000010100011110001111;
        x_t[32] = 26'b00000000011001101101101110;
        x_t[33] = 26'b00000000010110111011100011;
        x_t[34] = 26'b00000000010011010000101101;
        x_t[35] = 26'b00000000010000110101111010;
        x_t[36] = 26'b00000000001100101001011111;
        x_t[37] = 26'b00000000001001001110100110;
        x_t[38] = 26'b00000000011001110011001101;
        x_t[39] = 26'b00000000000000110011110000;
        x_t[40] = 26'b00000000011100000010011110;
        x_t[41] = 26'b00000000000000100011100110;
        x_t[42] = 26'b00000000011010111100110101;
        x_t[43] = 26'b00000000010000111011001110;
        x_t[44] = 26'b00000000011101111010101100;
        x_t[45] = 26'b00000000000001111010000000;
        x_t[46] = 26'b00000000011100111100000011;
        x_t[47] = 26'b00000000011011011101110011;
        x_t[48] = 26'b00000000010101100111011110;
        x_t[49] = 26'b00000000010110000001101001;
        x_t[50] = 26'b00000000011100000111011001;
        x_t[51] = 26'b00000000011101101110100000;
        x_t[52] = 26'b00000000011001101110010110;
        x_t[53] = 26'b00000000010101011110010100;
        x_t[54] = 26'b00000000010000110010111001;
        x_t[55] = 26'b00000000010010101101100100;
        x_t[56] = 26'b00000000010111111110010110;
        x_t[57] = 26'b00000000010111000010101101;
        x_t[58] = 26'b00000000011010101011001100;
        x_t[59] = 26'b00000000010010101100111110;
        x_t[60] = 26'b00000000010011000111010111;
        x_t[61] = 26'b00000000010111001111010101;
        x_t[62] = 26'b00000000010001000100011110;
        x_t[63] = 26'b00000000010111000111101110;
        
        h_t_prev[0] = 26'b00000000011111101101011000;
        h_t_prev[1] = 26'b00000000100001100000000111;
        h_t_prev[2] = 26'b00000000100000010001011011;
        h_t_prev[3] = 26'b00000000011111110111110100;
        h_t_prev[4] = 26'b00000000011011011010001111;
        h_t_prev[5] = 26'b00000000010110010111110100;
        h_t_prev[6] = 26'b00000000001110111110000001;
        h_t_prev[7] = 26'b00000000011000110110001101;
        h_t_prev[8] = 26'b00000000100000111110101101;
        h_t_prev[9] = 26'b00000000100000101100000000;
        h_t_prev[10] = 26'b00000000100000001001001010;
        h_t_prev[11] = 26'b00000000100001101101010000;
        h_t_prev[12] = 26'b00000000011010001011010100;
        h_t_prev[13] = 26'b00000000000110111100010111;
        h_t_prev[14] = 26'b00000000100000010101010011;
        h_t_prev[15] = 26'b00000000100001001110000111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 3 timeout!");
                $fdisplay(fd_cycles, "Test Vector   3: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   3: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 3");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 4
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000010110011101011101;
        x_t[1] = 26'b00000000010111101101101001;
        x_t[2] = 26'b00000000011010001100111101;
        x_t[3] = 26'b00000000011100110110011100;
        x_t[4] = 26'b00000000011000010000001010;
        x_t[5] = 26'b00000000010010001101100100;
        x_t[6] = 26'b00000000001101110011010101;
        x_t[7] = 26'b00000000001111010011011101;
        x_t[8] = 26'b00000000011000010001101110;
        x_t[9] = 26'b00000000011010101111001010;
        x_t[10] = 26'b00000000011011110111001011;
        x_t[11] = 26'b00000000011101111000101010;
        x_t[12] = 26'b00000000010101011010111101;
        x_t[13] = 26'b00000000001000101001011001;
        x_t[14] = 26'b00000000010111000110101011;
        x_t[15] = 26'b00000000011010110111010010;
        x_t[16] = 26'b00000000011010011011000001;
        x_t[17] = 26'b00000000011011000100110111;
        x_t[18] = 26'b00000000011011100001100000;
        x_t[19] = 26'b00000000011001000010011011;
        x_t[20] = 26'b00000000001101110011000100;
        x_t[21] = 26'b00000000001101101000011001;
        x_t[22] = 26'b00000000001100101100100100;
        x_t[23] = 26'b00000000001111010110010111;
        x_t[24] = 26'b00000000010000000110101001;
        x_t[25] = 26'b00000000010001000111000000;
        x_t[26] = 26'b00000000010011001111001000;
        x_t[27] = 26'b00000000010001000011001111;
        x_t[28] = 26'b00000000010001111011101010;
        x_t[29] = 26'b00000000010000101011110111;
        x_t[30] = 26'b00000000001111101110000011;
        x_t[31] = 26'b00000000010100001100100000;
        x_t[32] = 26'b00000000011000010010110111;
        x_t[33] = 26'b00000000011000000101100011;
        x_t[34] = 26'b00000000010101111100001011;
        x_t[35] = 26'b00000000010010011000100110;
        x_t[36] = 26'b00000000010001100111100100;
        x_t[37] = 26'b00000000001101100011110101;
        x_t[38] = 26'b00000000001110001000111011;
        x_t[39] = 26'b00000000001110001000010000;
        x_t[40] = 26'b00000000011000010011010110;
        x_t[41] = 26'b00000000010110010010100000;
        x_t[42] = 26'b00000000010000100100110001;
        x_t[43] = 26'b00000000000110101000111011;
        x_t[44] = 26'b00000000010000111111111110;
        x_t[45] = 26'b00000000000111101101011011;
        x_t[46] = 26'b00000000010001100110110000;
        x_t[47] = 26'b00000000010100010100010000;
        x_t[48] = 26'b00000000010001011100101001;
        x_t[49] = 26'b00000000010001111110001011;
        x_t[50] = 26'b00000000010110001011010010;
        x_t[51] = 26'b00000000010111000101100000;
        x_t[52] = 26'b00000000010011101001100011;
        x_t[53] = 26'b00000000010001111111101000;
        x_t[54] = 26'b00000000001111101010111110;
        x_t[55] = 26'b00000000001110101010100111;
        x_t[56] = 26'b00000000010011101011010111;
        x_t[57] = 26'b00000000010011100101000010;
        x_t[58] = 26'b00000000010110000010100110;
        x_t[59] = 26'b00000000010000101110101010;
        x_t[60] = 26'b00000000001110100100000000;
        x_t[61] = 26'b00000000010011010111000010;
        x_t[62] = 26'b00000000001101001000111101;
        x_t[63] = 26'b00000000010110110110000111;
        
        h_t_prev[0] = 26'b00000000010110011101011101;
        h_t_prev[1] = 26'b00000000010111101101101001;
        h_t_prev[2] = 26'b00000000011010001100111101;
        h_t_prev[3] = 26'b00000000011100110110011100;
        h_t_prev[4] = 26'b00000000011000010000001010;
        h_t_prev[5] = 26'b00000000010010001101100100;
        h_t_prev[6] = 26'b00000000001101110011010101;
        h_t_prev[7] = 26'b00000000001111010011011101;
        h_t_prev[8] = 26'b00000000011000010001101110;
        h_t_prev[9] = 26'b00000000011010101111001010;
        h_t_prev[10] = 26'b00000000011011110111001011;
        h_t_prev[11] = 26'b00000000011101111000101010;
        h_t_prev[12] = 26'b00000000010101011010111101;
        h_t_prev[13] = 26'b00000000001000101001011001;
        h_t_prev[14] = 26'b00000000010111000110101011;
        h_t_prev[15] = 26'b00000000011010110111010010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 4 timeout!");
                $fdisplay(fd_cycles, "Test Vector   4: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   4: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 4");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 5
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001110001000101110;
        x_t[1] = 26'b00000000010010110100011010;
        x_t[2] = 26'b00000000010100101111010110;
        x_t[3] = 26'b00000000011000100111101111;
        x_t[4] = 26'b00000000010110000010101101;
        x_t[5] = 26'b00000000010000001000011011;
        x_t[6] = 26'b00000000001110100101000111;
        x_t[7] = 26'b00000000001010001101101101;
        x_t[8] = 26'b00000000010000100010100111;
        x_t[9] = 26'b00000000010011100010001000;
        x_t[10] = 26'b00000000010101001000101001;
        x_t[11] = 26'b00000000011000001001110000;
        x_t[12] = 26'b00000000010000010011001011;
        x_t[13] = 26'b00000000000111110010111000;
        x_t[14] = 26'b00000000010001001010111111;
        x_t[15] = 26'b00000000010100001100000111;
        x_t[16] = 26'b00000000010011111010101001;
        x_t[17] = 26'b00000000010011111110110110;
        x_t[18] = 26'b00000000010011100111011111;
        x_t[19] = 26'b00000000010000110011001101;
        x_t[20] = 26'b00000000001001000110101110;
        x_t[21] = 26'b00000000001111010110111010;
        x_t[22] = 26'b00000000001010100000111100;
        x_t[23] = 26'b00000000001101100010010110;
        x_t[24] = 26'b00000000001010110001100111;
        x_t[25] = 26'b00000000001011010010000011;
        x_t[26] = 26'b00000000010000000100010111;
        x_t[27] = 26'b00000000001110100110000010;
        x_t[28] = 26'b00000000001111100100100001;
        x_t[29] = 26'b00000000000111000100010001;
        x_t[30] = 26'b00000000001100100011000111;
        x_t[31] = 26'b00000000010000100101110110;
        x_t[32] = 26'b00000000010011110000000110;
        x_t[33] = 26'b00000000010011001011000000;
        x_t[34] = 26'b00000000010010010111100011;
        x_t[35] = 26'b00000000001101011100110011;
        x_t[36] = 26'b00000000001100111101010111;
        x_t[37] = 26'b00000000001001111111100001;
        x_t[38] = 26'b00000000000101111100100001;
        x_t[39] = 26'b00000000000110110001111010;
        x_t[40] = 26'b00000000000011001111100011;
        x_t[41] = 26'b00000000000110001101001111;
        x_t[42] = 26'b00000000000001110000000111;
        x_t[43] = 26'b11111111111101101110011010;
        x_t[44] = 26'b00000000001000100111101111;
        x_t[45] = 26'b00000000000001111010000000;
        x_t[46] = 26'b00000000001110101100010000;
        x_t[47] = 26'b00000000010010001001000000;
        x_t[48] = 26'b00000000001110011110000011;
        x_t[49] = 26'b00000000001111010111010111;
        x_t[50] = 26'b00000000010010010100001110;
        x_t[51] = 26'b00000000010010100011101110;
        x_t[52] = 26'b00000000001110100010001001;
        x_t[53] = 26'b00000000001101000111110110;
        x_t[54] = 26'b00000000001001101011011011;
        x_t[55] = 26'b00000000001101000011000010;
        x_t[56] = 26'b00000000010001110011000011;
        x_t[57] = 26'b00000000010001101101101010;
        x_t[58] = 26'b00000000010010011111110001;
        x_t[59] = 26'b00000000001100110010000010;
        x_t[60] = 26'b00000000001100001010101010;
        x_t[61] = 26'b00000000010000010000011000;
        x_t[62] = 26'b00000000001001001101011100;
        x_t[63] = 26'b00000000010101001100100000;
        
        h_t_prev[0] = 26'b00000000001110001000101110;
        h_t_prev[1] = 26'b00000000010010110100011010;
        h_t_prev[2] = 26'b00000000010100101111010110;
        h_t_prev[3] = 26'b00000000011000100111101111;
        h_t_prev[4] = 26'b00000000010110000010101101;
        h_t_prev[5] = 26'b00000000010000001000011011;
        h_t_prev[6] = 26'b00000000001110100101000111;
        h_t_prev[7] = 26'b00000000001010001101101101;
        h_t_prev[8] = 26'b00000000010000100010100111;
        h_t_prev[9] = 26'b00000000010011100010001000;
        h_t_prev[10] = 26'b00000000010101001000101001;
        h_t_prev[11] = 26'b00000000011000001001110000;
        h_t_prev[12] = 26'b00000000010000010011001011;
        h_t_prev[13] = 26'b00000000000111110010111000;
        h_t_prev[14] = 26'b00000000010001001010111111;
        h_t_prev[15] = 26'b00000000010100001100000111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 5 timeout!");
                $fdisplay(fd_cycles, "Test Vector   5: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   5: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 5");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 6
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001001100000110000;
        x_t[1] = 26'b00000000001111011101000011;
        x_t[2] = 26'b00000000010010000000100010;
        x_t[3] = 26'b00000000010101111001101110;
        x_t[4] = 26'b00000000010010100100011011;
        x_t[5] = 26'b00000000001011010001110011;
        x_t[6] = 26'b00000000001010010011010010;
        x_t[7] = 26'b00000000000101011100010101;
        x_t[8] = 26'b00000000001110010010001110;
        x_t[9] = 26'b00000000010010100110000000;
        x_t[10] = 26'b00000000010100001101111100;
        x_t[11] = 26'b00000000010111100000111111;
        x_t[12] = 26'b00000000001111001100111100;
        x_t[13] = 26'b00000000000110100001000111;
        x_t[14] = 26'b00000000001111110110100111;
        x_t[15] = 26'b00000000010011100011011011;
        x_t[16] = 26'b00000000010011100110110100;
        x_t[17] = 26'b00000000010100100110010100;
        x_t[18] = 26'b00000000010011010010011010;
        x_t[19] = 26'b00000000010010001011000101;
        x_t[20] = 26'b00000000001010010001110100;
        x_t[21] = 26'b00000000001001101010001110;
        x_t[22] = 26'b00000000001000001000101000;
        x_t[23] = 26'b00000000001001000000010100;
        x_t[24] = 26'b00000000001001000100000000;
        x_t[25] = 26'b00000000001001010101101111;
        x_t[26] = 26'b00000000001100111001100110;
        x_t[27] = 26'b00000000001001101011100110;
        x_t[28] = 26'b00000000001001011110000101;
        x_t[29] = 26'b00000000000110000001101101;
        x_t[30] = 26'b00000000001110101111100110;
        x_t[31] = 26'b00000000001110111011011000;
        x_t[32] = 26'b00000000010011110000000110;
        x_t[33] = 26'b00000000010010010011100000;
        x_t[34] = 26'b00000000010000010010001100;
        x_t[35] = 26'b00000000001100110101010100;
        x_t[36] = 26'b00000000001001110110100101;
        x_t[37] = 26'b00000000000110011011001110;
        x_t[38] = 26'b00000000000101010100001011;
        x_t[39] = 26'b00000000000100011110111011;
        x_t[40] = 26'b00000000001000101011010111;
        x_t[41] = 26'b00000000000010101110101100;
        x_t[42] = 26'b00000000001010101001010011;
        x_t[43] = 26'b00000000001101011111110010;
        x_t[44] = 26'b00000000001100110011110111;
        x_t[45] = 26'b00000000000100110011101101;
        x_t[46] = 26'b00000000001100101111111011;
        x_t[47] = 26'b00000000001110101110001011;
        x_t[48] = 26'b00000000001010100110010011;
        x_t[49] = 26'b00000000001101111010101101;
        x_t[50] = 26'b00000000010010010100001110;
        x_t[51] = 26'b00000000010100010111101001;
        x_t[52] = 26'b00000000010010000011001111;
        x_t[53] = 26'b00000000010010101100001010;
        x_t[54] = 26'b00000000001101011011001001;
        x_t[55] = 26'b00000000001000101110110100;
        x_t[56] = 26'b00000000001101110001010000;
        x_t[57] = 26'b00000000001111100101001111;
        x_t[58] = 26'b00000000010011010100000111;
        x_t[59] = 26'b00000000001100100010001111;
        x_t[60] = 26'b00000000001010000000101001;
        x_t[61] = 26'b00000000001101011010010010;
        x_t[62] = 26'b00000000000101100000101110;
        x_t[63] = 26'b00000000010001010110000100;
        
        h_t_prev[0] = 26'b00000000001001100000110000;
        h_t_prev[1] = 26'b00000000001111011101000011;
        h_t_prev[2] = 26'b00000000010010000000100010;
        h_t_prev[3] = 26'b00000000010101111001101110;
        h_t_prev[4] = 26'b00000000010010100100011011;
        h_t_prev[5] = 26'b00000000001011010001110011;
        h_t_prev[6] = 26'b00000000001010010011010010;
        h_t_prev[7] = 26'b00000000000101011100010101;
        h_t_prev[8] = 26'b00000000001110010010001110;
        h_t_prev[9] = 26'b00000000010010100110000000;
        h_t_prev[10] = 26'b00000000010100001101111100;
        h_t_prev[11] = 26'b00000000010111100000111111;
        h_t_prev[12] = 26'b00000000001111001100111100;
        h_t_prev[13] = 26'b00000000000110100001000111;
        h_t_prev[14] = 26'b00000000001111110110100111;
        h_t_prev[15] = 26'b00000000010011100011011011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 6 timeout!");
                $fdisplay(fd_cycles, "Test Vector   6: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   6: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 6");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 7
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001100010010010101;
        x_t[1] = 26'b00000000010010100000110101;
        x_t[2] = 26'b00000000010101111101000010;
        x_t[3] = 26'b00000000011010011011110000;
        x_t[4] = 26'b00000000010111010011100010;
        x_t[5] = 26'b00000000010001001011000000;
        x_t[6] = 26'b00000000001110001100001110;
        x_t[7] = 26'b00000000000011001101110100;
        x_t[8] = 26'b00000000010000001101111111;
        x_t[9] = 26'b00000000010101011010011001;
        x_t[10] = 26'b00000000011000011111111010;
        x_t[11] = 26'b00000000011101001111111001;
        x_t[12] = 26'b00000000010111010000000001;
        x_t[13] = 26'b00000000001110001011101111;
        x_t[14] = 26'b00000000001001100101110100;
        x_t[15] = 26'b00000000010010010010000100;
        x_t[16] = 26'b00000000010100001110011110;
        x_t[17] = 26'b00000000010101001101110011;
        x_t[18] = 26'b00000000010110111010010101;
        x_t[19] = 26'b00000000011001000010011011;
        x_t[20] = 26'b00000000010100011100100010;
        x_t[21] = 26'b00000000001000010001110100;
        x_t[22] = 26'b00000000000111010101110111;
        x_t[23] = 26'b00000000000111100011100000;
        x_t[24] = 26'b00000000001011001001111110;
        x_t[25] = 26'b00000000001011011110011111;
        x_t[26] = 26'b00000000001110101111111000;
        x_t[27] = 26'b00000000001011001001111011;
        x_t[28] = 26'b00000000001001000100111001;
        x_t[29] = 26'b00000000001000101000000110;
        x_t[30] = 26'b00000000010001111010100010;
        x_t[31] = 26'b00000000010001011011000100;
        x_t[32] = 26'b00000000010101001010111101;
        x_t[33] = 26'b00000000010100111010000001;
        x_t[34] = 26'b00000000010010111101101010;
        x_t[35] = 26'b00000000010000001110011100;
        x_t[36] = 26'b00000000001110100000110001;
        x_t[37] = 26'b00000000001001111111100001;
        x_t[38] = 26'b00000000001001101110100011;
        x_t[39] = 26'b00000000001001100010010010;
        x_t[40] = 26'b00000000010000001001100111;
        x_t[41] = 26'b00000000001001101011110010;
        x_t[42] = 26'b00000000001010101001010011;
        x_t[43] = 26'b00000000100100110011111010;
        x_t[44] = 26'b00000000001100011101100001;
        x_t[45] = 26'b00000000010000011010100100;
        x_t[46] = 26'b00000000001001100000101101;
        x_t[47] = 26'b00000000001010101011100100;
        x_t[48] = 26'b00000000000110101110100010;
        x_t[49] = 26'b00000000001010001001110001;
        x_t[50] = 26'b00000000010001011011001101;
        x_t[51] = 26'b00000000010110011110110111;
        x_t[52] = 26'b00000000010111011111000110;
        x_t[53] = 26'b00000000011001101001100011;
        x_t[54] = 26'b00000000010111100010011000;
        x_t[55] = 26'b00000000000100011010100110;
        x_t[56] = 26'b00000000001010010001110101;
        x_t[57] = 26'b00000000001101011100110101;
        x_t[58] = 26'b00000000010110010100000010;
        x_t[59] = 26'b00000000001111111111010010;
        x_t[60] = 26'b00000000000110111001010010;
        x_t[61] = 26'b00000000001001110010100010;
        x_t[62] = 26'b00000000000011011011100100;
        x_t[63] = 26'b00000000001011110110000000;
        
        h_t_prev[0] = 26'b00000000001100010010010101;
        h_t_prev[1] = 26'b00000000010010100000110101;
        h_t_prev[2] = 26'b00000000010101111101000010;
        h_t_prev[3] = 26'b00000000011010011011110000;
        h_t_prev[4] = 26'b00000000010111010011100010;
        h_t_prev[5] = 26'b00000000010001001011000000;
        h_t_prev[6] = 26'b00000000001110001100001110;
        h_t_prev[7] = 26'b00000000000011001101110100;
        h_t_prev[8] = 26'b00000000010000001101111111;
        h_t_prev[9] = 26'b00000000010101011010011001;
        h_t_prev[10] = 26'b00000000011000011111111010;
        h_t_prev[11] = 26'b00000000011101001111111001;
        h_t_prev[12] = 26'b00000000010111010000000001;
        h_t_prev[13] = 26'b00000000001110001011101111;
        h_t_prev[14] = 26'b00000000001001100101110100;
        h_t_prev[15] = 26'b00000000010010010010000100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 7 timeout!");
                $fdisplay(fd_cycles, "Test Vector   7: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   7: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 7");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 8
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001100010010010101;
        x_t[1] = 26'b00000000010001010010100001;
        x_t[2] = 26'b00000000010100101111010110;
        x_t[3] = 26'b00000000011010101111000110;
        x_t[4] = 26'b00000000011000100100011000;
        x_t[5] = 26'b00000000010011100110010100;
        x_t[6] = 26'b00000000010010110110111101;
        x_t[7] = 26'b00000000000100011111010000;
        x_t[8] = 26'b00000000001101111101100101;
        x_t[9] = 26'b00000000010010010001111101;
        x_t[10] = 26'b00000000010110111110000100;
        x_t[11] = 26'b00000000011101001111111001;
        x_t[12] = 26'b00000000011001011100011111;
        x_t[13] = 26'b00000000010011010010110101;
        x_t[14] = 26'b00000000001001010000101110;
        x_t[15] = 26'b00000000010000000011101011;
        x_t[16] = 26'b00000000010001001000001101;
        x_t[17] = 26'b00000000010011000011101000;
        x_t[18] = 26'b00000000010110111010010101;
        x_t[19] = 26'b00000000011010000100010100;
        x_t[20] = 26'b00000000010111111101110010;
        x_t[21] = 26'b00000000001011001101101011;
        x_t[22] = 26'b00000000001000111011011010;
        x_t[23] = 26'b00000000001010011101001000;
        x_t[24] = 26'b00000000001011001001111110;
        x_t[25] = 26'b00000000001011110111010110;
        x_t[26] = 26'b00000000010000010101010001;
        x_t[27] = 26'b00000000001101100111001001;
        x_t[28] = 26'b00000000001100000001110100;
        x_t[29] = 26'b00000000001000101000000110;
        x_t[30] = 26'b00000000010000101100011111;
        x_t[31] = 26'b00000000010011000101100001;
        x_t[32] = 26'b00000000010101011101001000;
        x_t[33] = 26'b00000000010100100111100001;
        x_t[34] = 26'b00000000010011010000101101;
        x_t[35] = 26'b00000000010000100010001011;
        x_t[36] = 26'b00000000010001010011101011;
        x_t[37] = 26'b00000000001101110100001001;
        x_t[38] = 26'b00000000000110010000101100;
        x_t[39] = 26'b00000000001011110101010001;
        x_t[40] = 26'b00000000001100000100110000;
        x_t[41] = 26'b00000000001100010010101100;
        x_t[42] = 26'b00000000000110111100001001;
        x_t[43] = 26'b00000000010101000010100010;
        x_t[44] = 26'b00000000000110111000000001;
        x_t[45] = 26'b00000000010001110111011010;
        x_t[46] = 26'b00000000000110100110001100;
        x_t[47] = 26'b00000000001001001000000111;
        x_t[48] = 26'b00000000000101100010010011;
        x_t[49] = 26'b00000000001001010010001010;
        x_t[50] = 26'b00000000010000100010001100;
        x_t[51] = 26'b00000000010101111000001110;
        x_t[52] = 26'b00000000010101100100010101;
        x_t[53] = 26'b00000000011000010000011110;
        x_t[54] = 26'b00000000010100111010100101;
        x_t[55] = 26'b00000000000100101011110111;
        x_t[56] = 26'b00000000001010000000101001;
        x_t[57] = 26'b00000000001101001011110001;
        x_t[58] = 26'b00000000010011110111000000;
        x_t[59] = 26'b00000000001011100011000101;
        x_t[60] = 26'b00000000000100011111111100;
        x_t[61] = 26'b00000000000110111100011101;
        x_t[62] = 26'b00000000000001100101001101;
        x_t[63] = 26'b00000000000101110010110000;
        
        h_t_prev[0] = 26'b00000000001100010010010101;
        h_t_prev[1] = 26'b00000000010001010010100001;
        h_t_prev[2] = 26'b00000000010100101111010110;
        h_t_prev[3] = 26'b00000000011010101111000110;
        h_t_prev[4] = 26'b00000000011000100100011000;
        h_t_prev[5] = 26'b00000000010011100110010100;
        h_t_prev[6] = 26'b00000000010010110110111101;
        h_t_prev[7] = 26'b00000000000100011111010000;
        h_t_prev[8] = 26'b00000000001101111101100101;
        h_t_prev[9] = 26'b00000000010010010001111101;
        h_t_prev[10] = 26'b00000000010110111110000100;
        h_t_prev[11] = 26'b00000000011101001111111001;
        h_t_prev[12] = 26'b00000000011001011100011111;
        h_t_prev[13] = 26'b00000000010011010010110101;
        h_t_prev[14] = 26'b00000000001001010000101110;
        h_t_prev[15] = 26'b00000000010000000011101011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 8 timeout!");
                $fdisplay(fd_cycles, "Test Vector   8: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   8: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 8");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 9
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001011101010111000;
        x_t[1] = 26'b00000000001110110101111010;
        x_t[2] = 26'b00000000010010111010110011;
        x_t[3] = 26'b00000000010111101101101111;
        x_t[4] = 26'b00000000010101101110100000;
        x_t[5] = 26'b00000000010001110111011000;
        x_t[6] = 26'b00000000010010110110111101;
        x_t[7] = 26'b00000000000010111001011101;
        x_t[8] = 26'b00000000001010011010101010;
        x_t[9] = 26'b00000000001110100001011011;
        x_t[10] = 26'b00000000010010101100000101;
        x_t[11] = 26'b00000000011010000100000011;
        x_t[12] = 26'b00000000010110001001110010;
        x_t[13] = 26'b00000000010100100100100110;
        x_t[14] = 26'b00000000000110111101000100;
        x_t[15] = 26'b00000000001100001111100100;
        x_t[16] = 26'b00000000001101101110000110;
        x_t[17] = 26'b00000000010000100101101101;
        x_t[18] = 26'b00000000010011010010011010;
        x_t[19] = 26'b00000000010101111100101110;
        x_t[20] = 26'b00000000010100000011100000;
        x_t[21] = 26'b00000000001101011101010110;
        x_t[22] = 26'b00000000001001010100110010;
        x_t[23] = 26'b00000000001011001011100010;
        x_t[24] = 26'b00000000001100101011011010;
        x_t[25] = 26'b00000000001101100111001111;
        x_t[26] = 26'b00000000010000100110001010;
        x_t[27] = 26'b00000000001100110111111110;
        x_t[28] = 26'b00000000001000111000010011;
        x_t[29] = 26'b00000000001001011010000000;
        x_t[30] = 26'b00000000010000101100011111;
        x_t[31] = 26'b00000000010001001001010101;
        x_t[32] = 26'b00000000010100100110100111;
        x_t[33] = 26'b00000000010010111000100000;
        x_t[34] = 26'b00000000010001011110011001;
        x_t[35] = 26'b00000000001111010011001110;
        x_t[36] = 26'b00000000001100010101100111;
        x_t[37] = 26'b00000000001011010001000100;
        x_t[38] = 26'b00000000001000001001101101;
        x_t[39] = 26'b00000000000110110001111010;
        x_t[40] = 26'b00000000001011011001010001;
        x_t[41] = 26'b00000000000110101001000011;
        x_t[42] = 26'b00000000000110111100001001;
        x_t[43] = 26'b00000000010010010010111111;
        x_t[44] = 26'b00000000000001101000111000;
        x_t[45] = 26'b00000000001000001100011000;
        x_t[46] = 26'b00000000001000110111010000;
        x_t[47] = 26'b00000000001010111111011110;
        x_t[48] = 26'b00000000000110001000011010;
        x_t[49] = 26'b00000000001010011100010011;
        x_t[50] = 26'b00000000001111000011001010;
        x_t[51] = 26'b00000000010011001010010111;
        x_t[52] = 26'b00000000010000110001011001;
        x_t[53] = 26'b00000000010001101001010110;
        x_t[54] = 26'b00000000001111010011000000;
        x_t[55] = 26'b00000000001010100111101010;
        x_t[56] = 26'b00000000001110010011101000;
        x_t[57] = 26'b00000000001111000011001001;
        x_t[58] = 26'b00000000010001011001111111;
        x_t[59] = 26'b00000000001000110101011010;
        x_t[60] = 26'b00000000000110011010101000;
        x_t[61] = 26'b00000000000111001101000000;
        x_t[62] = 26'b00000000000000101010000010;
        x_t[63] = 26'b00000000000101100001001001;
        
        h_t_prev[0] = 26'b00000000001011101010111000;
        h_t_prev[1] = 26'b00000000001110110101111010;
        h_t_prev[2] = 26'b00000000010010111010110011;
        h_t_prev[3] = 26'b00000000010111101101101111;
        h_t_prev[4] = 26'b00000000010101101110100000;
        h_t_prev[5] = 26'b00000000010001110111011000;
        h_t_prev[6] = 26'b00000000010010110110111101;
        h_t_prev[7] = 26'b00000000000010111001011101;
        h_t_prev[8] = 26'b00000000001010011010101010;
        h_t_prev[9] = 26'b00000000001110100001011011;
        h_t_prev[10] = 26'b00000000010010101100000101;
        h_t_prev[11] = 26'b00000000011010000100000011;
        h_t_prev[12] = 26'b00000000010110001001110010;
        h_t_prev[13] = 26'b00000000010100100100100110;
        h_t_prev[14] = 26'b00000000000110111101000100;
        h_t_prev[15] = 26'b00000000001100001111100100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 9 timeout!");
                $fdisplay(fd_cycles, "Test Vector   9: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector   9: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 9");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 10
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001000100101100100;
        x_t[1] = 26'b00000000001001101001000101;
        x_t[2] = 26'b00000000001100110110010110;
        x_t[3] = 26'b00000000010001000100010101;
        x_t[4] = 26'b00000000001111011010010110;
        x_t[5] = 26'b00000000001001100010110111;
        x_t[6] = 26'b00000000000111001100001000;
        x_t[7] = 26'b00000000000100001010111001;
        x_t[8] = 26'b00000000000111110101101000;
        x_t[9] = 26'b00000000001010001000110011;
        x_t[10] = 26'b00000000001101001011110101;
        x_t[11] = 26'b00000000010010011010110110;
        x_t[12] = 26'b00000000001101000000011110;
        x_t[13] = 26'b00000000000100011000110101;
        x_t[14] = 26'b00000000001001010000101110;
        x_t[15] = 26'b00000000001100111000010000;
        x_t[16] = 26'b00000000001100011110110010;
        x_t[17] = 26'b00000000001101001100100100;
        x_t[18] = 26'b00000000001101010110111001;
        x_t[19] = 26'b00000000001110000011011110;
        x_t[20] = 26'b00000000001001011111110000;
        x_t[21] = 26'b00000000001010000000010100;
        x_t[22] = 26'b00000000000101111101000001;
        x_t[23] = 26'b00000000000111010111111001;
        x_t[24] = 26'b00000000000110011001011111;
        x_t[25] = 26'b00000000000111011001011011;
        x_t[26] = 26'b00000000001001101110110110;
        x_t[27] = 26'b00000000000110101110111011;
        x_t[28] = 26'b00000000001000010010100000;
        x_t[29] = 26'b00000000000011101011111110;
        x_t[30] = 26'b00000000001001011000001011;
        x_t[31] = 26'b00000000000111101110000101;
        x_t[32] = 26'b00000000001010111100110001;
        x_t[33] = 26'b00000000001001101000011011;
        x_t[34] = 26'b00000000001000001111110010;
        x_t[35] = 26'b00000000000100100000011010;
        x_t[36] = 26'b00000000000000110110000100;
        x_t[37] = 26'b00000000000100101001000100;
        x_t[38] = 26'b00000000000011101111010101;
        x_t[39] = 26'b11111111111101001000100101;
        x_t[40] = 26'b00000000000100100110100000;
        x_t[41] = 26'b11111111111110011000100000;
        x_t[42] = 26'b00000000000110001100101101;
        x_t[43] = 26'b00000000010001100111000110;
        x_t[44] = 26'b00000000001100000111001011;
        x_t[45] = 26'b00000000001001101001001111;
        x_t[46] = 26'b00000000010101001010101101;
        x_t[47] = 26'b00000000010001001101010101;
        x_t[48] = 26'b00000000001001011010000100;
        x_t[49] = 26'b00000000001101101000001011;
        x_t[50] = 26'b00000000001110011101001001;
        x_t[51] = 26'b00000000001111100010100011;
        x_t[52] = 26'b00000000001100100111011000;
        x_t[53] = 26'b00000000001101110100011001;
        x_t[54] = 26'b00000000001101110011000111;
        x_t[55] = 26'b00000000010001010111001111;
        x_t[56] = 26'b00000000010101000001010011;
        x_t[57] = 26'b00000000010001001011100100;
        x_t[58] = 26'b00000000010000010100001100;
        x_t[59] = 26'b00000000001010100011111011;
        x_t[60] = 26'b00000000001100001010101010;
        x_t[61] = 26'b00000000001100011000000101;
        x_t[62] = 26'b00000000000011001100110001;
        x_t[63] = 26'b00000000001100011001001101;
        
        h_t_prev[0] = 26'b00000000001000100101100100;
        h_t_prev[1] = 26'b00000000001001101001000101;
        h_t_prev[2] = 26'b00000000001100110110010110;
        h_t_prev[3] = 26'b00000000010001000100010101;
        h_t_prev[4] = 26'b00000000001111011010010110;
        h_t_prev[5] = 26'b00000000001001100010110111;
        h_t_prev[6] = 26'b00000000000111001100001000;
        h_t_prev[7] = 26'b00000000000100001010111001;
        h_t_prev[8] = 26'b00000000000111110101101000;
        h_t_prev[9] = 26'b00000000001010001000110011;
        h_t_prev[10] = 26'b00000000001101001011110101;
        h_t_prev[11] = 26'b00000000010010011010110110;
        h_t_prev[12] = 26'b00000000001101000000011110;
        h_t_prev[13] = 26'b00000000000100011000110101;
        h_t_prev[14] = 26'b00000000001001010000101110;
        h_t_prev[15] = 26'b00000000001100111000010000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 10 timeout!");
                $fdisplay(fd_cycles, "Test Vector  10: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  10: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 10");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 11
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000011000010011010;
        x_t[1] = 26'b00000000000011100001100011;
        x_t[2] = 26'b00000000000101010000110001;
        x_t[3] = 26'b00000000001000010011100110;
        x_t[4] = 26'b00000000000110100100100001;
        x_t[5] = 26'b11111111111111110101100101;
        x_t[6] = 26'b11111111111101110110101011;
        x_t[7] = 26'b11111111111111101101111000;
        x_t[8] = 26'b00000000000110001110011111;
        x_t[9] = 26'b00000000000111010100011001;
        x_t[10] = 26'b00000000001000100110010010;
        x_t[11] = 26'b00000000001000110111010110;
        x_t[12] = 26'b00000000000101101100001101;
        x_t[13] = 26'b11111111111101111111111110;
        x_t[14] = 26'b00000000001100001110100101;
        x_t[15] = 26'b00000000001110001001100111;
        x_t[16] = 26'b00000000001100001010111110;
        x_t[17] = 26'b00000000001011010110001000;
        x_t[18] = 26'b00000000001000101111101110;
        x_t[19] = 26'b00000000001000100100000000;
        x_t[20] = 26'b00000000000101100101011110;
        x_t[21] = 26'b00000000000011100111011011;
        x_t[22] = 26'b00000000000001001100011001;
        x_t[23] = 26'b00000000000011000001011101;
        x_t[24] = 26'b00000000000011100010110011;
        x_t[25] = 26'b00000000000100000110000101;
        x_t[26] = 26'b00000000000010000100110101;
        x_t[27] = 26'b11111111111110110111110101;
        x_t[28] = 26'b00000000000011100100001110;
        x_t[29] = 26'b00000000000001010110001110;
        x_t[30] = 26'b00000000000111011011010010;
        x_t[31] = 26'b00000000000011000000011101;
        x_t[32] = 26'b00000000000110011010000001;
        x_t[33] = 26'b00000000000100001000111000;
        x_t[34] = 26'b00000000000001101100101000;
        x_t[35] = 26'b11111111111110111101001000;
        x_t[36] = 26'b11111111111010111100010111;
        x_t[37] = 26'b11111111111111110011001110;
        x_t[38] = 26'b00000000000110111001000001;
        x_t[39] = 26'b11111111111001011101011010;
        x_t[40] = 26'b00000000001110110010101010;
        x_t[41] = 26'b00000000001000110100001001;
        x_t[42] = 26'b00000000010000100100110001;
        x_t[43] = 26'b00000000000011001101100000;
        x_t[44] = 26'b00000000010011011100011000;
        x_t[45] = 26'b00000000000111101101011011;
        x_t[46] = 26'b00000000010110011101100110;
        x_t[47] = 26'b00000000010100010100010000;
        x_t[48] = 26'b00000000001011011111011110;
        x_t[49] = 26'b00000000001111010111010111;
        x_t[50] = 26'b00000000001101110111001001;
        x_t[51] = 26'b00000000001101011011010100;
        x_t[52] = 26'b00000000001010000011101011;
        x_t[53] = 26'b00000000001100000101000011;
        x_t[54] = 26'b00000000001101000011001011;
        x_t[55] = 26'b00000000010101101011011101;
        x_t[56] = 26'b00000000011000001111100010;
        x_t[57] = 26'b00000000010010110001111000;
        x_t[58] = 26'b00000000001111001110011010;
        x_t[59] = 26'b00000000001010110011101110;
        x_t[60] = 26'b00000000010010111000000010;
        x_t[61] = 26'b00000000010010010100110100;
        x_t[62] = 26'b00000000000110001101000111;
        x_t[63] = 26'b00000000010101001100100000;
        
        h_t_prev[0] = 26'b00000000000011000010011010;
        h_t_prev[1] = 26'b00000000000011100001100011;
        h_t_prev[2] = 26'b00000000000101010000110001;
        h_t_prev[3] = 26'b00000000001000010011100110;
        h_t_prev[4] = 26'b00000000000110100100100001;
        h_t_prev[5] = 26'b11111111111111110101100101;
        h_t_prev[6] = 26'b11111111111101110110101011;
        h_t_prev[7] = 26'b11111111111111101101111000;
        h_t_prev[8] = 26'b00000000000110001110011111;
        h_t_prev[9] = 26'b00000000000111010100011001;
        h_t_prev[10] = 26'b00000000001000100110010010;
        h_t_prev[11] = 26'b00000000001000110111010110;
        h_t_prev[12] = 26'b00000000000101101100001101;
        h_t_prev[13] = 26'b11111111111101111111111110;
        h_t_prev[14] = 26'b00000000001100001110100101;
        h_t_prev[15] = 26'b00000000001110001001100111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 11 timeout!");
                $fdisplay(fd_cycles, "Test Vector  11: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  11: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 11");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 12
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001010011011111101;
        x_t[1] = 26'b00000000001000000111001101;
        x_t[2] = 26'b00000000000111111111100101;
        x_t[3] = 26'b00000000001000010011100110;
        x_t[4] = 26'b00000000000110010000010100;
        x_t[5] = 26'b11111111111110011100110101;
        x_t[6] = 26'b11111111111101011101110001;
        x_t[7] = 26'b00000000000110101101110001;
        x_t[8] = 26'b00000000001001110001011010;
        x_t[9] = 26'b00000000001000100100100101;
        x_t[10] = 26'b00000000000111000100011100;
        x_t[11] = 26'b00000000000111100101110100;
        x_t[12] = 26'b00000000000011001000010101;
        x_t[13] = 26'b11111111111101100100101101;
        x_t[14] = 26'b00000000010000001011101101;
        x_t[15] = 26'b00000000001111101111010101;
        x_t[16] = 26'b00000000001011110111001001;
        x_t[17] = 26'b00000000001000100100011110;
        x_t[18] = 26'b00000000000101011100111000;
        x_t[19] = 26'b00000000000110001010001111;
        x_t[20] = 26'b00000000000010110110010010;
        x_t[21] = 26'b00000000000101100000111111;
        x_t[22] = 26'b00000000000001111111001010;
        x_t[23] = 26'b00000000000001110000010000;
        x_t[24] = 26'b00000000000110001101010100;
        x_t[25] = 26'b00000000000110100111101100;
        x_t[26] = 26'b00000000000011001000011011;
        x_t[27] = 26'b11111111111111010111010001;
        x_t[28] = 26'b00000000000010001100000100;
        x_t[29] = 26'b00000000000111110110001011;
        x_t[30] = 26'b00000000001000101001010101;
        x_t[31] = 26'b00000000000011010010001100;
        x_t[32] = 26'b00000000001000111101100100;
        x_t[33] = 26'b00000000000111000001111001;
        x_t[34] = 26'b00000000000011110010000000;
        x_t[35] = 26'b00000000000001011011000010;
        x_t[36] = 26'b11111111111100001011111000;
        x_t[37] = 26'b00000000000000110100011101;
        x_t[38] = 26'b00000000001001011010011000;
        x_t[39] = 26'b11111111110111001010011011;
        x_t[40] = 26'b00000000010011001101010001;
        x_t[41] = 26'b11111111111100001101011011;
        x_t[42] = 26'b00000000010110100000001110;
        x_t[43] = 26'b11111111110100110011111001;
        x_t[44] = 26'b00000000010011110010101110;
        x_t[45] = 26'b11111111111111111110001100;
        x_t[46] = 26'b00000000010100110101111111;
        x_t[47] = 26'b00000000010100010100010000;
        x_t[48] = 26'b00000000001011011111011110;
        x_t[49] = 26'b00000000001101101000001011;
        x_t[50] = 26'b00000000001011001100000110;
        x_t[51] = 26'b00000000001010000110110100;
        x_t[52] = 26'b00000000000101010000101111;
        x_t[53] = 26'b00000000000110110111000000;
        x_t[54] = 26'b00000000000101111011101101;
        x_t[55] = 26'b00000000010101001000111011;
        x_t[56] = 26'b00000000010111001010110010;
        x_t[57] = 26'b00000000010001101101101010;
        x_t[58] = 26'b00000000001011001000101100;
        x_t[59] = 26'b00000000000101001000100100;
        x_t[60] = 26'b00000000010101010001011000;
        x_t[61] = 26'b00000000010100001000101100;
        x_t[62] = 26'b00000000000101111110010100;
        x_t[63] = 26'b00000000010111101010111011;
        
        h_t_prev[0] = 26'b00000000001010011011111101;
        h_t_prev[1] = 26'b00000000001000000111001101;
        h_t_prev[2] = 26'b00000000000111111111100101;
        h_t_prev[3] = 26'b00000000001000010011100110;
        h_t_prev[4] = 26'b00000000000110010000010100;
        h_t_prev[5] = 26'b11111111111110011100110101;
        h_t_prev[6] = 26'b11111111111101011101110001;
        h_t_prev[7] = 26'b00000000000110101101110001;
        h_t_prev[8] = 26'b00000000001001110001011010;
        h_t_prev[9] = 26'b00000000001000100100100101;
        h_t_prev[10] = 26'b00000000000111000100011100;
        h_t_prev[11] = 26'b00000000000111100101110100;
        h_t_prev[12] = 26'b00000000000011001000010101;
        h_t_prev[13] = 26'b11111111111101100100101101;
        h_t_prev[14] = 26'b00000000010000001011101101;
        h_t_prev[15] = 26'b00000000001111101111010101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 12 timeout!");
                $fdisplay(fd_cycles, "Test Vector  12: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  12: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 12");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 13
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001010101111101011;
        x_t[1] = 26'b00000000001001000001111100;
        x_t[2] = 26'b00000000001000100110011011;
        x_t[3] = 26'b00000000001000111010010001;
        x_t[4] = 26'b00000000000100111111011110;
        x_t[5] = 26'b11111111111100010111101101;
        x_t[6] = 26'b11111111111011111010001101;
        x_t[7] = 26'b00000000000111111111001101;
        x_t[8] = 26'b00000000001001001000001001;
        x_t[9] = 26'b00000000000111000000010110;
        x_t[10] = 26'b00000000000110011101010011;
        x_t[11] = 26'b00000000000110010100010001;
        x_t[12] = 26'b11111111111111110101100111;
        x_t[13] = 26'b11111111111000111000111000;
        x_t[14] = 26'b00000000001111110110100111;
        x_t[15] = 26'b00000000001101110101010010;
        x_t[16] = 26'b00000000001010000000001011;
        x_t[17] = 26'b00000000000110000110100011;
        x_t[18] = 26'b00000000000100011101101000;
        x_t[19] = 26'b00000000000100011100011001;
        x_t[20] = 26'b00000000000000000111000110;
        x_t[21] = 26'b00000000000110000010001001;
        x_t[22] = 26'b00000000000000011001100111;
        x_t[23] = 26'b00000000000001000001110101;
        x_t[24] = 26'b00000000000111100010100100;
        x_t[25] = 26'b00000000001000001011001001;
        x_t[26] = 26'b00000000000001110011111100;
        x_t[27] = 26'b11111111111111000111100011;
        x_t[28] = 26'b00000000000001111111011110;
        x_t[29] = 26'b00000000001010111101110101;
        x_t[30] = 26'b00000000000101101110000000;
        x_t[31] = 26'b00000000000011000000011101;
        x_t[32] = 26'b00000000000111100010101101;
        x_t[33] = 26'b00000000000100101101111000;
        x_t[34] = 26'b00000000000001101100101000;
        x_t[35] = 26'b11111111111110000001111010;
        x_t[36] = 26'b11111111111011010000001111;
        x_t[37] = 26'b00000000000001000100110001;
        x_t[38] = 26'b00000000001100001111111010;
        x_t[39] = 26'b11111111110011011111010000;
        x_t[40] = 26'b00000000010101100101011100;
        x_t[41] = 26'b11111111110000111010001001;
        x_t[42] = 26'b00000000010010110011000100;
        x_t[43] = 26'b00000000010111110010000101;
        x_t[44] = 26'b00000000010011011100011000;
        x_t[45] = 26'b11111111111110100001010101;
        x_t[46] = 26'b00000000010010100100111011;
        x_t[47] = 26'b00000000010000111001011011;
        x_t[48] = 26'b00000000001000110011111100;
        x_t[49] = 26'b00000000001100001011100000;
        x_t[50] = 26'b00000000001010100110000101;
        x_t[51] = 26'b00000000001001100000001011;
        x_t[52] = 26'b00000000000100111100010001;
        x_t[53] = 26'b00000000000101011101111011;
        x_t[54] = 26'b00000000000010001100000000;
        x_t[55] = 26'b00000000001110101010100111;
        x_t[56] = 26'b00000000010010000100001111;
        x_t[57] = 26'b00000000001110001111111111;
        x_t[58] = 26'b00000000001000001000110001;
        x_t[59] = 26'b00000000000000111100001010;
        x_t[60] = 26'b00000000010010001010000001;
        x_t[61] = 26'b00000000010000010000011000;
        x_t[62] = 26'b00000000000001110100000000;
        x_t[63] = 26'b00000000001111111110000011;
        
        h_t_prev[0] = 26'b00000000001010101111101011;
        h_t_prev[1] = 26'b00000000001001000001111100;
        h_t_prev[2] = 26'b00000000001000100110011011;
        h_t_prev[3] = 26'b00000000001000111010010001;
        h_t_prev[4] = 26'b00000000000100111111011110;
        h_t_prev[5] = 26'b11111111111100010111101101;
        h_t_prev[6] = 26'b11111111111011111010001101;
        h_t_prev[7] = 26'b00000000000111111111001101;
        h_t_prev[8] = 26'b00000000001001001000001001;
        h_t_prev[9] = 26'b00000000000111000000010110;
        h_t_prev[10] = 26'b00000000000110011101010011;
        h_t_prev[11] = 26'b00000000000110010100010001;
        h_t_prev[12] = 26'b11111111111111110101100111;
        h_t_prev[13] = 26'b11111111111000111000111000;
        h_t_prev[14] = 26'b00000000001111110110100111;
        h_t_prev[15] = 26'b00000000001101110101010010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 13 timeout!");
                $fdisplay(fd_cycles, "Test Vector  13: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  13: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 13");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 14
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000111101010011000;
        x_t[1] = 26'b00000000000010111010011001;
        x_t[2] = 26'b00000000000100000011000101;
        x_t[3] = 26'b00000000000110011111100100;
        x_t[4] = 26'b11111111111110111111100001;
        x_t[5] = 26'b11111111110110011110100000;
        x_t[6] = 26'b11111111110110110110100101;
        x_t[7] = 26'b00000000000000010110100110;
        x_t[8] = 26'b00000000000011010100110100;
        x_t[9] = 26'b00000000000011001111110100;
        x_t[10] = 26'b00000000000100000000101111;
        x_t[11] = 26'b00000000000001110110111010;
        x_t[12] = 26'b11111111111010101101110101;
        x_t[13] = 26'b11111111110101111010000101;
        x_t[14] = 26'b00000000000111100111010000;
        x_t[15] = 26'b00000000000111011110011100;
        x_t[16] = 26'b00000000000100011011010010;
        x_t[17] = 26'b00000000000010011001101011;
        x_t[18] = 26'b00000000000001001010110010;
        x_t[19] = 26'b00000000000000010100110010;
        x_t[20] = 26'b11111111111011011010110000;
        x_t[21] = 26'b00000000000011010001010101;
        x_t[22] = 26'b11111111111010011100110101;
        x_t[23] = 26'b11111111111011011010001100;
        x_t[24] = 26'b00000000000101101000110001;
        x_t[25] = 26'b00000000000110001110110101;
        x_t[26] = 26'b11111111111001111001000010;
        x_t[27] = 26'b11111111110111000000101111;
        x_t[28] = 26'b11111111111011011111110101;
        x_t[29] = 26'b00000000000111000100010001;
        x_t[30] = 26'b00000000000010100011000100;
        x_t[31] = 26'b11111111111100010110101000;
        x_t[32] = 26'b00000000000001110111010001;
        x_t[33] = 26'b11111111111100100111110011;
        x_t[34] = 26'b11111111111001000100000111;
        x_t[35] = 26'b11111111110111100011011011;
        x_t[36] = 26'b11111111110010100011101000;
        x_t[37] = 26'b11111111111010011100110001;
        x_t[38] = 26'b00000000001010111111001110;
        x_t[39] = 26'b11111111101101000011101101;
        x_t[40] = 26'b00000000010010001100000011;
        x_t[41] = 26'b11111111110100011000101100;
        x_t[42] = 26'b00000000000101110100111111;
        x_t[43] = 26'b00000000010101101110011011;
        x_t[44] = 26'b00000000000111111011000011;
        x_t[45] = 26'b11111111101100101000000111;
        x_t[46] = 26'b00000000000111001111101001;
        x_t[47] = 26'b00000000000111100100101001;
        x_t[48] = 26'b00000000000001000100011010;
        x_t[49] = 26'b00000000000100010111000110;
        x_t[50] = 26'b00000000000011011101111101;
        x_t[51] = 26'b00000000000010100011110110;
        x_t[52] = 26'b11111111111101100101101001;
        x_t[53] = 26'b11111111111100000100101001;
        x_t[54] = 26'b11111111110101011100111101;
        x_t[55] = 26'b00000000000101110000111010;
        x_t[56] = 26'b00000000001001101111011101;
        x_t[57] = 26'b00000000000111010100101000;
        x_t[58] = 26'b00000000000000110001101100;
        x_t[59] = 26'b11111111111010110001011011;
        x_t[60] = 26'b00000000001010011111010100;
        x_t[61] = 26'b00000000001000001111001110;
        x_t[62] = 26'b11111111111010001011110001;
        x_t[63] = 26'b00000000000100001001001000;
        
        h_t_prev[0] = 26'b00000000000111101010011000;
        h_t_prev[1] = 26'b00000000000010111010011001;
        h_t_prev[2] = 26'b00000000000100000011000101;
        h_t_prev[3] = 26'b00000000000110011111100100;
        h_t_prev[4] = 26'b11111111111110111111100001;
        h_t_prev[5] = 26'b11111111110110011110100000;
        h_t_prev[6] = 26'b11111111110110110110100101;
        h_t_prev[7] = 26'b00000000000000010110100110;
        h_t_prev[8] = 26'b00000000000011010100110100;
        h_t_prev[9] = 26'b00000000000011001111110100;
        h_t_prev[10] = 26'b00000000000100000000101111;
        h_t_prev[11] = 26'b00000000000001110110111010;
        h_t_prev[12] = 26'b11111111111010101101110101;
        h_t_prev[13] = 26'b11111111110101111010000101;
        h_t_prev[14] = 26'b00000000000111100111010000;
        h_t_prev[15] = 26'b00000000000111011110011100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 14 timeout!");
                $fdisplay(fd_cycles, "Test Vector  14: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  14: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 14");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 15
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001001110100011111;
        x_t[1] = 26'b00000000000101101010100101;
        x_t[2] = 26'b00000000000101100100001100;
        x_t[3] = 26'b00000000000110110010111010;
        x_t[4] = 26'b00000000000000100100100100;
        x_t[5] = 26'b11111111110111001010111000;
        x_t[6] = 26'b11111111110011101111011011;
        x_t[7] = 26'b00000000000110101101110001;
        x_t[8] = 26'b00000000000111110101101000;
        x_t[9] = 26'b00000000001000010000100010;
        x_t[10] = 26'b00000000001001100001000000;
        x_t[11] = 26'b00000000001000100010111101;
        x_t[12] = 26'b11111111111110010111111101;
        x_t[13] = 26'b11111111111000000010011000;
        x_t[14] = 26'b00000000001010100101000111;
        x_t[15] = 26'b00000000001100100011111010;
        x_t[16] = 26'b00000000001001101100010110;
        x_t[17] = 26'b00000000001000100100011110;
        x_t[18] = 26'b00000000000111110000011110;
        x_t[19] = 26'b00000000000110110110001010;
        x_t[20] = 26'b11111111111111101110000100;
        x_t[21] = 26'b00000000000001100010110100;
        x_t[22] = 26'b11111111111011101000111111;
        x_t[23] = 26'b11111111111101011001110011;
        x_t[24] = 26'b00000000000100010011100001;
        x_t[25] = 26'b00000000000101011101000111;
        x_t[26] = 26'b11111111111110011000010010;
        x_t[27] = 26'b11111111111001101101101011;
        x_t[28] = 26'b11111111111101101010011000;
        x_t[29] = 26'b00000000000111100101100010;
        x_t[30] = 26'b00000000000011100001100001;
        x_t[31] = 26'b00000000000010001011001110;
        x_t[32] = 26'b00000000001001001111101111;
        x_t[33] = 26'b00000000000101010010111000;
        x_t[34] = 26'b00000000000001000110100010;
        x_t[35] = 26'b11111111111110111101001000;
        x_t[36] = 26'b11111111111000110001001101;
        x_t[37] = 26'b00000000000011000111001110;
        x_t[38] = 26'b00000000001110001000111011;
        x_t[39] = 26'b11111111111000000101001110;
        x_t[40] = 26'b00000000010000001001100111;
        x_t[41] = 26'b00000000000101110001011010;
        x_t[42] = 26'b00000000001100011111111000;
        x_t[43] = 26'b00000000001101011111110010;
        x_t[44] = 26'b00000000001011011010011111;
        x_t[45] = 26'b00000000000101110001100111;
        x_t[46] = 26'b00000000001100101111111011;
        x_t[47] = 26'b00000000001110011010010010;
        x_t[48] = 26'b00000000001000100000111000;
        x_t[49] = 26'b00000000001101000011000110;
        x_t[50] = 26'b00000000001101010001001000;
        x_t[51] = 26'b00000000001100100001010111;
        x_t[52] = 26'b00000000001000011101010111;
        x_t[53] = 26'b00000000000111111001110100;
        x_t[54] = 26'b00000000000110010011101100;
        x_t[55] = 26'b00000000001011111101111110;
        x_t[56] = 26'b00000000010000011101000111;
        x_t[57] = 26'b00000000001110100001000010;
        x_t[58] = 26'b00000000001000111101000111;
        x_t[59] = 26'b00000000000010011010111001;
        x_t[60] = 26'b00000000001000010101010011;
        x_t[61] = 26'b00000000000111011101100011;
        x_t[62] = 26'b11111111111001011111011001;
        x_t[63] = 26'b00000000000100001001001000;
        
        h_t_prev[0] = 26'b00000000001001110100011111;
        h_t_prev[1] = 26'b00000000000101101010100101;
        h_t_prev[2] = 26'b00000000000101100100001100;
        h_t_prev[3] = 26'b00000000000110110010111010;
        h_t_prev[4] = 26'b00000000000000100100100100;
        h_t_prev[5] = 26'b11111111110111001010111000;
        h_t_prev[6] = 26'b11111111110011101111011011;
        h_t_prev[7] = 26'b00000000000110101101110001;
        h_t_prev[8] = 26'b00000000000111110101101000;
        h_t_prev[9] = 26'b00000000001000010000100010;
        h_t_prev[10] = 26'b00000000001001100001000000;
        h_t_prev[11] = 26'b00000000001000100010111101;
        h_t_prev[12] = 26'b11111111111110010111111101;
        h_t_prev[13] = 26'b11111111111000000010011000;
        h_t_prev[14] = 26'b00000000001010100101000111;
        h_t_prev[15] = 26'b00000000001100100011111010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 15 timeout!");
                $fdisplay(fd_cycles, "Test Vector  15: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  15: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 15");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 16
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001101001101100010;
        x_t[1] = 26'b00000000001100101100110111;
        x_t[2] = 26'b00000000001101110000100111;
        x_t[3] = 26'b00000000001111110110111111;
        x_t[4] = 26'b00000000001100010000010000;
        x_t[5] = 26'b00000000000010010000111010;
        x_t[6] = 26'b11111111111110101000011101;
        x_t[7] = 26'b00000000001011011111001001;
        x_t[8] = 26'b00000000001110100110110110;
        x_t[9] = 26'b00000000001111001001100000;
        x_t[10] = 26'b00000000010001011101110100;
        x_t[11] = 26'b00000000010010000110011110;
        x_t[12] = 26'b00000000001011100010110100;
        x_t[13] = 26'b00000000000100011000110101;
        x_t[14] = 26'b00000000010010011111010111;
        x_t[15] = 26'b00000000010001111101101110;
        x_t[16] = 26'b00000000010001011100000010;
        x_t[17] = 26'b00000000010000010001111101;
        x_t[18] = 26'b00000000010000010100101001;
        x_t[19] = 26'b00000000001111110001010100;
        x_t[20] = 26'b00000000001001011111110000;
        x_t[21] = 26'b00000000000011111101100010;
        x_t[22] = 26'b00000000000000011001100111;
        x_t[23] = 26'b00000000000001001101011100;
        x_t[24] = 26'b00000000000100101011111000;
        x_t[25] = 26'b00000000000110001110110101;
        x_t[26] = 26'b00000000000011111011000111;
        x_t[27] = 26'b11111111111101111000111100;
        x_t[28] = 26'b00000000000000001110000111;
        x_t[29] = 26'b00000000000110110011101000;
        x_t[30] = 26'b00000000000011010001111010;
        x_t[31] = 26'b00000000000101100000001000;
        x_t[32] = 26'b00000000001010111100110001;
        x_t[33] = 26'b00000000001000001011111010;
        x_t[34] = 26'b00000000000100111110001101;
        x_t[35] = 26'b00000000000000110011100011;
        x_t[36] = 26'b11111111111100001011111000;
        x_t[37] = 26'b00000000000101101010010011;
        x_t[38] = 26'b00000000000110100100110110;
        x_t[39] = 26'b11111111111100001101110010;
        x_t[40] = 26'b00000000000111101010001001;
        x_t[41] = 26'b00000000000101110001011010;
        x_t[42] = 26'b00000000001100011111111000;
        x_t[43] = 26'b00000000001110110111100100;
        x_t[44] = 26'b00000000001010101101110011;
        x_t[45] = 26'b00000000001010100111001000;
        x_t[46] = 26'b00000000001111010101101101;
        x_t[47] = 26'b00000000010000111001011011;
        x_t[48] = 26'b00000000001000110011111100;
        x_t[49] = 26'b00000000001110110010010011;
        x_t[50] = 26'b00000000001111000011001010;
        x_t[51] = 26'b00000000001110101000100101;
        x_t[52] = 26'b00000000001011010101100001;
        x_t[53] = 26'b00000000001001010010111001;
        x_t[54] = 26'b00000000000101001011110001;
        x_t[55] = 26'b00000000001110101010100111;
        x_t[56] = 26'b00000000010010010101011011;
        x_t[57] = 26'b00000000010000000111010110;
        x_t[58] = 26'b00000000001011001000101100;
        x_t[59] = 26'b00000000000010111010011110;
        x_t[60] = 26'b00000000001100101001010101;
        x_t[61] = 26'b00000000001100011000000101;
        x_t[62] = 26'b11111111111111010001010000;
        x_t[63] = 26'b00000000001010011101111111;
        
        h_t_prev[0] = 26'b00000000001101001101100010;
        h_t_prev[1] = 26'b00000000001100101100110111;
        h_t_prev[2] = 26'b00000000001101110000100111;
        h_t_prev[3] = 26'b00000000001111110110111111;
        h_t_prev[4] = 26'b00000000001100010000010000;
        h_t_prev[5] = 26'b00000000000010010000111010;
        h_t_prev[6] = 26'b11111111111110101000011101;
        h_t_prev[7] = 26'b00000000001011011111001001;
        h_t_prev[8] = 26'b00000000001110100110110110;
        h_t_prev[9] = 26'b00000000001111001001100000;
        h_t_prev[10] = 26'b00000000010001011101110100;
        h_t_prev[11] = 26'b00000000010010000110011110;
        h_t_prev[12] = 26'b00000000001011100010110100;
        h_t_prev[13] = 26'b00000000000100011000110101;
        h_t_prev[14] = 26'b00000000010010011111010111;
        h_t_prev[15] = 26'b00000000010001111101101110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 16 timeout!");
                $fdisplay(fd_cycles, "Test Vector  16: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  16: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 16");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 17
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000010011010111100;
        x_t[1] = 26'b00000000000011100001100011;
        x_t[2] = 26'b11111111110011111101101010;
        x_t[3] = 26'b11111111110111111111011100;
        x_t[4] = 26'b11111111110110011101111010;
        x_t[5] = 26'b11111111110100011001011000;
        x_t[6] = 26'b11111111111001111101101110;
        x_t[7] = 26'b00000000001000100111111011;
        x_t[8] = 26'b00000000000000011011001010;
        x_t[9] = 26'b11111111111010001010100010;
        x_t[10] = 26'b11111111110101111100100010;
        x_t[11] = 26'b11111111101111011000101010;
        x_t[12] = 26'b11111111110000110101101100;
        x_t[13] = 26'b11111111110010111011010010;
        x_t[14] = 26'b00000000001100001110100101;
        x_t[15] = 26'b00000000000100010011000010;
        x_t[16] = 26'b11111111111011110000000111;
        x_t[17] = 26'b11111111110111111010100001;
        x_t[18] = 26'b11111111101111011000010001;
        x_t[19] = 26'b11111111101111110110010111;
        x_t[20] = 26'b11111111110100110001010010;
        x_t[21] = 26'b11111111111111011110001101;
        x_t[22] = 26'b00000000000011110001011001;
        x_t[23] = 26'b00000000000101000001000101;
        x_t[24] = 26'b00000000000010110010000101;
        x_t[25] = 26'b00000000000010010110001100;
        x_t[26] = 26'b11111111111000100100100011;
        x_t[27] = 26'b11111111111011111011001011;
        x_t[28] = 26'b00000000000111100000001000;
        x_t[29] = 26'b00000000000001100110110111;
        x_t[30] = 26'b00000000001000111000111100;
        x_t[31] = 26'b11111111111110110110010100;
        x_t[32] = 26'b11111111111100011110000000;
        x_t[33] = 26'b11111111111010100110010010;
        x_t[34] = 26'b11111111111001010111001011;
        x_t[35] = 26'b11111111110110111011111100;
        x_t[36] = 26'b11111111111110111110110011;
        x_t[37] = 26'b11111111101100011011110111;
        x_t[38] = 26'b00000000000100010111101010;
        x_t[39] = 26'b00000000000010001011111100;
        x_t[40] = 26'b00000000001000101011010111;
        x_t[41] = 26'b00000000000011100110010101;
        x_t[42] = 26'b00000000001100001000001011;
        x_t[43] = 26'b11111111111111000110001100;
        x_t[44] = 26'b00000000001101110110111001;
        x_t[45] = 26'b11111111111111111110001100;
        x_t[46] = 26'b00000000001101101110000110;
        x_t[47] = 26'b00000000001010111111011110;
        x_t[48] = 26'b00000000000111000001100101;
        x_t[49] = 26'b00000000000010100111111001;
        x_t[50] = 26'b11111111111010100011110011;
        x_t[51] = 26'b11111111110111101100011001;
        x_t[52] = 26'b11111111111000011110001111;
        x_t[53] = 26'b11111111111011101110011000;
        x_t[54] = 26'b00000000000100110011110011;
        x_t[55] = 26'b00000000000111000111001111;
        x_t[56] = 26'b00000000001010010001110101;
        x_t[57] = 26'b11111111111101001100101000;
        x_t[58] = 26'b11111111111100101011111110;
        x_t[59] = 26'b00000000001010100011111011;
        x_t[60] = 26'b00000000000001011000100110;
        x_t[61] = 26'b11111111111101000111011010;
        x_t[62] = 26'b11111111111110010110000101;
        x_t[63] = 26'b00000000000011110111100001;
        
        h_t_prev[0] = 26'b00000000000010011010111100;
        h_t_prev[1] = 26'b00000000000011100001100011;
        h_t_prev[2] = 26'b11111111110011111101101010;
        h_t_prev[3] = 26'b11111111110111111111011100;
        h_t_prev[4] = 26'b11111111110110011101111010;
        h_t_prev[5] = 26'b11111111110100011001011000;
        h_t_prev[6] = 26'b11111111111001111101101110;
        h_t_prev[7] = 26'b00000000001000100111111011;
        h_t_prev[8] = 26'b00000000000000011011001010;
        h_t_prev[9] = 26'b11111111111010001010100010;
        h_t_prev[10] = 26'b11111111110101111100100010;
        h_t_prev[11] = 26'b11111111101111011000101010;
        h_t_prev[12] = 26'b11111111110000110101101100;
        h_t_prev[13] = 26'b11111111110010111011010010;
        h_t_prev[14] = 26'b00000000001100001110100101;
        h_t_prev[15] = 26'b00000000000100010011000010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 17 timeout!");
                $fdisplay(fd_cycles, "Test Vector  17: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  17: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 17");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 18
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001010011011111101;
        x_t[1] = 26'b00000000001100000101101101;
        x_t[2] = 26'b00000000000000000110100101;
        x_t[3] = 26'b00000000000010100100001101;
        x_t[4] = 26'b11111111111110101011010100;
        x_t[5] = 26'b11111111111100010111101101;
        x_t[6] = 26'b11111111111111000001010110;
        x_t[7] = 26'b00000000010010110011011001;
        x_t[8] = 26'b00000000001001001000001001;
        x_t[9] = 26'b00000000000011100011110111;
        x_t[10] = 26'b00000000000000000010010101;
        x_t[11] = 26'b11111111111010110110011110;
        x_t[12] = 26'b11111111111100001011011111;
        x_t[13] = 26'b11111111111101100100101101;
        x_t[14] = 26'b00000000001100001110100101;
        x_t[15] = 26'b00000000001010000001001011;
        x_t[16] = 26'b00000000000011110011101000;
        x_t[17] = 26'b00000000000011000001001001;
        x_t[18] = 26'b11111111111011001111010010;
        x_t[19] = 26'b11111111111100111001000111;
        x_t[20] = 26'b00000000000000000111000110;
        x_t[21] = 26'b00000000000000101011100100;
        x_t[22] = 26'b00000000000101001010001111;
        x_t[23] = 26'b00000000000110010010010010;
        x_t[24] = 26'b00000000000101101000110001;
        x_t[25] = 26'b00000000000101011101000111;
        x_t[26] = 26'b11111111111110000111011000;
        x_t[27] = 26'b11111111111111100111000000;
        x_t[28] = 26'b00000000001000000101111010;
        x_t[29] = 26'b00000000000111100101100010;
        x_t[30] = 26'b00000000001111001110110101;
        x_t[31] = 26'b00000000000011110101101011;
        x_t[32] = 26'b00000000000100011010110100;
        x_t[33] = 26'b00000000000001001111110110;
        x_t[34] = 26'b11111111111110101110000111;
        x_t[35] = 26'b11111111111101011010011100;
        x_t[36] = 26'b00000000000001001001111101;
        x_t[37] = 26'b11111111101010101001101101;
        x_t[38] = 26'b00000000001110011101000110;
        x_t[39] = 26'b00000000000011000110101111;
        x_t[40] = 26'b00000000010011100011000000;
        x_t[41] = 26'b11111111111001100110100000;
        x_t[42] = 26'b00000000001100011111111000;
        x_t[43] = 26'b00000000001010000100010111;
        x_t[44] = 26'b00000000001101110110111001;
        x_t[45] = 26'b00000000000100110011101101;
        x_t[46] = 26'b00000000001000001101110100;
        x_t[47] = 26'b00000000001001101111111001;
        x_t[48] = 26'b00000000000111000001100101;
        x_t[49] = 26'b00000000000100010111000110;
        x_t[50] = 26'b00000000000000110010111010;
        x_t[51] = 26'b00000000000000011100101000;
        x_t[52] = 26'b00000000000000110010010001;
        x_t[53] = 26'b00000000000001111111001110;
        x_t[54] = 26'b00000000001000111011011111;
        x_t[55] = 26'b00000000000100011010100110;
        x_t[56] = 26'b00000000000111100101111101;
        x_t[57] = 26'b00000000000000001000001101;
        x_t[58] = 26'b00000000000100110111011001;
        x_t[59] = 26'b00000000001010110011101110;
        x_t[60] = 26'b11111111111101110010100100;
        x_t[61] = 26'b11111111111110101010101111;
        x_t[62] = 26'b00000000000100010110110000;
        x_t[63] = 26'b11111111111011010101110110;
        
        h_t_prev[0] = 26'b00000000001010011011111101;
        h_t_prev[1] = 26'b00000000001100000101101101;
        h_t_prev[2] = 26'b00000000000000000110100101;
        h_t_prev[3] = 26'b00000000000010100100001101;
        h_t_prev[4] = 26'b11111111111110101011010100;
        h_t_prev[5] = 26'b11111111111100010111101101;
        h_t_prev[6] = 26'b11111111111111000001010110;
        h_t_prev[7] = 26'b00000000010010110011011001;
        h_t_prev[8] = 26'b00000000001001001000001001;
        h_t_prev[9] = 26'b00000000000011100011110111;
        h_t_prev[10] = 26'b00000000000000000010010101;
        h_t_prev[11] = 26'b11111111111010110110011110;
        h_t_prev[12] = 26'b11111111111100001011011111;
        h_t_prev[13] = 26'b11111111111101100100101101;
        h_t_prev[14] = 26'b00000000001100001110100101;
        h_t_prev[15] = 26'b00000000001010000001001011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 18 timeout!");
                $fdisplay(fd_cycles, "Test Vector  18: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  18: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 18");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 19
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000010010011100111101;
        x_t[1] = 26'b00000000010000101011010111;
        x_t[2] = 26'b00000000000100111101010110;
        x_t[3] = 26'b00000000000101100101100100;
        x_t[4] = 26'b00000000000000010000010111;
        x_t[5] = 26'b11111111111110011100110101;
        x_t[6] = 26'b11111111111110101000011101;
        x_t[7] = 26'b00000000010101000001111010;
        x_t[8] = 26'b00000000001010000110000010;
        x_t[9] = 26'b00000000000110000100001110;
        x_t[10] = 26'b00000000000001110111110000;
        x_t[11] = 26'b00000000000000010000111111;
        x_t[12] = 26'b00000000000000111011110110;
        x_t[13] = 26'b11111111111101100100101101;
        x_t[14] = 26'b00000000001110001101001001;
        x_t[15] = 26'b00000000001010111110001101;
        x_t[16] = 26'b00000000000101101010100110;
        x_t[17] = 26'b00000000000110101110000010;
        x_t[18] = 26'b00000000000010011111001000;
        x_t[19] = 26'b00000000000101011110010011;
        x_t[20] = 26'b00000000000111001001100101;
        x_t[21] = 26'b00000000001010001011011000;
        x_t[22] = 26'b00000000001100011111111000;
        x_t[23] = 26'b00000000001010111111111011;
        x_t[24] = 26'b00000000010001110100010000;
        x_t[25] = 26'b00000000010001000111000000;
        x_t[26] = 26'b00000000000100001100000000;
        x_t[27] = 26'b00000000000010110011011000;
        x_t[28] = 26'b00000000001001010001011111;
        x_t[29] = 26'b00000000010011110011100001;
        x_t[30] = 26'b00000000011011101010111110;
        x_t[31] = 26'b00000000001010011111100000;
        x_t[32] = 26'b00000000001100000101011101;
        x_t[33] = 26'b00000000000111010100011010;
        x_t[34] = 26'b00000000000100011000000110;
        x_t[35] = 26'b00000000000010111101101110;
        x_t[36] = 26'b00000000000001011101110101;
        x_t[37] = 26'b11111111100111000101011001;
        x_t[38] = 26'b00000000011100010100100100;
        x_t[39] = 26'b11111111111110111110001011;
        x_t[40] = 26'b00000000011011101100101111;
        x_t[41] = 26'b11111111110000011110010101;
        x_t[42] = 26'b00000000010111001111101010;
        x_t[43] = 26'b00000000000000011101111101;
        x_t[44] = 26'b00000000010100011111011010;
        x_t[45] = 26'b00000000010100110001001000;
        x_t[46] = 26'b00000000001111000000111111;
        x_t[47] = 26'b00000000001111111101110000;
        x_t[48] = 26'b00000000001111111101010110;
        x_t[49] = 26'b00000000001101010101101000;
        x_t[50] = 26'b00000000001101110111001001;
        x_t[51] = 26'b00000000010001101001110001;
        x_t[52] = 26'b00000000010011111110000001;
        x_t[53] = 26'b00000000010100011011100000;
        x_t[54] = 26'b00000000010111111010010111;
        x_t[55] = 26'b00000000001011011011011100;
        x_t[56] = 26'b00000000001110100100110100;
        x_t[57] = 26'b00000000001101111110111011;
        x_t[58] = 26'b00000000010111111100101110;
        x_t[59] = 26'b00000000010111001001001011;
        x_t[60] = 26'b11111111111110000001111010;
        x_t[61] = 26'b00000000000001110001011000;
        x_t[62] = 26'b00000000000111110100101011;
        x_t[63] = 26'b11111111110100001100001011;
        
        h_t_prev[0] = 26'b00000000010010011100111101;
        h_t_prev[1] = 26'b00000000010000101011010111;
        h_t_prev[2] = 26'b00000000000100111101010110;
        h_t_prev[3] = 26'b00000000000101100101100100;
        h_t_prev[4] = 26'b00000000000000010000010111;
        h_t_prev[5] = 26'b11111111111110011100110101;
        h_t_prev[6] = 26'b11111111111110101000011101;
        h_t_prev[7] = 26'b00000000010101000001111010;
        h_t_prev[8] = 26'b00000000001010000110000010;
        h_t_prev[9] = 26'b00000000000110000100001110;
        h_t_prev[10] = 26'b00000000000001110111110000;
        h_t_prev[11] = 26'b00000000000000010000111111;
        h_t_prev[12] = 26'b00000000000000111011110110;
        h_t_prev[13] = 26'b11111111111101100100101101;
        h_t_prev[14] = 26'b00000000001110001101001001;
        h_t_prev[15] = 26'b00000000001010111110001101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 19 timeout!");
                $fdisplay(fd_cycles, "Test Vector  19: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  19: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 19");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 20
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000011100101000000101;
        x_t[1] = 26'b00000000011010110001011011;
        x_t[2] = 26'b00000000001111010001101111;
        x_t[3] = 26'b00000000001110000010111110;
        x_t[4] = 26'b00000000001011100111110110;
        x_t[5] = 26'b00000000001010111011100111;
        x_t[6] = 26'b00000000000111111101111011;
        x_t[7] = 26'b00000000011101010011001111;
        x_t[8] = 26'b00000000010101000011011011;
        x_t[9] = 26'b00000000010010100110000000;
        x_t[10] = 26'b00000000010000100011000110;
        x_t[11] = 26'b00000000001110010001110111;
        x_t[12] = 26'b00000000010011001110011110;
        x_t[13] = 26'b00000000001111111000110001;
        x_t[14] = 26'b00000000011000011011000011;
        x_t[15] = 26'b00000000010111101011110111;
        x_t[16] = 26'b00000000010010101011010101;
        x_t[17] = 26'b00000000010011010111010111;
        x_t[18] = 26'b00000000010100111011110100;
        x_t[19] = 26'b00000000011001101110010110;
        x_t[20] = 26'b00000000011100101010000111;
        x_t[21] = 26'b00000000001100001111111111;
        x_t[22] = 26'b00000000001100101100100100;
        x_t[23] = 26'b00000000001011001011100010;
        x_t[24] = 26'b00000000010001011011111001;
        x_t[25] = 26'b00000000010001010011011100;
        x_t[26] = 26'b00000000000111111000100100;
        x_t[27] = 26'b00000000000101010000100110;
        x_t[28] = 26'b00000000001010000011110111;
        x_t[29] = 26'b00000000001111011000101011;
        x_t[30] = 26'b00000000011011111010100101;
        x_t[31] = 26'b00000000001100011011101101;
        x_t[32] = 26'b00000000001101001110001001;
        x_t[33] = 26'b00000000001001111010111011;
        x_t[34] = 26'b00000000000111101001101011;
        x_t[35] = 26'b00000000000101101111010111;
        x_t[36] = 26'b00000000000101100000010001;
        x_t[37] = 26'b11111111101011001010010100;
        x_t[38] = 26'b00000000010110101001100000;
        x_t[39] = 26'b00000000001001100010010010;
        x_t[40] = 26'b00000000010110010000111010;
        x_t[41] = 26'b00000000000111000100110111;
        x_t[42] = 26'b00000000010100010001111011;
        x_t[43] = 26'b11111111111111000110001100;
        x_t[44] = 26'b00000000010101111000110010;
        x_t[45] = 26'b00000000100001010101111000;
        x_t[46] = 26'b00000000010010111001101001;
        x_t[47] = 26'b00000000010010001001000000;
        x_t[48] = 26'b00000000010001101111101101;
        x_t[49] = 26'b00000000010001101011101001;
        x_t[50] = 26'b00000000010010111010001110;
        x_t[51] = 26'b00000000011011111010100110;
        x_t[52] = 26'b00000000011110100001010010;
        x_t[53] = 26'b00000000011111001101110111;
        x_t[54] = 26'b00000000100000001001101111;
        x_t[55] = 26'b00000000001100100000100000;
        x_t[56] = 26'b00000000001110000010011100;
        x_t[57] = 26'b00000000010011010011111110;
        x_t[58] = 26'b00000000100010000010010010;
        x_t[59] = 26'b00000000011100110100010100;
        x_t[60] = 26'b00000000000010000110100110;
        x_t[61] = 26'b00000000001010100100001101;
        x_t[62] = 26'b00000000010000011000000101;
        x_t[63] = 26'b11111111111010001111011011;
        
        h_t_prev[0] = 26'b00000000011100101000000101;
        h_t_prev[1] = 26'b00000000011010110001011011;
        h_t_prev[2] = 26'b00000000001111010001101111;
        h_t_prev[3] = 26'b00000000001110000010111110;
        h_t_prev[4] = 26'b00000000001011100111110110;
        h_t_prev[5] = 26'b00000000001010111011100111;
        h_t_prev[6] = 26'b00000000000111111101111011;
        h_t_prev[7] = 26'b00000000011101010011001111;
        h_t_prev[8] = 26'b00000000010101000011011011;
        h_t_prev[9] = 26'b00000000010010100110000000;
        h_t_prev[10] = 26'b00000000010000100011000110;
        h_t_prev[11] = 26'b00000000001110010001110111;
        h_t_prev[12] = 26'b00000000010011001110011110;
        h_t_prev[13] = 26'b00000000001111111000110001;
        h_t_prev[14] = 26'b00000000011000011011000011;
        h_t_prev[15] = 26'b00000000010111101011110111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 20 timeout!");
                $fdisplay(fd_cycles, "Test Vector  20: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  20: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 20");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 21
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001011101010111000;
        x_t[1] = 26'b00000000001100101100110111;
        x_t[2] = 26'b00000000000100000011000101;
        x_t[3] = 26'b00000000000100011000001110;
        x_t[4] = 26'b00000000000110010000010100;
        x_t[5] = 26'b00000000000111110011111010;
        x_t[6] = 26'b00000000001010010011010010;
        x_t[7] = 26'b00000000001100110000100101;
        x_t[8] = 26'b00000000001000001010010000;
        x_t[9] = 26'b00000000000111000000010110;
        x_t[10] = 26'b00000000000110110000110111;
        x_t[11] = 26'b00000000000111111010001100;
        x_t[12] = 26'b00000000010001110000110101;
        x_t[13] = 26'b00000000010010110111100100;
        x_t[14] = 26'b00000000001100001110100101;
        x_t[15] = 26'b00000000001011100110111001;
        x_t[16] = 26'b00000000001000110000110111;
        x_t[17] = 26'b00000000001011101001110111;
        x_t[18] = 26'b00000000001110101011001110;
        x_t[19] = 26'b00000000010101010000110010;
        x_t[20] = 26'b00000000011011000110000000;
        x_t[21] = 26'b11111111111011101011000101;
        x_t[22] = 26'b00000000000000100110010100;
        x_t[23] = 26'b00000000000101100011111000;
        x_t[24] = 26'b11111111111100111000100001;
        x_t[25] = 26'b11111111111100111010000111;
        x_t[26] = 26'b11111111111100010001000111;
        x_t[27] = 26'b00000000000000100101111000;
        x_t[28] = 26'b00000000000110101101110000;
        x_t[29] = 26'b11111111111010110110010001;
        x_t[30] = 26'b00000000000100011111111101;
        x_t[31] = 26'b00000000000011100011111100;
        x_t[32] = 26'b11111111111101100110101100;
        x_t[33] = 26'b11111111111101011111010100;
        x_t[34] = 26'b11111111111111000001001010;
        x_t[35] = 26'b11111111111011100100000001;
        x_t[36] = 26'b00000000000101100000010001;
        x_t[37] = 26'b11111111101101111101101101;
        x_t[38] = 26'b11111111111110011000011100;
        x_t[39] = 26'b00000000001011110101010001;
        x_t[40] = 26'b00000000001001010110110110;
        x_t[41] = 26'b00000000001011011011000011;
        x_t[42] = 26'b00000000000010000111110101;
        x_t[43] = 26'b00000000010011101010110000;
        x_t[44] = 26'b00000000001000100111101111;
        x_t[45] = 26'b00000000011000101000101111;
        x_t[46] = 26'b00000000001000110111010000;
        x_t[47] = 26'b00000000001000110100001110;
        x_t[48] = 26'b00000000001000100000111000;
        x_t[49] = 26'b00000000001001100100101101;
        x_t[50] = 26'b00000000001101010001001000;
        x_t[51] = 26'b00000000010110011110110111;
        x_t[52] = 26'b00000000011000001000000010;
        x_t[53] = 26'b00000000011000010000011110;
        x_t[54] = 26'b00000000010100111010100101;
        x_t[55] = 26'b00000000000111011000100000;
        x_t[56] = 26'b00000000001001011110010001;
        x_t[57] = 26'b00000000010000101001011101;
        x_t[58] = 26'b00000000011100100101010101;
        x_t[59] = 26'b00000000010111001001001011;
        x_t[60] = 26'b00000000000011100010100110;
        x_t[61] = 26'b00000000010000110001011111;
        x_t[62] = 26'b00000000010110011000110000;
        x_t[63] = 26'b00000000000001101010101101;
        
        h_t_prev[0] = 26'b00000000001011101010111000;
        h_t_prev[1] = 26'b00000000001100101100110111;
        h_t_prev[2] = 26'b00000000000100000011000101;
        h_t_prev[3] = 26'b00000000000100011000001110;
        h_t_prev[4] = 26'b00000000000110010000010100;
        h_t_prev[5] = 26'b00000000000111110011111010;
        h_t_prev[6] = 26'b00000000001010010011010010;
        h_t_prev[7] = 26'b00000000001100110000100101;
        h_t_prev[8] = 26'b00000000001000001010010000;
        h_t_prev[9] = 26'b00000000000111000000010110;
        h_t_prev[10] = 26'b00000000000110110000110111;
        h_t_prev[11] = 26'b00000000000111111010001100;
        h_t_prev[12] = 26'b00000000010001110000110101;
        h_t_prev[13] = 26'b00000000010010110111100100;
        h_t_prev[14] = 26'b00000000001100001110100101;
        h_t_prev[15] = 26'b00000000001011100110111001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 21 timeout!");
                $fdisplay(fd_cycles, "Test Vector  21: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  21: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 21");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 22
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000011000010011010;
        x_t[1] = 26'b00000000000101101010100101;
        x_t[2] = 26'b11111111111110100101011101;
        x_t[3] = 26'b00000000000001000011100001;
        x_t[4] = 26'b00000000000100010111000100;
        x_t[5] = 26'b00000000000111000111100010;
        x_t[6] = 26'b00000000001010010011010010;
        x_t[7] = 26'b00000000001010110110011011;
        x_t[8] = 26'b00000000000011101001011101;
        x_t[9] = 26'b00000000000100001011111101;
        x_t[10] = 26'b00000000000101100010100101;
        x_t[11] = 26'b00000000001000001110100101;
        x_t[12] = 26'b00000000001111100100010110;
        x_t[13] = 26'b00000000010011010010110101;
        x_t[14] = 26'b00000000001011001111010011;
        x_t[15] = 26'b00000000001001101100110101;
        x_t[16] = 26'b00000000000111001101101110;
        x_t[17] = 26'b00000000001010101110101001;
        x_t[18] = 26'b00000000001100101100101110;
        x_t[19] = 26'b00000000010010001011000101;
        x_t[20] = 26'b00000000011000101111110101;
        x_t[21] = 26'b00000000000001100010110100;
        x_t[22] = 26'b00000000000100110000110111;
        x_t[23] = 26'b00000000000111000000101100;
        x_t[24] = 26'b00000000000110011001011111;
        x_t[25] = 26'b00000000000101011101000111;
        x_t[26] = 26'b11111111111110111010000101;
        x_t[27] = 26'b00000000000010000100001110;
        x_t[28] = 26'b00000000001000010010100000;
        x_t[29] = 26'b00000000000111110110001011;
        x_t[30] = 26'b00000000001111101110000011;
        x_t[31] = 26'b00000000000111001010100110;
        x_t[32] = 26'b00000000000010011011100111;
        x_t[33] = 26'b00000000000001110100110110;
        x_t[34] = 26'b00000000000001101100101000;
        x_t[35] = 26'b00000000000000001100000101;
        x_t[36] = 26'b00000000000110101111110010;
        x_t[37] = 26'b11111111101001111000110010;
        x_t[38] = 26'b00000000010000010110000111;
        x_t[39] = 26'b00000000001000001010000110;
        x_t[40] = 26'b00000000001101110001011100;
        x_t[41] = 26'b00000000000111111100100000;
        x_t[42] = 26'b00000000010111100111011000;
        x_t[43] = 26'b11111111111111000110001100;
        x_t[44] = 26'b00000000001110111001111011;
        x_t[45] = 26'b00000000010001011000011101;
        x_t[46] = 26'b00000000010001111011011111;
        x_t[47] = 26'b00000000010010001001000000;
        x_t[48] = 26'b00000000001111010111001111;
        x_t[49] = 26'b00000000001111101001111010;
        x_t[50] = 26'b00000000010001001000001100;
        x_t[51] = 26'b00000000010111101100001001;
        x_t[52] = 26'b00000000010111110011100100;
        x_t[53] = 26'b00000000010110100001001000;
        x_t[54] = 26'b00000000010011011010101100;
        x_t[55] = 26'b00000000010010101101100100;
        x_t[56] = 26'b00000000010011011010001011;
        x_t[57] = 26'b00000000010101011100011001;
        x_t[58] = 26'b00000000011100110110110010;
        x_t[59] = 26'b00000000010111001001001011;
        x_t[60] = 26'b00000000001000010101010011;
        x_t[61] = 26'b00000000010110001101000111;
        x_t[62] = 26'b00000000011001001010010011;
        x_t[63] = 26'b00000000001101001110000001;
        
        h_t_prev[0] = 26'b00000000000011000010011010;
        h_t_prev[1] = 26'b00000000000101101010100101;
        h_t_prev[2] = 26'b11111111111110100101011101;
        h_t_prev[3] = 26'b00000000000001000011100001;
        h_t_prev[4] = 26'b00000000000100010111000100;
        h_t_prev[5] = 26'b00000000000111000111100010;
        h_t_prev[6] = 26'b00000000001010010011010010;
        h_t_prev[7] = 26'b00000000001010110110011011;
        h_t_prev[8] = 26'b00000000000011101001011101;
        h_t_prev[9] = 26'b00000000000100001011111101;
        h_t_prev[10] = 26'b00000000000101100010100101;
        h_t_prev[11] = 26'b00000000001000001110100101;
        h_t_prev[12] = 26'b00000000001111100100010110;
        h_t_prev[13] = 26'b00000000010011010010110101;
        h_t_prev[14] = 26'b00000000001011001111010011;
        h_t_prev[15] = 26'b00000000001001101100110101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 22 timeout!");
                $fdisplay(fd_cycles, "Test Vector  22: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  22: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 22");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 23
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000010011000100011010;
        x_t[1] = 26'b00000000010000101011010111;
        x_t[2] = 26'b00000000000101100100001100;
        x_t[3] = 26'b00000000001000010011100110;
        x_t[4] = 26'b00000000000110100100100001;
        x_t[5] = 26'b00000000000111000111100010;
        x_t[6] = 26'b00000000001001111010011001;
        x_t[7] = 26'b00000000011010110000010111;
        x_t[8] = 26'b00000000001110010010001110;
        x_t[9] = 26'b00000000001010110000111001;
        x_t[10] = 26'b00000000001010101111010001;
        x_t[11] = 26'b00000000001001100000000111;
        x_t[12] = 26'b00000000001100101001000011;
        x_t[13] = 26'b00000000001110001011101111;
        x_t[14] = 26'b00000000011000011011000011;
        x_t[15] = 26'b00000000010001111101101110;
        x_t[16] = 26'b00000000001110000001111011;
        x_t[17] = 26'b00000000001110101111010001;
        x_t[18] = 26'b00000000001101010110111001;
        x_t[19] = 26'b00000000010001001001001011;
        x_t[20] = 26'b00000000010100011100100010;
        x_t[21] = 26'b00000000000111001111100000;
        x_t[22] = 26'b00000000001010101101101001;
        x_t[23] = 26'b00000000001011101110010101;
        x_t[24] = 26'b00000000001011101110100001;
        x_t[25] = 26'b00000000001011011110011111;
        x_t[26] = 26'b00000000000001010010001001;
        x_t[27] = 26'b00000000000100110001001010;
        x_t[28] = 26'b00000000001110110010001001;
        x_t[29] = 26'b00000000001101000010111100;
        x_t[30] = 26'b00000000010011100111110100;
        x_t[31] = 26'b00000000000101110001111000;
        x_t[32] = 26'b00000000000100101100111111;
        x_t[33] = 26'b00000000000010111110110111;
        x_t[34] = 26'b00000000000001101100101000;
        x_t[35] = 26'b11111111111111100100100110;
        x_t[36] = 26'b00000000000110001000000001;
        x_t[37] = 26'b11111111101111101111110110;
        x_t[38] = 26'b00000000010000101010010010;
        x_t[39] = 26'b00000000001001000100111001;
        x_t[40] = 26'b00000000010011100011000000;
        x_t[41] = 26'b00000000000011001010100000;
        x_t[42] = 26'b00000000010110110111111100;
        x_t[43] = 26'b00000000000101111101000011;
        x_t[44] = 26'b00000000011011000111111100;
        x_t[45] = 26'b00000000001101000001111001;
        x_t[46] = 26'b00000000011010000001100011;
        x_t[47] = 26'b00000000010101100011110101;
        x_t[48] = 26'b00000000010000110110100010;
        x_t[49] = 26'b00000000001111101001111010;
        x_t[50] = 26'b00000000001111010110001010;
        x_t[51] = 26'b00000000010100010111101001;
        x_t[52] = 26'b00000000010011101001100011;
        x_t[53] = 26'b00000000010010101100001010;
        x_t[54] = 26'b00000000010010010010110010;
        x_t[55] = 26'b00000000010011100001010110;
        x_t[56] = 26'b00000000010010100110100111;
        x_t[57] = 26'b00000000010010100000110100;
        x_t[58] = 26'b00000000011010001000010011;
        x_t[59] = 26'b00000000010110001010000001;
        x_t[60] = 26'b00000000001101010111010101;
        x_t[61] = 26'b00000000011001100100010100;
        x_t[62] = 26'b00000000011000111011100000;
        x_t[63] = 26'b00000000010100111010111001;
        
        h_t_prev[0] = 26'b00000000010011000100011010;
        h_t_prev[1] = 26'b00000000010000101011010111;
        h_t_prev[2] = 26'b00000000000101100100001100;
        h_t_prev[3] = 26'b00000000001000010011100110;
        h_t_prev[4] = 26'b00000000000110100100100001;
        h_t_prev[5] = 26'b00000000000111000111100010;
        h_t_prev[6] = 26'b00000000001001111010011001;
        h_t_prev[7] = 26'b00000000011010110000010111;
        h_t_prev[8] = 26'b00000000001110010010001110;
        h_t_prev[9] = 26'b00000000001010110000111001;
        h_t_prev[10] = 26'b00000000001010101111010001;
        h_t_prev[11] = 26'b00000000001001100000000111;
        h_t_prev[12] = 26'b00000000001100101001000011;
        h_t_prev[13] = 26'b00000000001110001011101111;
        h_t_prev[14] = 26'b00000000011000011011000011;
        h_t_prev[15] = 26'b00000000010001111101101110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 23 timeout!");
                $fdisplay(fd_cycles, "Test Vector  23: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  23: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 23");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 24
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000100010001010101;
        x_t[1] = 26'b00000000000110111000111001;
        x_t[2] = 26'b11111111111111011111101111;
        x_t[3] = 26'b00000000000011011110001101;
        x_t[4] = 26'b11111111111111100111111100;
        x_t[5] = 26'b11111111111110000110101001;
        x_t[6] = 26'b00000000000001101111100111;
        x_t[7] = 26'b00000000001100110000100101;
        x_t[8] = 26'b00000000000101100101001110;
        x_t[9] = 26'b00000000000101110000001011;
        x_t[10] = 26'b00000000000110001001101110;
        x_t[11] = 26'b00000000000000100101011000;
        x_t[12] = 26'b00000000000011110111001001;
        x_t[13] = 26'b00000000000001011010000010;
        x_t[14] = 26'b00000000010001110101001011;
        x_t[15] = 26'b00000000001100001111100100;
        x_t[16] = 26'b00000000001001000100101100;
        x_t[17] = 26'b00000000001010101110101001;
        x_t[18] = 26'b00000000000111011011011000;
        x_t[19] = 26'b00000000001010010001110101;
        x_t[20] = 26'b00000000001100001110111100;
        x_t[21] = 26'b11111111111010101000110010;
        x_t[22] = 26'b11111111111111001101011101;
        x_t[23] = 26'b00000000000010011110101010;
        x_t[24] = 26'b11111111111101000100101101;
        x_t[25] = 26'b11111111111101000110100011;
        x_t[26] = 26'b11111111110111010000000100;
        x_t[27] = 26'b11111111111010101100100100;
        x_t[28] = 26'b00000000000100111100011001;
        x_t[29] = 26'b11111111111100001001011110;
        x_t[30] = 26'b00000000000110011100110110;
        x_t[31] = 26'b11111111111110000001000101;
        x_t[32] = 26'b11111111111100110000001011;
        x_t[33] = 26'b11111111111010111000110010;
        x_t[34] = 26'b11111111111000110001000100;
        x_t[35] = 26'b11111111110101101101000000;
        x_t[36] = 26'b11111111111010000000101110;
        x_t[37] = 26'b11111111101010011001011001;
        x_t[38] = 26'b11111111111111101001000111;
        x_t[39] = 26'b11111111111101100101111111;
        x_t[40] = 26'b00000000010100111001111101;
        x_t[41] = 26'b11111111101110010011001111;
        x_t[42] = 26'b00000000010100101001101001;
        x_t[43] = 26'b00000000001000101100100101;
        x_t[44] = 26'b00000000011010110001100110;
        x_t[45] = 26'b00000000010001110111011010;
        x_t[46] = 26'b00000000011000101110101010;
        x_t[47] = 26'b00000000010011011000100101;
        x_t[48] = 26'b00000000010000010000011010;
        x_t[49] = 26'b00000000001110110010010011;
        x_t[50] = 26'b00000000001110001010001001;
        x_t[51] = 26'b00000000010011110001000000;
        x_t[52] = 26'b00000000010011101001100011;
        x_t[53] = 26'b00000000010011000010011011;
        x_t[54] = 26'b00000000010110011010011110;
        x_t[55] = 26'b00000000001111101111101010;
        x_t[56] = 26'b00000000010000101110010011;
        x_t[57] = 26'b00000000010001011100100111;
        x_t[58] = 26'b00000000011010111100101001;
        x_t[59] = 26'b00000000011001100111000100;
        x_t[60] = 26'b00000000001101100110101010;
        x_t[61] = 26'b00000000011001100100010100;
        x_t[62] = 26'b00000000011000000000010100;
        x_t[63] = 26'b00000000010100101001010011;
        
        h_t_prev[0] = 26'b00000000000100010001010101;
        h_t_prev[1] = 26'b00000000000110111000111001;
        h_t_prev[2] = 26'b11111111111111011111101111;
        h_t_prev[3] = 26'b00000000000011011110001101;
        h_t_prev[4] = 26'b11111111111111100111111100;
        h_t_prev[5] = 26'b11111111111110000110101001;
        h_t_prev[6] = 26'b00000000000001101111100111;
        h_t_prev[7] = 26'b00000000001100110000100101;
        h_t_prev[8] = 26'b00000000000101100101001110;
        h_t_prev[9] = 26'b00000000000101110000001011;
        h_t_prev[10] = 26'b00000000000110001001101110;
        h_t_prev[11] = 26'b00000000000000100101011000;
        h_t_prev[12] = 26'b00000000000011110111001001;
        h_t_prev[13] = 26'b00000000000001011010000010;
        h_t_prev[14] = 26'b00000000010001110101001011;
        h_t_prev[15] = 26'b00000000001100001111100100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 24 timeout!");
                $fdisplay(fd_cycles, "Test Vector  24: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  24: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 24");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 25
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000100100101000100;
        x_t[1] = 26'b00000000001001000001111100;
        x_t[2] = 26'b00000000000001111011000111;
        x_t[3] = 26'b00000000000100111110111001;
        x_t[4] = 26'b11111111111111111100001001;
        x_t[5] = 26'b11111111111100010111101101;
        x_t[6] = 26'b11111111111010101111100001;
        x_t[7] = 26'b00000000010101000001111010;
        x_t[8] = 26'b00000000001011000011111011;
        x_t[9] = 26'b00000000001010110000111001;
        x_t[10] = 26'b00000000001010001000001000;
        x_t[11] = 26'b00000000000101000010101111;
        x_t[12] = 26'b00000000000101101100001101;
        x_t[13] = 26'b11111111111111010001101111;
        x_t[14] = 26'b00000000011000011011000011;
        x_t[15] = 26'b00000000010011100011011011;
        x_t[16] = 26'b00000000001110000001111011;
        x_t[17] = 26'b00000000001111010110101111;
        x_t[18] = 26'b00000000001011000011010011;
        x_t[19] = 26'b00000000001100101011100111;
        x_t[20] = 26'b00000000001110100101000111;
        x_t[21] = 26'b11111111111110111101000011;
        x_t[22] = 26'b00000000000000100110010100;
        x_t[23] = 26'b00000000000010011110101010;
        x_t[24] = 26'b00000000000011010110101000;
        x_t[25] = 26'b00000000000010100010101000;
        x_t[26] = 26'b11111111111011101111010100;
        x_t[27] = 26'b11111111111010111100010010;
        x_t[28] = 26'b00000000000001111111011110;
        x_t[29] = 26'b00000000000000000011000010;
        x_t[30] = 26'b00000000001011110100010001;
        x_t[31] = 26'b00000000000001111001011110;
        x_t[32] = 26'b00000000000100001000101001;
        x_t[33] = 26'b00000000000010000111010110;
        x_t[34] = 26'b11111111111101100001111001;
        x_t[35] = 26'b11111111111011010000010001;
        x_t[36] = 26'b11111111111011010000001111;
        x_t[37] = 26'b11111111101010001001000101;
        x_t[38] = 26'b00000000000101101000010110;
        x_t[39] = 26'b11111111111011010011000000;
        x_t[40] = 26'b00000000001001101100100101;
        x_t[41] = 26'b11111111110010001101100110;
        x_t[42] = 26'b00000000001111000101111001;
        x_t[43] = 26'b00000000001010000100010111;
        x_t[44] = 26'b00000000010001010110010100;
        x_t[45] = 26'b00000000010100010010001011;
        x_t[46] = 26'b00000000010101011111011011;
        x_t[47] = 26'b00000000010101100011110101;
        x_t[48] = 26'b00000000010011100010000011;
        x_t[49] = 26'b00000000010010010000101101;
        x_t[50] = 26'b00000000010010000001001101;
        x_t[51] = 26'b00000000010100111110010001;
        x_t[52] = 26'b00000000010100010010011110;
        x_t[53] = 26'b00000000010011011000101101;
        x_t[54] = 26'b00000000010100111010100101;
        x_t[55] = 26'b00000000010001101000100000;
        x_t[56] = 26'b00000000010001100001110111;
        x_t[57] = 26'b00000000010001011100100111;
        x_t[58] = 26'b00000000011010001000010011;
        x_t[59] = 26'b00000000010111001001001011;
        x_t[60] = 26'b00000000001100011001111111;
        x_t[61] = 26'b00000000010111110000011100;
        x_t[62] = 26'b00000000010110001001111101;
        x_t[63] = 26'b00000000010001010110000100;
        
        h_t_prev[0] = 26'b00000000000100100101000100;
        h_t_prev[1] = 26'b00000000001001000001111100;
        h_t_prev[2] = 26'b00000000000001111011000111;
        h_t_prev[3] = 26'b00000000000100111110111001;
        h_t_prev[4] = 26'b11111111111111111100001001;
        h_t_prev[5] = 26'b11111111111100010111101101;
        h_t_prev[6] = 26'b11111111111010101111100001;
        h_t_prev[7] = 26'b00000000010101000001111010;
        h_t_prev[8] = 26'b00000000001011000011111011;
        h_t_prev[9] = 26'b00000000001010110000111001;
        h_t_prev[10] = 26'b00000000001010001000001000;
        h_t_prev[11] = 26'b00000000000101000010101111;
        h_t_prev[12] = 26'b00000000000101101100001101;
        h_t_prev[13] = 26'b11111111111111010001101111;
        h_t_prev[14] = 26'b00000000011000011011000011;
        h_t_prev[15] = 26'b00000000010011100011011011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 25 timeout!");
                $fdisplay(fd_cycles, "Test Vector  25: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  25: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 25");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 26
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000101001100100001;
        x_t[1] = 26'b00000000001100011001010010;
        x_t[2] = 26'b00000000000111000101010011;
        x_t[3] = 26'b00000000001011000001100111;
        x_t[4] = 26'b00000000000100111111011110;
        x_t[5] = 26'b00000000000010111101010010;
        x_t[6] = 26'b00000000000001010110101110;
        x_t[7] = 26'b00000000010000010000100001;
        x_t[8] = 26'b00000000001011011000100011;
        x_t[9] = 26'b00000000001011011000111110;
        x_t[10] = 26'b00000000001010101111010001;
        x_t[11] = 26'b00000000000111100101110100;
        x_t[12] = 26'b00000000001000100111100001;
        x_t[13] = 26'b00000000000011000111000011;
        x_t[14] = 26'b00000000010000001011101101;
        x_t[15] = 26'b00000000001101100000111100;
        x_t[16] = 26'b00000000001011001111011111;
        x_t[17] = 26'b00000000001101110100000011;
        x_t[18] = 26'b00000000001010000100000011;
        x_t[19] = 26'b00000000001010111101110001;
        x_t[20] = 26'b00000000001101000001000000;
        x_t[21] = 26'b11111111111100001100001111;
        x_t[22] = 26'b11111111111111011010001010;
        x_t[23] = 26'b00000000000001111011110110;
        x_t[24] = 26'b11111111111110000001100110;
        x_t[25] = 26'b11111111111110011101100100;
        x_t[26] = 26'b11111111111110000111011000;
        x_t[27] = 26'b11111111111101001001110010;
        x_t[28] = 26'b00000000000010111110011100;
        x_t[29] = 26'b11111111110101101001100001;
        x_t[30] = 26'b00000000000101111101100111;
        x_t[31] = 26'b00000000000001010101111111;
        x_t[32] = 26'b00000000000010111111111101;
        x_t[33] = 26'b00000000000010000111010110;
        x_t[34] = 26'b11111111111110101110000111;
        x_t[35] = 26'b11111111111010010101000100;
        x_t[36] = 26'b11111111111101101111010010;
        x_t[37] = 26'b11111111101011011010101000;
        x_t[38] = 26'b11111111111010010010001111;
        x_t[39] = 26'b00000000000000010110010111;
        x_t[40] = 26'b00000000000000100001101000;
        x_t[41] = 26'b11111111111010111001111101;
        x_t[42] = 26'b00000000000101110100111111;
        x_t[43] = 26'b11111111110111100011011100;
        x_t[44] = 26'b00000000001000111110000101;
        x_t[45] = 26'b00000000001010100111001000;
        x_t[46] = 26'b00000000001001001011111110;
        x_t[47] = 26'b00000000001001001000000111;
        x_t[48] = 26'b00000000001010010011001111;
        x_t[49] = 26'b00000000001000011010100100;
        x_t[50] = 26'b00000000001010010011000101;
        x_t[51] = 26'b00000000001101001000000000;
        x_t[52] = 26'b00000000001100100111011000;
        x_t[53] = 26'b00000000001011011000100000;
        x_t[54] = 26'b00000000001100101011001101;
        x_t[55] = 26'b00000000001000001100010010;
        x_t[56] = 26'b00000000001001001101000101;
        x_t[57] = 26'b00000000001001001011111111;
        x_t[58] = 26'b00000000010001111100111000;
        x_t[59] = 26'b00000000001111011111101101;
        x_t[60] = 26'b00000000000111100111010011;
        x_t[61] = 26'b00000000010001010010100110;
        x_t[62] = 26'b00000000001110010010111011;
        x_t[63] = 26'b00000000000111111111100100;
        
        h_t_prev[0] = 26'b00000000000101001100100001;
        h_t_prev[1] = 26'b00000000001100011001010010;
        h_t_prev[2] = 26'b00000000000111000101010011;
        h_t_prev[3] = 26'b00000000001011000001100111;
        h_t_prev[4] = 26'b00000000000100111111011110;
        h_t_prev[5] = 26'b00000000000010111101010010;
        h_t_prev[6] = 26'b00000000000001010110101110;
        h_t_prev[7] = 26'b00000000010000010000100001;
        h_t_prev[8] = 26'b00000000001011011000100011;
        h_t_prev[9] = 26'b00000000001011011000111110;
        h_t_prev[10] = 26'b00000000001010101111010001;
        h_t_prev[11] = 26'b00000000000111100101110100;
        h_t_prev[12] = 26'b00000000001000100111100001;
        h_t_prev[13] = 26'b00000000000011000111000011;
        h_t_prev[14] = 26'b00000000010000001011101101;
        h_t_prev[15] = 26'b00000000001101100000111100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 26 timeout!");
                $fdisplay(fd_cycles, "Test Vector  26: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  26: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 26");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 27
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111111100110111110010;
        x_t[1] = 26'b00000000000010111010011001;
        x_t[2] = 26'b00000000000000011010000000;
        x_t[3] = 26'b00000000000100101011100011;
        x_t[4] = 26'b11111111111111111100001001;
        x_t[5] = 26'b11111111111111001001001101;
        x_t[6] = 26'b00000000000000100100111011;
        x_t[7] = 26'b00000000000010010000110000;
        x_t[8] = 26'b11111111111111011101010001;
        x_t[9] = 26'b00000000000011110111111010;
        x_t[10] = 26'b00000000000100010100010100;
        x_t[11] = 26'b00000000000000010000111111;
        x_t[12] = 26'b00000000000010110000111010;
        x_t[13] = 26'b00000000000001011010000010;
        x_t[14] = 26'b00000000000010101010110110;
        x_t[15] = 26'b00000000000100100111011000;
        x_t[16] = 26'b00000000000011110011101000;
        x_t[17] = 26'b00000000000111010101100000;
        x_t[18] = 26'b00000000000011001001010011;
        x_t[19] = 26'b00000000000100011100011001;
        x_t[20] = 26'b00000000001001011111110000;
        x_t[21] = 26'b11111111111110110010000000;
        x_t[22] = 26'b00000000000010001011110110;
        x_t[23] = 26'b00000000000101001100101011;
        x_t[24] = 26'b00000000000000101100000111;
        x_t[25] = 26'b00000000000000100110010100;
        x_t[26] = 26'b11111111111101100101100110;
        x_t[27] = 26'b11111111111110011000011001;
        x_t[28] = 26'b00000000000110000111111101;
        x_t[29] = 26'b11111111111101011100101010;
        x_t[30] = 26'b00000000000110001101001111;
        x_t[31] = 26'b00000000000000110010100000;
        x_t[32] = 26'b00000000000000001010001111;
        x_t[33] = 26'b11111111111111110011010101;
        x_t[34] = 26'b11111111111100010101101100;
        x_t[35] = 26'b11111111111001000110000111;
        x_t[36] = 26'b11111111111111010010101011;
        x_t[37] = 26'b11111111101111101111110110;
        x_t[38] = 26'b00000000000010001010011110;
        x_t[39] = 26'b00000000000011100100001001;
        x_t[40] = 26'b00000000001010101101110011;
        x_t[41] = 26'b11111111110111011011011011;
        x_t[42] = 26'b00000000001000110010101110;
        x_t[43] = 26'b11111111111010010010111111;
        x_t[44] = 26'b00000000001000100111101111;
        x_t[45] = 26'b00000000010001110111011010;
        x_t[46] = 26'b00000000000111111001000101;
        x_t[47] = 26'b00000000000111111000100010;
        x_t[48] = 26'b00000000001010100110010011;
        x_t[49] = 26'b00000000001000001000000010;
        x_t[50] = 26'b00000000000111010101000001;
        x_t[51] = 26'b00000000001001100000001011;
        x_t[52] = 26'b00000000001000110001110101;
        x_t[53] = 26'b00000000001000111100100111;
        x_t[54] = 26'b00000000001110111011000010;
        x_t[55] = 26'b00000000001000101110110100;
        x_t[56] = 26'b00000000001011010110100100;
        x_t[57] = 26'b00000000001000011000110101;
        x_t[58] = 26'b00000000001110011010000100;
        x_t[59] = 26'b00000000001110000000111110;
        x_t[60] = 26'b00000000000100101111010010;
        x_t[61] = 26'b00000000001101001001101111;
        x_t[62] = 26'b00000000001000101111110110;
        x_t[63] = 26'b00000000000100001001001000;
        
        h_t_prev[0] = 26'b11111111111100110111110010;
        h_t_prev[1] = 26'b00000000000010111010011001;
        h_t_prev[2] = 26'b00000000000000011010000000;
        h_t_prev[3] = 26'b00000000000100101011100011;
        h_t_prev[4] = 26'b11111111111111111100001001;
        h_t_prev[5] = 26'b11111111111111001001001101;
        h_t_prev[6] = 26'b00000000000000100100111011;
        h_t_prev[7] = 26'b00000000000010010000110000;
        h_t_prev[8] = 26'b11111111111111011101010001;
        h_t_prev[9] = 26'b00000000000011110111111010;
        h_t_prev[10] = 26'b00000000000100010100010100;
        h_t_prev[11] = 26'b00000000000000010000111111;
        h_t_prev[12] = 26'b00000000000010110000111010;
        h_t_prev[13] = 26'b00000000000001011010000010;
        h_t_prev[14] = 26'b00000000000010101010110110;
        h_t_prev[15] = 26'b00000000000100100111011000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 27 timeout!");
                $fdisplay(fd_cycles, "Test Vector  27: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  27: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 27");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 28
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000100010001010101;
        x_t[1] = 26'b00000000000100011100010001;
        x_t[2] = 26'b11111111111111001100010011;
        x_t[3] = 26'b00000000000000011100110110;
        x_t[4] = 26'b11111111111011110101011100;
        x_t[5] = 26'b11111111111011010101001001;
        x_t[6] = 26'b11111111111110001111100100;
        x_t[7] = 26'b00000000001100000111110111;
        x_t[8] = 26'b00000000000011000000001100;
        x_t[9] = 26'b00000000000100100000000000;
        x_t[10] = 26'b00000000000100010100010100;
        x_t[11] = 26'b11111111111101011001100010;
        x_t[12] = 26'b11111111111110010111111101;
        x_t[13] = 26'b11111111111100010010111100;
        x_t[14] = 26'b00000000001001010000101110;
        x_t[15] = 26'b00000000001000011011011110;
        x_t[16] = 26'b00000000000101111110011011;
        x_t[17] = 26'b00000000000111101001010000;
        x_t[18] = 26'b11111111111111110110011101;
        x_t[19] = 26'b11111111111111010010111001;
        x_t[20] = 26'b00000000000100110011011011;
        x_t[21] = 26'b00000000000010011010000101;
        x_t[22] = 26'b00000000000101001010001111;
        x_t[23] = 26'b00000000000110110101000110;
        x_t[24] = 26'b00000000000101010000011010;
        x_t[25] = 26'b00000000000101010000101011;
        x_t[26] = 26'b11111111111011101111010100;
        x_t[27] = 26'b11111111111100111010000011;
        x_t[28] = 26'b00000000000011110000110100;
        x_t[29] = 26'b00000000000001000101100101;
        x_t[30] = 26'b00000000001010100110001110;
        x_t[31] = 26'b11111111111101001011110110;
        x_t[32] = 26'b11111111111100110000001011;
        x_t[33] = 26'b11111111111100010101010011;
        x_t[34] = 26'b11111111111000110001000100;
        x_t[35] = 26'b11111111110110000000101111;
        x_t[36] = 26'b11111111111010111100010111;
        x_t[37] = 26'b11111111101110001110000000;
        x_t[38] = 26'b00000000000111110101100010;
        x_t[39] = 26'b11111111111010110101100110;
        x_t[40] = 26'b00000000001101000101111110;
        x_t[41] = 26'b11111111110001110001110010;
        x_t[42] = 26'b00000000000111010011110111;
        x_t[43] = 26'b00000000001100001000000001;
        x_t[44] = 26'b00000000001011000100001001;
        x_t[45] = 26'b00000000001000001100011000;
        x_t[46] = 26'b00000000001010110011100110;
        x_t[47] = 26'b00000000001010000011110010;
        x_t[48] = 26'b00000000001010010011001111;
        x_t[49] = 26'b00000000000111010000011011;
        x_t[50] = 26'b00000000000010010001111100;
        x_t[51] = 26'b00000000000001010110100101;
        x_t[52] = 26'b11111111111110110111011111;
        x_t[53] = 26'b11111111111110100000100010;
        x_t[54] = 26'b00000000000100110011110011;
        x_t[55] = 26'b00000000001011001010001100;
        x_t[56] = 26'b00000000001100101100100000;
        x_t[57] = 26'b00000000000100011001000011;
        x_t[58] = 26'b00000000000100010100100000;
        x_t[59] = 26'b00000000000100001001011010;
        x_t[60] = 26'b00000000000101001101111100;
        x_t[61] = 26'b00000000001011000101010100;
        x_t[62] = 26'b00000000000100110100010110;
        x_t[63] = 26'b00000000000100101100010101;
        
        h_t_prev[0] = 26'b00000000000100010001010101;
        h_t_prev[1] = 26'b00000000000100011100010001;
        h_t_prev[2] = 26'b11111111111111001100010011;
        h_t_prev[3] = 26'b00000000000000011100110110;
        h_t_prev[4] = 26'b11111111111011110101011100;
        h_t_prev[5] = 26'b11111111111011010101001001;
        h_t_prev[6] = 26'b11111111111110001111100100;
        h_t_prev[7] = 26'b00000000001100000111110111;
        h_t_prev[8] = 26'b00000000000011000000001100;
        h_t_prev[9] = 26'b00000000000100100000000000;
        h_t_prev[10] = 26'b00000000000100010100010100;
        h_t_prev[11] = 26'b11111111111101011001100010;
        h_t_prev[12] = 26'b11111111111110010111111101;
        h_t_prev[13] = 26'b11111111111100010010111100;
        h_t_prev[14] = 26'b00000000001001010000101110;
        h_t_prev[15] = 26'b00000000001000011011011110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 28 timeout!");
                $fdisplay(fd_cycles, "Test Vector  28: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  28: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 28");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 29
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000101001100100001;
        x_t[1] = 26'b00000000000101000011011011;
        x_t[2] = 26'b11111111111101101011001100;
        x_t[3] = 26'b11111111111110010101100000;
        x_t[4] = 26'b11111111111000000010111100;
        x_t[5] = 26'b11111111110100011001011000;
        x_t[6] = 26'b11111111111000000001010000;
        x_t[7] = 26'b00000000001101101101101010;
        x_t[8] = 26'b00000000000110100011000111;
        x_t[9] = 26'b00000000000100001011111101;
        x_t[10] = 26'b00000000000001100100001011;
        x_t[11] = 26'b11111111111100110000110001;
        x_t[12] = 26'b11111111111000001001111100;
        x_t[13] = 26'b11111111110101000011100100;
        x_t[14] = 26'b00000000001011001111010011;
        x_t[15] = 26'b00000000001000000111001000;
        x_t[16] = 26'b00000000000101010110110001;
        x_t[17] = 26'b00000000000101001011010101;
        x_t[18] = 26'b11111111111011100100010111;
        x_t[19] = 26'b11111111111001000111011111;
        x_t[20] = 26'b11111111111100100101110110;
        x_t[21] = 26'b00000000000000101011100100;
        x_t[22] = 26'b00000000000011011000000000;
        x_t[23] = 26'b00000000000100010010101011;
        x_t[24] = 26'b00000000000100010011100001;
        x_t[25] = 26'b00000000000100010010100001;
        x_t[26] = 26'b11111111111101000011110011;
        x_t[27] = 26'b11111111111011111011001011;
        x_t[28] = 26'b00000000000001011001101011;
        x_t[29] = 26'b00000000000011011011010101;
        x_t[30] = 26'b00000000001001011000001011;
        x_t[31] = 26'b11111111111111011001110011;
        x_t[32] = 26'b11111111111111010011101110;
        x_t[33] = 26'b00000000000000000101110101;
        x_t[34] = 26'b11111111111011101111100101;
        x_t[35] = 26'b11111111110111100011011011;
        x_t[36] = 26'b11111111111011111000000000;
        x_t[37] = 26'b11111111101101111101101101;
        x_t[38] = 26'b00000000001001011010011000;
        x_t[39] = 26'b11111111111011010011000000;
        x_t[40] = 26'b00000000001110011100111011;
        x_t[41] = 26'b00000000000010010010111000;
        x_t[42] = 26'b00000000010101110000110011;
        x_t[43] = 26'b11111111111101000010100010;
        x_t[44] = 26'b00000000010010011001010110;
        x_t[45] = 26'b00000000000001111010000000;
        x_t[46] = 26'b00000000010000111101010100;
        x_t[47] = 26'b00000000001101011110100111;
        x_t[48] = 26'b00000000001100111110110001;
        x_t[49] = 26'b00000000001001010010001010;
        x_t[50] = 26'b00000000000100111100111111;
        x_t[51] = 26'b00000000000000001001010011;
        x_t[52] = 26'b11111111111110001110100100;
        x_t[53] = 26'b11111111111011101110011000;
        x_t[54] = 26'b00000000000000010100001001;
        x_t[55] = 26'b00000000010000010010001100;
        x_t[56] = 26'b00000000010000101110010011;
        x_t[57] = 26'b00000000000100111011001010;
        x_t[58] = 26'b11111111111110110111100011;
        x_t[59] = 26'b11111111111111111101000000;
        x_t[60] = 26'b00000000001000110011111110;
        x_t[61] = 26'b00000000001010110100110000;
        x_t[62] = 26'b00000000000000101010000010;
        x_t[63] = 26'b00000000000101110010110000;
        
        h_t_prev[0] = 26'b00000000000101001100100001;
        h_t_prev[1] = 26'b00000000000101000011011011;
        h_t_prev[2] = 26'b11111111111101101011001100;
        h_t_prev[3] = 26'b11111111111110010101100000;
        h_t_prev[4] = 26'b11111111111000000010111100;
        h_t_prev[5] = 26'b11111111110100011001011000;
        h_t_prev[6] = 26'b11111111111000000001010000;
        h_t_prev[7] = 26'b00000000001101101101101010;
        h_t_prev[8] = 26'b00000000000110100011000111;
        h_t_prev[9] = 26'b00000000000100001011111101;
        h_t_prev[10] = 26'b00000000000001100100001011;
        h_t_prev[11] = 26'b11111111111100110000110001;
        h_t_prev[12] = 26'b11111111111000001001111100;
        h_t_prev[13] = 26'b11111111110101000011100100;
        h_t_prev[14] = 26'b00000000001011001111010011;
        h_t_prev[15] = 26'b00000000001000000111001000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 29 timeout!");
                $fdisplay(fd_cycles, "Test Vector  29: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  29: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 29");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 30
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001011111110100111;
        x_t[1] = 26'b00000000001110001110110000;
        x_t[2] = 26'b00000000000110011110011101;
        x_t[3] = 26'b00000000000111101100111011;
        x_t[4] = 26'b00000000000011011010011100;
        x_t[5] = 26'b11111111111110011100110101;
        x_t[6] = 26'b00000000000010111010010011;
        x_t[7] = 26'b00000000010110010011010110;
        x_t[8] = 26'b00000000001110100110110110;
        x_t[9] = 26'b00000000001100101001001010;
        x_t[10] = 26'b00000000001010101111010001;
        x_t[11] = 26'b00000000000100101110010111;
        x_t[12] = 26'b00000000000000001101000001;
        x_t[13] = 26'b00000000000011100010010100;
        x_t[14] = 26'b00000000010000100000110011;
        x_t[15] = 26'b00000000001110001001100111;
        x_t[16] = 26'b00000000001010111011101010;
        x_t[17] = 26'b00000000001011010110001000;
        x_t[18] = 26'b00000000000001110100111101;
        x_t[19] = 26'b11111111111101001111000101;
        x_t[20] = 26'b00000000000000111001001001;
        x_t[21] = 26'b00000000001001101010001110;
        x_t[22] = 26'b00000000001100011111111000;
        x_t[23] = 26'b00000000001011111001111100;
        x_t[24] = 26'b00000000001110001100110110;
        x_t[25] = 26'b00000000001101110011101011;
        x_t[26] = 26'b00000000000110110100111110;
        x_t[27] = 26'b00000000000101010000100110;
        x_t[28] = 26'b00000000001001110111010001;
        x_t[29] = 26'b00000000001111001000000010;
        x_t[30] = 26'b00000000010001011011010100;
        x_t[31] = 26'b00000000001000100011010011;
        x_t[32] = 26'b00000000001001001111101111;
        x_t[33] = 26'b00000000001001111010111011;
        x_t[34] = 26'b00000000000110001010011010;
        x_t[35] = 26'b00000000000001101110110001;
        x_t[36] = 26'b00000000000101001100011000;
        x_t[37] = 26'b11111111110101100110111011;
        x_t[38] = 26'b00000000010010001111001000;
        x_t[39] = 26'b00000000001000100111100000;
        x_t[40] = 26'b00000000010010100001110010;
        x_t[41] = 26'b00000000001000011000010100;
        x_t[42] = 26'b00000000011110101001111111;
        x_t[43] = 26'b11111111111010010010111111;
        x_t[44] = 26'b00000000010111101000100000;
        x_t[45] = 26'b11111111111101100011011011;
        x_t[46] = 26'b00000000010110001000111000;
        x_t[47] = 26'b00000000001111010101111110;
        x_t[48] = 26'b00000000001101010001110100;
        x_t[49] = 26'b00000000001000111111101000;
        x_t[50] = 26'b00000000000001111110111011;
        x_t[51] = 26'b11111111110111000101110000;
        x_t[52] = 26'b11111111110100111101001001;
        x_t[53] = 26'b11111111110000100101110000;
        x_t[54] = 26'b11111111110110001100111001;
        x_t[55] = 26'b00000000010001111001110001;
        x_t[56] = 26'b00000000010000001011111011;
        x_t[57] = 26'b11111111111101101110101111;
        x_t[58] = 26'b11111111101101101100010111;
        x_t[59] = 26'b11111111110011000111111110;
        x_t[60] = 26'b00000000001100001010101010;
        x_t[61] = 26'b00000000001000110000010101;
        x_t[62] = 26'b11111111111000000110100111;
        x_t[63] = 26'b00000000000110100111100011;
        
        h_t_prev[0] = 26'b00000000001011111110100111;
        h_t_prev[1] = 26'b00000000001110001110110000;
        h_t_prev[2] = 26'b00000000000110011110011101;
        h_t_prev[3] = 26'b00000000000111101100111011;
        h_t_prev[4] = 26'b00000000000011011010011100;
        h_t_prev[5] = 26'b11111111111110011100110101;
        h_t_prev[6] = 26'b00000000000010111010010011;
        h_t_prev[7] = 26'b00000000010110010011010110;
        h_t_prev[8] = 26'b00000000001110100110110110;
        h_t_prev[9] = 26'b00000000001100101001001010;
        h_t_prev[10] = 26'b00000000001010101111010001;
        h_t_prev[11] = 26'b00000000000100101110010111;
        h_t_prev[12] = 26'b00000000000000001101000001;
        h_t_prev[13] = 26'b00000000000011100010010100;
        h_t_prev[14] = 26'b00000000010000100000110011;
        h_t_prev[15] = 26'b00000000001110001001100111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 30 timeout!");
                $fdisplay(fd_cycles, "Test Vector  30: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  30: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 30");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 31
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001111101011011000;
        x_t[1] = 26'b00000000010000000100001101;
        x_t[2] = 26'b00000000000111000101010011;
        x_t[3] = 26'b00000000001011010100111101;
        x_t[4] = 26'b00000000000101010011101100;
        x_t[5] = 26'b11111111111111110101100101;
        x_t[6] = 26'b00000000000000001100000010;
        x_t[7] = 26'b00000000010100011001001100;
        x_t[8] = 26'b00000000001100010110011100;
        x_t[9] = 26'b00000000001010110000111001;
        x_t[10] = 26'b00000000001000111001110111;
        x_t[11] = 26'b11111111111111010011110101;
        x_t[12] = 26'b11111111111011011100101010;
        x_t[13] = 26'b11111111111000111000111000;
        x_t[14] = 26'b00000000001110110111010101;
        x_t[15] = 26'b00000000001001101100110101;
        x_t[16] = 26'b00000000000101111110011011;
        x_t[17] = 26'b00000000000100010000000111;
        x_t[18] = 26'b11111111111010100101000111;
        x_t[19] = 26'b11111111110011111101111110;
        x_t[20] = 26'b11111111110100011000010000;
        x_t[21] = 26'b00000000001010001011011000;
        x_t[22] = 26'b00000000001101000101111101;
        x_t[23] = 26'b00000000001101100010010110;
        x_t[24] = 26'b00000000001011101110100001;
        x_t[25] = 26'b00000000001011110111010110;
        x_t[26] = 26'b00000000000101110001011001;
        x_t[27] = 26'b00000000000101000000111000;
        x_t[28] = 26'b00000000001001011110000101;
        x_t[29] = 26'b00000000001011011111000111;
        x_t[30] = 26'b00000000001100100011000111;
        x_t[31] = 26'b00000000000101001110011001;
        x_t[32] = 26'b00000000000110101100001100;
        x_t[33] = 26'b00000000000111000001111001;
        x_t[34] = 26'b00000000000100000101000011;
        x_t[35] = 26'b11111111111110111101001000;
        x_t[36] = 26'b00000000000010000101100110;
        x_t[37] = 26'b11111111110000110001000101;
        x_t[38] = 26'b00000000001010000010101110;
        x_t[39] = 26'b11111111111111011011100100;
        x_t[40] = 26'b00000000010001001010110101;
        x_t[41] = 26'b11111111101100001000001001;
        x_t[42] = 26'b00000000010100010001111011;
        x_t[43] = 26'b00000000001010000100010111;
        x_t[44] = 26'b00000000010101001100000110;
        x_t[45] = 26'b11111111110101010101010000;
        x_t[46] = 26'b00000000010100001100100010;
        x_t[47] = 26'b00000000001001001000000111;
        x_t[48] = 26'b00000000000100000011000000;
        x_t[49] = 26'b00000000000000010011101000;
        x_t[50] = 26'b11111111110111010010101111;
        x_t[51] = 26'b11111111101010101101101101;
        x_t[52] = 26'b11111111101000001010101001;
        x_t[53] = 26'b11111111100101110011011010;
        x_t[54] = 26'b11111111101111011101011010;
        x_t[55] = 26'b00000000001101100101100011;
        x_t[56] = 26'b00000000001010100011000001;
        x_t[57] = 26'b11111111110100111100000001;
        x_t[58] = 26'b11111111100001011011001111;
        x_t[59] = 26'b11111111101011111110000101;
        x_t[60] = 26'b00000000001010101110101001;
        x_t[61] = 26'b00000000000010010010011111;
        x_t[62] = 26'b11111111101101000000011101;
        x_t[63] = 26'b00000000000110100111100011;
        
        h_t_prev[0] = 26'b00000000001111101011011000;
        h_t_prev[1] = 26'b00000000010000000100001101;
        h_t_prev[2] = 26'b00000000000111000101010011;
        h_t_prev[3] = 26'b00000000001011010100111101;
        h_t_prev[4] = 26'b00000000000101010011101100;
        h_t_prev[5] = 26'b11111111111111110101100101;
        h_t_prev[6] = 26'b00000000000000001100000010;
        h_t_prev[7] = 26'b00000000010100011001001100;
        h_t_prev[8] = 26'b00000000001100010110011100;
        h_t_prev[9] = 26'b00000000001010110000111001;
        h_t_prev[10] = 26'b00000000001000111001110111;
        h_t_prev[11] = 26'b11111111111111010011110101;
        h_t_prev[12] = 26'b11111111111011011100101010;
        h_t_prev[13] = 26'b11111111111000111000111000;
        h_t_prev[14] = 26'b00000000001110110111010101;
        h_t_prev[15] = 26'b00000000001001101100110101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 31 timeout!");
                $fdisplay(fd_cycles, "Test Vector  31: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  31: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 31");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 32
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000110000111101110;
        x_t[1] = 26'b00000000001010010000001111;
        x_t[2] = 26'b11111111111111001100010011;
        x_t[3] = 26'b00000000001001001101100110;
        x_t[4] = 26'b00000000000011000110001110;
        x_t[5] = 26'b11111111111100000001100001;
        x_t[6] = 26'b11111111111101011101110001;
        x_t[7] = 26'b00000000001110010110011000;
        x_t[8] = 26'b00000000000111001100011000;
        x_t[9] = 26'b00000000000110011000010001;
        x_t[10] = 26'b00000000000100010100010100;
        x_t[11] = 26'b11111111111101011001100010;
        x_t[12] = 26'b11111111111100001011011111;
        x_t[13] = 26'b11111111110110010101010110;
        x_t[14] = 26'b00000000001011001111010011;
        x_t[15] = 26'b00000000000101010000000011;
        x_t[16] = 26'b00000000000001000001001011;
        x_t[17] = 26'b11111111111111010100010001;
        x_t[18] = 26'b11111111111000100110100111;
        x_t[19] = 26'b11111111110110000001110001;
        x_t[20] = 26'b11111111110111100000011111;
        x_t[21] = 26'b00000000000100001000100101;
        x_t[22] = 26'b00000000001000001000101000;
        x_t[23] = 26'b00000000001001101110101110;
        x_t[24] = 26'b00000000000110110001110110;
        x_t[25] = 26'b00000000000111000000100100;
        x_t[26] = 26'b00000000000010010101101111;
        x_t[27] = 26'b00000000000000110101100111;
        x_t[28] = 26'b00000000000110100001001010;
        x_t[29] = 26'b00000000000010011000110010;
        x_t[30] = 26'b00000000000111101010111001;
        x_t[31] = 26'b00000000000100000111011011;
        x_t[32] = 26'b00000000000100111111001010;
        x_t[33] = 26'b00000000000111000001111001;
        x_t[34] = 26'b00000000000010010010101111;
        x_t[35] = 26'b11111111111100001011011111;
        x_t[36] = 26'b00000000000001011101110101;
        x_t[37] = 26'b11111111101110001110000000;
        x_t[38] = 26'b11111111111111010100111101;
        x_t[39] = 26'b00000000000011000110101111;
        x_t[40] = 26'b00000000001001101100100101;
        x_t[41] = 26'b11111111110110000111111110;
        x_t[42] = 26'b00000000001100110111100110;
        x_t[43] = 26'b11111111111000001111010101;
        x_t[44] = 26'b00000000001011110000110101;
        x_t[45] = 26'b11111111111110100001010101;
        x_t[46] = 26'b00000000001011110001110000;
        x_t[47] = 26'b00000000000110101000111110;
        x_t[48] = 26'b00000000000100000011000000;
        x_t[49] = 26'b11111111111101000111110000;
        x_t[50] = 26'b11111111110110111111101111;
        x_t[51] = 26'b11111111101101011011100100;
        x_t[52] = 26'b11111111101100010100101010;
        x_t[53] = 26'b11111111101010101011001011;
        x_t[54] = 26'b11111111110001101101001111;
        x_t[55] = 26'b00000000001010111000111011;
        x_t[56] = 26'b00000000000111100101111101;
        x_t[57] = 26'b11111111110010100010100011;
        x_t[58] = 26'b11111111100100011011001010;
        x_t[59] = 26'b11111111101100011101101010;
        x_t[60] = 26'b00000000000111010111111101;
        x_t[61] = 26'b11111111111100000101001100;
        x_t[62] = 26'b11111111100110111111110010;
        x_t[63] = 26'b00000000000101100001001001;
        
        h_t_prev[0] = 26'b00000000000110000111101110;
        h_t_prev[1] = 26'b00000000001010010000001111;
        h_t_prev[2] = 26'b11111111111111001100010011;
        h_t_prev[3] = 26'b00000000001001001101100110;
        h_t_prev[4] = 26'b00000000000011000110001110;
        h_t_prev[5] = 26'b11111111111100000001100001;
        h_t_prev[6] = 26'b11111111111101011101110001;
        h_t_prev[7] = 26'b00000000001110010110011000;
        h_t_prev[8] = 26'b00000000000111001100011000;
        h_t_prev[9] = 26'b00000000000110011000010001;
        h_t_prev[10] = 26'b00000000000100010100010100;
        h_t_prev[11] = 26'b11111111111101011001100010;
        h_t_prev[12] = 26'b11111111111100001011011111;
        h_t_prev[13] = 26'b11111111110110010101010110;
        h_t_prev[14] = 26'b00000000001011001111010011;
        h_t_prev[15] = 26'b00000000000101010000000011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 32 timeout!");
                $fdisplay(fd_cycles, "Test Vector  32: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  32: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 32");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 33
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111111010101101101011;
        x_t[1] = 26'b11111111111010010110001110;
        x_t[2] = 26'b11111111111000001101100101;
        x_t[3] = 26'b11111111111000100110000111;
        x_t[4] = 26'b11111111110101110101011111;
        x_t[5] = 26'b11111111101101110011110011;
        x_t[6] = 26'b11111111101011111101100010;
        x_t[7] = 26'b11111111111110011100011100;
        x_t[8] = 26'b11111111111000010111011011;
        x_t[9] = 26'b11111111110110011010000000;
        x_t[10] = 26'b11111111110101111100100010;
        x_t[11] = 26'b11111111110010100100100000;
        x_t[12] = 26'b11111111101110010001110011;
        x_t[13] = 26'b11111111100100000001010010;
        x_t[14] = 26'b11111111111110101101101110;
        x_t[15] = 26'b11111111111001011111011011;
        x_t[16] = 26'b11111111110111000110101101;
        x_t[17] = 26'b11111111110100100001011000;
        x_t[18] = 26'b11111111110100101001100111;
        x_t[19] = 26'b11111111110010100110000111;
        x_t[20] = 26'b11111111110000011101111111;
        x_t[21] = 26'b11111111111010111110111000;
        x_t[22] = 26'b11111111110101000110001000;
        x_t[23] = 26'b11111111111000101100001010;
        x_t[24] = 26'b11111111111010100110011000;
        x_t[25] = 26'b11111111111011001010001110;
        x_t[26] = 26'b11111111110011000001101110;
        x_t[27] = 26'b11111111110101000010111101;
        x_t[28] = 26'b11111111110101001100110010;
        x_t[29] = 26'b11111111111011010111100011;
        x_t[30] = 26'b11111111110100101001010001;
        x_t[31] = 26'b11111111111010111101111010;
        x_t[32] = 26'b11111111111000011111100110;
        x_t[33] = 26'b11111111110100100001101111;
        x_t[34] = 26'b11111111110001100111110100;
        x_t[35] = 26'b11111111101110111010110001;
        x_t[36] = 26'b11111111101110001101010100;
        x_t[37] = 26'b11111111100001011110101000;
        x_t[38] = 26'b11111111111000101101011000;
        x_t[39] = 26'b11111111100011011010011000;
        x_t[40] = 26'b11111111111000000010001010;
        x_t[41] = 26'b11111111101010011000111000;
        x_t[42] = 26'b11111111111110000010111100;
        x_t[43] = 26'b11111111111010111110111000;
        x_t[44] = 26'b11111111101110000101101001;
        x_t[45] = 26'b11111111101100001001001010;
        x_t[46] = 26'b11111111111110110100110111;
        x_t[47] = 26'b11111111111100000100100110;
        x_t[48] = 26'b11111111111001100111111100;
        x_t[49] = 26'b11111111111101000111110000;
        x_t[50] = 26'b11111111111000011110110001;
        x_t[51] = 26'b11111111111001001100111111;
        x_t[52] = 26'b11111111111001000111001010;
        x_t[53] = 26'b11111111110100000100011101;
        x_t[54] = 26'b11111111110010000101001101;
        x_t[55] = 26'b11111111111011110010001011;
        x_t[56] = 26'b11111111111110111111111111;
        x_t[57] = 26'b11111111111111000100000000;
        x_t[58] = 26'b00000000000000110001101100;
        x_t[59] = 26'b00000000000000101100010111;
        x_t[60] = 26'b11111111111010111010100011;
        x_t[61] = 26'b11111111110110111010000111;
        x_t[62] = 26'b11111111111010001011110001;
        x_t[63] = 26'b11111111110000010101101111;
        
        h_t_prev[0] = 26'b11111111111010101101101011;
        h_t_prev[1] = 26'b11111111111010010110001110;
        h_t_prev[2] = 26'b11111111111000001101100101;
        h_t_prev[3] = 26'b11111111111000100110000111;
        h_t_prev[4] = 26'b11111111110101110101011111;
        h_t_prev[5] = 26'b11111111101101110011110011;
        h_t_prev[6] = 26'b11111111101011111101100010;
        h_t_prev[7] = 26'b11111111111110011100011100;
        h_t_prev[8] = 26'b11111111111000010111011011;
        h_t_prev[9] = 26'b11111111110110011010000000;
        h_t_prev[10] = 26'b11111111110101111100100010;
        h_t_prev[11] = 26'b11111111110010100100100000;
        h_t_prev[12] = 26'b11111111101110010001110011;
        h_t_prev[13] = 26'b11111111100100000001010010;
        h_t_prev[14] = 26'b11111111111110101101101110;
        h_t_prev[15] = 26'b11111111111001011111011011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 33 timeout!");
                $fdisplay(fd_cycles, "Test Vector  33: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  33: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 33");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 34
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111110001110001011110;
        x_t[1] = 26'b11111111110001110010000100;
        x_t[2] = 26'b11111111101111011010010011;
        x_t[3] = 26'b11111111101110101000000001;
        x_t[4] = 26'b11111111101101101000000101;
        x_t[5] = 26'b11111111100111100100011010;
        x_t[6] = 26'b11111111100111101011101101;
        x_t[7] = 26'b11111111111010101000001001;
        x_t[8] = 26'b11111111110011110110101000;
        x_t[9] = 26'b11111111110001000101001111;
        x_t[10] = 26'b11111111110001000011011010;
        x_t[11] = 26'b11111111110000000001011011;
        x_t[12] = 26'b11111111101111000000101000;
        x_t[13] = 26'b11111111101000101101000111;
        x_t[14] = 26'b11111111111011000101101100;
        x_t[15] = 26'b11111111110110111100101100;
        x_t[16] = 26'b11111111110100010100010000;
        x_t[17] = 26'b11111111110010010111001100;
        x_t[18] = 26'b11111111110100111110101100;
        x_t[19] = 26'b11111111110110010111101111;
        x_t[20] = 26'b11111111110101001010010100;
        x_t[21] = 26'b11111111110100111100000110;
        x_t[22] = 26'b11111111101111010110000011;
        x_t[23] = 26'b11111111110010111000111010;
        x_t[24] = 26'b11111111110101010001010110;
        x_t[25] = 26'b11111111110101100001101101;
        x_t[26] = 26'b11111111101011000110110100;
        x_t[27] = 26'b11111111101101011011100101;
        x_t[28] = 26'b11111111101111000110010110;
        x_t[29] = 26'b11111111110100000101101100;
        x_t[30] = 26'b11111111101101000101010101;
        x_t[31] = 26'b11111111110011110000100110;
        x_t[32] = 26'b11111111101111111110011011;
        x_t[33] = 26'b11111111101100001001001010;
        x_t[34] = 26'b11111111101001010010010110;
        x_t[35] = 26'b11111111100110100101110110;
        x_t[36] = 26'b11111111100111010111111101;
        x_t[37] = 26'b11111111100001111111010000;
        x_t[38] = 26'b11111111110001011101011111;
        x_t[39] = 26'b11111111100110001010110000;
        x_t[40] = 26'b11111111110001111010110111;
        x_t[41] = 26'b11111111110011000101001111;
        x_t[42] = 26'b11111111110000010101011100;
        x_t[43] = 26'b11111111100101000010100001;
        x_t[44] = 26'b11111111100111011101000111;
        x_t[45] = 26'b11111111110100010111010110;
        x_t[46] = 26'b11111111111000111111110111;
        x_t[47] = 26'b11111111111011110000101101;
        x_t[48] = 26'b11111111111100010011011110;
        x_t[49] = 26'b00000000000001110000010011;
        x_t[50] = 26'b11111111111100101000110101;
        x_t[51] = 26'b11111111111111100010101011;
        x_t[52] = 26'b11111111111111110100111000;
        x_t[53] = 26'b11111111111011101110011000;
        x_t[54] = 26'b11111111111010101100100100;
        x_t[55] = 26'b11111111111110110000000100;
        x_t[56] = 26'b00000000000011000001110010;
        x_t[57] = 26'b00000000000101101110010100;
        x_t[58] = 26'b00000000000111010100011011;
        x_t[59] = 26'b00000000001000000110000010;
        x_t[60] = 26'b11111111111101000100100100;
        x_t[61] = 26'b11111111111011010011100010;
        x_t[62] = 26'b00000000000000101010000010;
        x_t[63] = 26'b11111111110110101010100110;
        
        h_t_prev[0] = 26'b11111111110001110001011110;
        h_t_prev[1] = 26'b11111111110001110010000100;
        h_t_prev[2] = 26'b11111111101111011010010011;
        h_t_prev[3] = 26'b11111111101110101000000001;
        h_t_prev[4] = 26'b11111111101101101000000101;
        h_t_prev[5] = 26'b11111111100111100100011010;
        h_t_prev[6] = 26'b11111111100111101011101101;
        h_t_prev[7] = 26'b11111111111010101000001001;
        h_t_prev[8] = 26'b11111111110011110110101000;
        h_t_prev[9] = 26'b11111111110001000101001111;
        h_t_prev[10] = 26'b11111111110001000011011010;
        h_t_prev[11] = 26'b11111111110000000001011011;
        h_t_prev[12] = 26'b11111111101111000000101000;
        h_t_prev[13] = 26'b11111111101000101101000111;
        h_t_prev[14] = 26'b11111111111011000101101100;
        h_t_prev[15] = 26'b11111111110110111100101100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 34 timeout!");
                $fdisplay(fd_cycles, "Test Vector  34: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  34: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 34");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 35
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111110000110110010010;
        x_t[1] = 26'b11111111110000010000001011;
        x_t[2] = 26'b11111111101101100101110001;
        x_t[3] = 26'b11111111101110101000000001;
        x_t[4] = 26'b11111111101101101000000101;
        x_t[5] = 26'b11111111101001101001100010;
        x_t[6] = 26'b11111111100110111001111010;
        x_t[7] = 26'b11111111111000101101111111;
        x_t[8] = 26'b11111111110100001011010000;
        x_t[9] = 26'b11111111110011100101100110;
        x_t[10] = 26'b11111111110110010000000110;
        x_t[11] = 26'b11111111110111010110010000;
        x_t[12] = 26'b11111111110101001110101001;
        x_t[13] = 26'b11111111110001001110010000;
        x_t[14] = 26'b11111111110111001000100100;
        x_t[15] = 26'b11111111111000100010011001;
        x_t[16] = 26'b11111111111000101001110110;
        x_t[17] = 26'b11111111110111010011000010;
        x_t[18] = 26'b11111111111010100101000111;
        x_t[19] = 26'b11111111111101001111000101;
        x_t[20] = 26'b11111111111100001100110100;
        x_t[21] = 26'b11111111110011101110101111;
        x_t[22] = 26'b11111111101101010111000111;
        x_t[23] = 26'b11111111110001010000100000;
        x_t[24] = 26'b11111111110100001000010001;
        x_t[25] = 26'b11111111110100010111000111;
        x_t[26] = 26'b11111111101100001010011010;
        x_t[27] = 26'b11111111101101101011010011;
        x_t[28] = 26'b11111111101100101111001101;
        x_t[29] = 26'b11111111110011010011110001;
        x_t[30] = 26'b11111111101100110101101110;
        x_t[31] = 26'b11111111110111101001000000;
        x_t[32] = 26'b11111111110100001111000001;
        x_t[33] = 26'b11111111110001000011101101;
        x_t[34] = 26'b11111111101110000011001100;
        x_t[35] = 26'b11111111101011001101111010;
        x_t[36] = 26'b11111111101100000010001010;
        x_t[37] = 26'b11111111100011000000011110;
        x_t[38] = 26'b11111111110101001111100001;
        x_t[39] = 26'b11111111101101100001000110;
        x_t[40] = 26'b11111111111001101110110111;
        x_t[41] = 26'b11111111111110110100010101;
        x_t[42] = 26'b11111111111010101101100000;
        x_t[43] = 26'b11111111011101011111110010;
        x_t[44] = 26'b11111111101101101111010011;
        x_t[45] = 26'b11111111111000101101111010;
        x_t[46] = 26'b00000000000000000111110000;
        x_t[47] = 26'b00000000000010010010011101;
        x_t[48] = 26'b00000000000011011100111000;
        x_t[49] = 26'b00000000001010011100010011;
        x_t[50] = 26'b00000000000100101001111110;
        x_t[51] = 26'b00000000000101100101000010;
        x_t[52] = 26'b00000000000100111100010001;
        x_t[53] = 26'b00000000000001101000111101;
        x_t[54] = 26'b00000000000010001100000000;
        x_t[55] = 26'b00000000000111011000100000;
        x_t[56] = 26'b00000000001011111000111100;
        x_t[57] = 26'b00000000001101101101111000;
        x_t[58] = 26'b00000000001011101011100101;
        x_t[59] = 26'b00000000001110000000111110;
        x_t[60] = 26'b00000000000101001101111100;
        x_t[61] = 26'b00000000000100000110010111;
        x_t[62] = 26'b00000000001000010010010001;
        x_t[63] = 26'b00000000000001101010101101;
        
        h_t_prev[0] = 26'b11111111110000110110010010;
        h_t_prev[1] = 26'b11111111110000010000001011;
        h_t_prev[2] = 26'b11111111101101100101110001;
        h_t_prev[3] = 26'b11111111101110101000000001;
        h_t_prev[4] = 26'b11111111101101101000000101;
        h_t_prev[5] = 26'b11111111101001101001100010;
        h_t_prev[6] = 26'b11111111100110111001111010;
        h_t_prev[7] = 26'b11111111111000101101111111;
        h_t_prev[8] = 26'b11111111110100001011010000;
        h_t_prev[9] = 26'b11111111110011100101100110;
        h_t_prev[10] = 26'b11111111110110010000000110;
        h_t_prev[11] = 26'b11111111110111010110010000;
        h_t_prev[12] = 26'b11111111110101001110101001;
        h_t_prev[13] = 26'b11111111110001001110010000;
        h_t_prev[14] = 26'b11111111110111001000100100;
        h_t_prev[15] = 26'b11111111111000100010011001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 35 timeout!");
                $fdisplay(fd_cycles, "Test Vector  35: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  35: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 35");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 36
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111110110011001011100;
        x_t[1] = 26'b11111111111010101001110011;
        x_t[2] = 26'b11111111111001011011010001;
        x_t[3] = 26'b11111111111010000110110010;
        x_t[4] = 26'b11111111111001010011110010;
        x_t[5] = 26'b11111111110101110010001000;
        x_t[6] = 26'b11111111110011101111011011;
        x_t[7] = 26'b00000000000010100101000110;
        x_t[8] = 26'b11111111111111001000101001;
        x_t[9] = 26'b11111111111111001011001111;
        x_t[10] = 26'b00000000000010001011010100;
        x_t[11] = 26'b00000000000010110100000011;
        x_t[12] = 26'b11111111111111011110001100;
        x_t[13] = 26'b11111111111001101111011001;
        x_t[14] = 26'b00000000000011111111001110;
        x_t[15] = 26'b00000000000011111110101100;
        x_t[16] = 26'b00000000000100000111011101;
        x_t[17] = 26'b00000000000010101101011010;
        x_t[18] = 26'b00000000000101000111110011;
        x_t[19] = 26'b00000000000101110100010001;
        x_t[20] = 26'b00000000000100011010011001;
        x_t[21] = 26'b11111111111001100110011110;
        x_t[22] = 26'b11111111110011101101010010;
        x_t[23] = 26'b11111111110101110010100010;
        x_t[24] = 26'b11111111111001101001011110;
        x_t[25] = 26'b11111111111010001100000100;
        x_t[26] = 26'b11111111110110001100011111;
        x_t[27] = 26'b11111111110110100001010010;
        x_t[28] = 26'b11111111110010110101101001;
        x_t[29] = 26'b11111111111000110001001011;
        x_t[30] = 26'b11111111110100001010000010;
        x_t[31] = 26'b00000000000000110010100000;
        x_t[32] = 26'b11111111111111010011101110;
        x_t[33] = 26'b11111111111011110000010011;
        x_t[34] = 26'b11111111110111110111111010;
        x_t[35] = 26'b11111111110110111011111100;
        x_t[36] = 26'b11111111110111100001101100;
        x_t[37] = 26'b11111111101001011000001010;
        x_t[38] = 26'b11111111111111101001000111;
        x_t[39] = 26'b11111111110011111100101010;
        x_t[40] = 26'b00000000000011001111100011;
        x_t[41] = 26'b11111111111101111100101100;
        x_t[42] = 26'b00000000000101000101100011;
        x_t[43] = 26'b11111111111010111110111000;
        x_t[44] = 26'b11111111111000111010010010;
        x_t[45] = 26'b11111111111110100001010101;
        x_t[46] = 26'b00000000001011110001110000;
        x_t[47] = 26'b00000000001110011010010010;
        x_t[48] = 26'b00000000001110001011000000;
        x_t[49] = 26'b00000000010100010010011100;
        x_t[50] = 26'b00000000001111010110001010;
        x_t[51] = 26'b00000000001101011011010100;
        x_t[52] = 26'b00000000001011010101100001;
        x_t[53] = 26'b00000000000111001101010001;
        x_t[54] = 26'b00000000001001010011011101;
        x_t[55] = 26'b00000000010010001011000010;
        x_t[56] = 26'b00000000010110000110000010;
        x_t[57] = 26'b00000000010111010011110001;
        x_t[58] = 26'b00000000010000110111000101;
        x_t[59] = 26'b00000000010001101101110100;
        x_t[60] = 26'b00000000010001011100000001;
        x_t[61] = 26'b00000000010000100000111100;
        x_t[62] = 26'b00000000010000100110111000;
        x_t[63] = 26'b00000000001111001001001111;
        
        h_t_prev[0] = 26'b11111111110110011001011100;
        h_t_prev[1] = 26'b11111111111010101001110011;
        h_t_prev[2] = 26'b11111111111001011011010001;
        h_t_prev[3] = 26'b11111111111010000110110010;
        h_t_prev[4] = 26'b11111111111001010011110010;
        h_t_prev[5] = 26'b11111111110101110010001000;
        h_t_prev[6] = 26'b11111111110011101111011011;
        h_t_prev[7] = 26'b00000000000010100101000110;
        h_t_prev[8] = 26'b11111111111111001000101001;
        h_t_prev[9] = 26'b11111111111111001011001111;
        h_t_prev[10] = 26'b00000000000010001011010100;
        h_t_prev[11] = 26'b00000000000010110100000011;
        h_t_prev[12] = 26'b11111111111111011110001100;
        h_t_prev[13] = 26'b11111111111001101111011001;
        h_t_prev[14] = 26'b00000000000011111111001110;
        h_t_prev[15] = 26'b00000000000011111110101100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 36 timeout!");
                $fdisplay(fd_cycles, "Test Vector  36: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  36: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 36");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 37
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111111110000110101101;
        x_t[1] = 26'b00000000000010111010011001;
        x_t[2] = 26'b11111111111111011111101111;
        x_t[3] = 26'b11111111111110000010001010;
        x_t[4] = 26'b11111111111100001001101010;
        x_t[5] = 26'b11111111111000100011101000;
        x_t[6] = 26'b11111111110111101000010111;
        x_t[7] = 26'b00000000001011110011100000;
        x_t[8] = 26'b00000000000101100101001110;
        x_t[9] = 26'b00000000000100001011111101;
        x_t[10] = 26'b00000000000100111011011101;
        x_t[11] = 26'b00000000000000111001110000;
        x_t[12] = 26'b11111111111110101111011000;
        x_t[13] = 26'b11111111110011010110100011;
        x_t[14] = 26'b00000000001011100100011001;
        x_t[15] = 26'b00000000001001101100110101;
        x_t[16] = 26'b00000000000111110101011000;
        x_t[17] = 26'b00000000000101011111000100;
        x_t[18] = 26'b00000000000110011100001000;
        x_t[19] = 26'b00000000000100110010010111;
        x_t[20] = 26'b00000000000000100000000111;
        x_t[21] = 26'b11111111111001010000011000;
        x_t[22] = 26'b11111111110101010010110101;
        x_t[23] = 26'b11111111110110111000001001;
        x_t[24] = 26'b11111111111001110101101010;
        x_t[25] = 26'b11111111111010110001010111;
        x_t[26] = 26'b11111111110110011101011000;
        x_t[27] = 26'b11111111111000001111010110;
        x_t[28] = 26'b11111111110100110011100110;
        x_t[29] = 26'b11111111111111010001001000;
        x_t[30] = 26'b11111111110000101111011111;
        x_t[31] = 26'b00000000000001111001011110;
        x_t[32] = 26'b11111111111111000001100011;
        x_t[33] = 26'b11111111111010000001010010;
        x_t[34] = 26'b11111111110110101011101101;
        x_t[35] = 26'b11111111110101011001010000;
        x_t[36] = 26'b11111111111000001001011101;
        x_t[37] = 26'b11111111101001111000110010;
        x_t[38] = 26'b00000000000001110110010011;
        x_t[39] = 26'b11111111110001101001101011;
        x_t[40] = 26'b00000000000110111110101011;
        x_t[41] = 26'b11111111110100110100100001;
        x_t[42] = 26'b00000000000011100110101100;
        x_t[43] = 26'b11111111110001011000011110;
        x_t[44] = 26'b11111111111011101101000010;
        x_t[45] = 26'b11111111111010101001101110;
        x_t[46] = 26'b00000000001111010101101101;
        x_t[47] = 26'b00000000010000111001011011;
        x_t[48] = 26'b00000000010000110110100010;
        x_t[49] = 26'b00000000010101001010000010;
        x_t[50] = 26'b00000000010000001111001011;
        x_t[51] = 26'b00000000001101001000000000;
        x_t[52] = 26'b00000000001010000011101011;
        x_t[53] = 26'b00000000000011101110100101;
        x_t[54] = 26'b00000000000010001100000000;
        x_t[55] = 26'b00000000010101111100101110;
        x_t[56] = 26'b00000000011000110001111010;
        x_t[57] = 26'b00000000011010110001011100;
        x_t[58] = 26'b00000000010000000010110000;
        x_t[59] = 26'b00000000001101100001011001;
        x_t[60] = 26'b00000000011011010000101111;
        x_t[61] = 26'b00000000011000100010000110;
        x_t[62] = 26'b00000000010011011000011011;
        x_t[63] = 26'b00000000010110000001010011;
        
        h_t_prev[0] = 26'b11111111111110000110101101;
        h_t_prev[1] = 26'b00000000000010111010011001;
        h_t_prev[2] = 26'b11111111111111011111101111;
        h_t_prev[3] = 26'b11111111111110000010001010;
        h_t_prev[4] = 26'b11111111111100001001101010;
        h_t_prev[5] = 26'b11111111111000100011101000;
        h_t_prev[6] = 26'b11111111110111101000010111;
        h_t_prev[7] = 26'b00000000001011110011100000;
        h_t_prev[8] = 26'b00000000000101100101001110;
        h_t_prev[9] = 26'b00000000000100001011111101;
        h_t_prev[10] = 26'b00000000000100111011011101;
        h_t_prev[11] = 26'b00000000000000111001110000;
        h_t_prev[12] = 26'b11111111111110101111011000;
        h_t_prev[13] = 26'b11111111110011010110100011;
        h_t_prev[14] = 26'b00000000001011100100011001;
        h_t_prev[15] = 26'b00000000001001101100110101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 37 timeout!");
                $fdisplay(fd_cycles, "Test Vector  37: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  37: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 37");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 38
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000001001100000001;
        x_t[1] = 26'b00000000000000110001010110;
        x_t[2] = 26'b11111111111100011101100000;
        x_t[3] = 26'b11111111111001001100110010;
        x_t[4] = 26'b11111111110110110010000111;
        x_t[5] = 26'b11111111110100000011001100;
        x_t[6] = 26'b11111111110100100001001101;
        x_t[7] = 26'b00000000001100011100001110;
        x_t[8] = 26'b00000000000100111011111110;
        x_t[9] = 26'b00000000000001010111100011;
        x_t[10] = 26'b11111111111111101110110001;
        x_t[11] = 26'b11111111111001010000100011;
        x_t[12] = 26'b11111111111001100111100110;
        x_t[13] = 26'b11111111110001101001100001;
        x_t[14] = 26'b00000000001101111000000011;
        x_t[15] = 26'b00000000001010010101100001;
        x_t[16] = 26'b00000000000110111001111001;
        x_t[17] = 26'b00000000000011111100010111;
        x_t[18] = 26'b00000000000100001000100011;
        x_t[19] = 26'b00000000000010000010101000;
        x_t[20] = 26'b11111111111111101110000100;
        x_t[21] = 26'b11111111111010101000110010;
        x_t[22] = 26'b11111111110110010010010010;
        x_t[23] = 26'b11111111111000101100001010;
        x_t[24] = 26'b11111111111100000111110011;
        x_t[25] = 26'b11111111111100111010000111;
        x_t[26] = 26'b11111111110110011101011000;
        x_t[27] = 26'b11111111111000111110100000;
        x_t[28] = 26'b11111111110110110001100011;
        x_t[29] = 26'b00000000000011011011010101;
        x_t[30] = 26'b11111111110110010110100010;
        x_t[31] = 26'b00000000000001111001011110;
        x_t[32] = 26'b00000000000000001010001111;
        x_t[33] = 26'b11111111111011011101110011;
        x_t[34] = 26'b11111111110111010001110011;
        x_t[35] = 26'b11111111110110111011111100;
        x_t[36] = 26'b11111111111000011101010101;
        x_t[37] = 26'b11111111101010111010000001;
        x_t[38] = 26'b00000000001011111011101111;
        x_t[39] = 26'b11111111110110001111101001;
        x_t[40] = 26'b00000000001110011100111011;
        x_t[41] = 26'b00000000000011001010100000;
        x_t[42] = 26'b00000000001011110000011101;
        x_t[43] = 26'b11111111101001110101101110;
        x_t[44] = 26'b00000000000000100101110110;
        x_t[45] = 26'b11111111111010001010110001;
        x_t[46] = 26'b00000000010110110010010100;
        x_t[47] = 26'b00000000010110110011011001;
        x_t[48] = 26'b00000000010101111010100001;
        x_t[49] = 26'b00000000011001100000000011;
        x_t[50] = 26'b00000000010010100111001110;
        x_t[51] = 26'b00000000001111001111001110;
        x_t[52] = 26'b00000000001100100111011000;
        x_t[53] = 26'b00000000000101011101111011;
        x_t[54] = 26'b00000000000001110100000001;
        x_t[55] = 26'b00000000011100101100010011;
        x_t[56] = 26'b00000000011101111000011101;
        x_t[57] = 26'b00000000011111000010010010;
        x_t[58] = 26'b00000000010001101011011011;
        x_t[59] = 26'b00000000001111000000001000;
        x_t[60] = 26'b00000000100001010000000111;
        x_t[61] = 26'b00000000011100101010111101;
        x_t[62] = 26'b00000000010010111010110101;
        x_t[63] = 26'b00000000010110110110000111;
        
        h_t_prev[0] = 26'b00000000000001001100000001;
        h_t_prev[1] = 26'b00000000000000110001010110;
        h_t_prev[2] = 26'b11111111111100011101100000;
        h_t_prev[3] = 26'b11111111111001001100110010;
        h_t_prev[4] = 26'b11111111110110110010000111;
        h_t_prev[5] = 26'b11111111110100000011001100;
        h_t_prev[6] = 26'b11111111110100100001001101;
        h_t_prev[7] = 26'b00000000001100011100001110;
        h_t_prev[8] = 26'b00000000000100111011111110;
        h_t_prev[9] = 26'b00000000000001010111100011;
        h_t_prev[10] = 26'b11111111111111101110110001;
        h_t_prev[11] = 26'b11111111111001010000100011;
        h_t_prev[12] = 26'b11111111111001100111100110;
        h_t_prev[13] = 26'b11111111110001101001100001;
        h_t_prev[14] = 26'b00000000001101111000000011;
        h_t_prev[15] = 26'b00000000001010010101100001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 38 timeout!");
                $fdisplay(fd_cycles, "Test Vector  38: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  38: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 38");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 39
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001001100000110000;
        x_t[1] = 26'b00000000001001000001111100;
        x_t[2] = 26'b00000000000010110101011000;
        x_t[3] = 26'b11111111111110101000110101;
        x_t[4] = 26'b11111111111011110101011100;
        x_t[5] = 26'b11111111110111100001000100;
        x_t[6] = 26'b11111111110111001111011110;
        x_t[7] = 26'b00000000010110010011010110;
        x_t[8] = 26'b00000000001110010010001110;
        x_t[9] = 26'b00000000001001100000101101;
        x_t[10] = 26'b00000000000101100010100101;
        x_t[11] = 26'b11111111111110101011000100;
        x_t[12] = 26'b11111111111101101001001000;
        x_t[13] = 26'b11111111110110110000100110;
        x_t[14] = 26'b00000000010111110000110111;
        x_t[15] = 26'b00000000010011110111110001;
        x_t[16] = 26'b00000000001110101001100101;
        x_t[17] = 26'b00000000001001110011011011;
        x_t[18] = 26'b00000000001001000100110011;
        x_t[19] = 26'b00000000000110110110001010;
        x_t[20] = 26'b00000000000100011010011001;
        x_t[21] = 26'b11111111111101111010110000;
        x_t[22] = 26'b11111111111000101010100110;
        x_t[23] = 26'b11111111111001110001110001;
        x_t[24] = 26'b11111111111110110010010100;
        x_t[25] = 26'b11111111111111011011101110;
        x_t[26] = 26'b11111111111001101000001001;
        x_t[27] = 26'b11111111111010011100110101;
        x_t[28] = 26'b11111111110110100100111101;
        x_t[29] = 26'b00000000000110010010010110;
        x_t[30] = 26'b11111111111100011100110011;
        x_t[31] = 26'b00000000000100101010111010;
        x_t[32] = 26'b00000000000100001000101001;
        x_t[33] = 26'b11111111111111001110010101;
        x_t[34] = 26'b11111111111011001001011111;
        x_t[35] = 26'b11111111111001011001110110;
        x_t[36] = 26'b11111111110110100110000011;
        x_t[37] = 26'b11111111101000100111001111;
        x_t[38] = 26'b00000000001110001000111011;
        x_t[39] = 26'b11111111110010100100011110;
        x_t[40] = 26'b00000000001101110001011100;
        x_t[41] = 26'b11111111111001100110100000;
        x_t[42] = 26'b00000000000110111100001001;
        x_t[43] = 26'b11111111101101010001001010;
        x_t[44] = 26'b00000000000111100100101101;
        x_t[45] = 26'b11111111111100000110100101;
        x_t[46] = 26'b00000000011010111111101101;
        x_t[47] = 26'b00000000011011011101110011;
        x_t[48] = 26'b00000000011010101011011110;
        x_t[49] = 26'b00000000011110001000100101;
        x_t[50] = 26'b00000000010110011110010011;
        x_t[51] = 26'b00000000010010010000011010;
        x_t[52] = 26'b00000000010000001000011101;
        x_t[53] = 26'b00000000001001010010111001;
        x_t[54] = 26'b00000000000110101011101010;
        x_t[55] = 26'b00000000011110010011111000;
        x_t[56] = 26'b00000000011111110000110001;
        x_t[57] = 26'b00000000100000101000100110;
        x_t[58] = 26'b00000000010100001000011101;
        x_t[59] = 26'b00000000010010101100111110;
        x_t[60] = 26'b00000000100100001000001000;
        x_t[61] = 26'b00000000011110111111111100;
        x_t[62] = 26'b00000000010100100010011001;
        x_t[63] = 26'b00000000011001100110001001;
        
        h_t_prev[0] = 26'b00000000001001100000110000;
        h_t_prev[1] = 26'b00000000001001000001111100;
        h_t_prev[2] = 26'b00000000000010110101011000;
        h_t_prev[3] = 26'b11111111111110101000110101;
        h_t_prev[4] = 26'b11111111111011110101011100;
        h_t_prev[5] = 26'b11111111110111100001000100;
        h_t_prev[6] = 26'b11111111110111001111011110;
        h_t_prev[7] = 26'b00000000010110010011010110;
        h_t_prev[8] = 26'b00000000001110010010001110;
        h_t_prev[9] = 26'b00000000001001100000101101;
        h_t_prev[10] = 26'b00000000000101100010100101;
        h_t_prev[11] = 26'b11111111111110101011000100;
        h_t_prev[12] = 26'b11111111111101101001001000;
        h_t_prev[13] = 26'b11111111110110110000100110;
        h_t_prev[14] = 26'b00000000010111110000110111;
        h_t_prev[15] = 26'b00000000010011110111110001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 39 timeout!");
                $fdisplay(fd_cycles, "Test Vector  39: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  39: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 39");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 40
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000111101010011000;
        x_t[1] = 26'b00000000001001010101100001;
        x_t[2] = 26'b00000000000010110101011000;
        x_t[3] = 26'b00000000000000011100110110;
        x_t[4] = 26'b11111111111101011010011111;
        x_t[5] = 26'b11111111111000001101011100;
        x_t[6] = 26'b11111111111000000001010000;
        x_t[7] = 26'b00000000010100101101100011;
        x_t[8] = 26'b00000000001111111001010111;
        x_t[9] = 26'b00000000001010110000111001;
        x_t[10] = 26'b00000000001001110100100100;
        x_t[11] = 26'b00000000000011001000011100;
        x_t[12] = 26'b00000000000001101010101011;
        x_t[13] = 26'b11111111111001101111011001;
        x_t[14] = 26'b00000000010101011101001101;
        x_t[15] = 26'b00000000010100110100110010;
        x_t[16] = 26'b00000000010001011100000010;
        x_t[17] = 26'b00000000001100100101000101;
        x_t[18] = 26'b00000000001011011000011001;
        x_t[19] = 26'b00000000001000111001111110;
        x_t[20] = 26'b00000000000101111110100000;
        x_t[21] = 26'b11111111111011100000000010;
        x_t[22] = 26'b11111111110101101100001101;
        x_t[23] = 26'b11111111110111000011110000;
        x_t[24] = 26'b11111111111011100011010001;
        x_t[25] = 26'b11111111111100010100110100;
        x_t[26] = 26'b11111111110100111000000000;
        x_t[27] = 26'b11111111110110010001100100;
        x_t[28] = 26'b11111111110011001110110101;
        x_t[29] = 26'b00000000000001100110110111;
        x_t[30] = 26'b11111111111001010001110111;
        x_t[31] = 26'b00000000000001000100010000;
        x_t[32] = 26'b11111111111110011101001101;
        x_t[33] = 26'b11111111111001011100010001;
        x_t[34] = 26'b11111111110110011000101001;
        x_t[35] = 26'b11111111110011100010110101;
        x_t[36] = 26'b11111111110011001011011000;
        x_t[37] = 26'b11111111100110110101000110;
        x_t[38] = 26'b00000000000111100001010111;
        x_t[39] = 26'b11111111101111110100000101;
        x_t[40] = 26'b00000000000101111101011101;
        x_t[41] = 26'b11111111111010011110001001;
        x_t[42] = 26'b00000000001001111001111000;
        x_t[43] = 26'b11111111100010111110110111;
        x_t[44] = 26'b00000000000111001110010111;
        x_t[45] = 26'b11111111111000101101111010;
        x_t[46] = 26'b00000000010011110111110100;
        x_t[47] = 26'b00000000010111000111010010;
        x_t[48] = 26'b00000000010111011001110100;
        x_t[49] = 26'b00000000011100000110110110;
        x_t[50] = 26'b00000000010100101100010000;
        x_t[51] = 26'b00000000001111100010100011;
        x_t[52] = 26'b00000000001100111011110101;
        x_t[53] = 26'b00000000000110001010011101;
        x_t[54] = 26'b00000000000101111011101101;
        x_t[55] = 26'b00000000011011010101111111;
        x_t[56] = 26'b00000000011101010110000101;
        x_t[57] = 26'b00000000011101011011111110;
        x_t[58] = 26'b00000000010001001000100010;
        x_t[59] = 26'b00000000001111011111101101;
        x_t[60] = 26'b00000000100100001000001000;
        x_t[61] = 26'b00000000011111100001000011;
        x_t[62] = 26'b00000000010111010011111100;
        x_t[63] = 26'b00000000011101001010111110;
        
        h_t_prev[0] = 26'b00000000000111101010011000;
        h_t_prev[1] = 26'b00000000001001010101100001;
        h_t_prev[2] = 26'b00000000000010110101011000;
        h_t_prev[3] = 26'b00000000000000011100110110;
        h_t_prev[4] = 26'b11111111111101011010011111;
        h_t_prev[5] = 26'b11111111111000001101011100;
        h_t_prev[6] = 26'b11111111111000000001010000;
        h_t_prev[7] = 26'b00000000010100101101100011;
        h_t_prev[8] = 26'b00000000001111111001010111;
        h_t_prev[9] = 26'b00000000001010110000111001;
        h_t_prev[10] = 26'b00000000001001110100100100;
        h_t_prev[11] = 26'b00000000000011001000011100;
        h_t_prev[12] = 26'b00000000000001101010101011;
        h_t_prev[13] = 26'b11111111111001101111011001;
        h_t_prev[14] = 26'b00000000010101011101001101;
        h_t_prev[15] = 26'b00000000010100110100110010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 40 timeout!");
                $fdisplay(fd_cycles, "Test Vector  40: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  40: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 40");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 41
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000001011111110000;
        x_t[1] = 26'b00000000000100011100010001;
        x_t[2] = 26'b00000000000001000000110110;
        x_t[3] = 26'b11111111111110101000110101;
        x_t[4] = 26'b11111111111100011101110111;
        x_t[5] = 26'b11111111110110011110100000;
        x_t[6] = 26'b11111111110101101011111001;
        x_t[7] = 26'b00000000001101101101101010;
        x_t[8] = 26'b00000000001100101011000100;
        x_t[9] = 26'b00000000001010001000110011;
        x_t[10] = 26'b00000000001010011011101101;
        x_t[11] = 26'b00000000000100011001111110;
        x_t[12] = 26'b11111111111111000110110010;
        x_t[13] = 26'b11111111110010000100110001;
        x_t[14] = 26'b00000000010010011111010111;
        x_t[15] = 26'b00000000010010111010101111;
        x_t[16] = 26'b00000000001111111000111001;
        x_t[17] = 26'b00000000001010101110101001;
        x_t[18] = 26'b00000000001001011001111001;
        x_t[19] = 26'b00000000000100110010010111;
        x_t[20] = 26'b11111111111110001001111101;
        x_t[21] = 26'b11111111111100000001001100;
        x_t[22] = 26'b11111111110110011110111111;
        x_t[23] = 26'b11111111110111011010111101;
        x_t[24] = 26'b11111111111100100000001010;
        x_t[25] = 26'b11111111111101010010111110;
        x_t[26] = 26'b11111111110110101110010001;
        x_t[27] = 26'b11111111110111111111100111;
        x_t[28] = 26'b11111111110101100101111110;
        x_t[29] = 26'b00000000000010111010000011;
        x_t[30] = 26'b11111111111011011110010111;
        x_t[31] = 26'b00000000000011010010001100;
        x_t[32] = 26'b00000000000010101101110010;
        x_t[33] = 26'b11111111111110000100010100;
        x_t[34] = 26'b11111111111001111101010001;
        x_t[35] = 26'b11111111111000011110101000;
        x_t[36] = 26'b11111111110110100110000011;
        x_t[37] = 26'b11111111101101101101011001;
        x_t[38] = 26'b00000000001000001001101101;
        x_t[39] = 26'b11111111110011011111010000;
        x_t[40] = 26'b00000000001010000010010100;
        x_t[41] = 26'b11111111110100011000101100;
        x_t[42] = 26'b00000000001101100111000010;
        x_t[43] = 26'b11111111110100001000000001;
        x_t[44] = 26'b00000000000110100001101011;
        x_t[45] = 26'b11111111110110110010000110;
        x_t[46] = 26'b00000000010011001110011000;
        x_t[47] = 26'b00000000010110011111100000;
        x_t[48] = 26'b00000000010110110011101101;
        x_t[49] = 26'b00000000011010000101000111;
        x_t[50] = 26'b00000000010100000110010000;
        x_t[51] = 26'b00000000001100110100101011;
        x_t[52] = 26'b00000000001001011010110000;
        x_t[53] = 26'b00000000000001010010101100;
        x_t[54] = 26'b00000000000001110100000001;
        x_t[55] = 26'b00000000011100101100010011;
        x_t[56] = 26'b00000000011101111000011101;
        x_t[57] = 26'b00000000011011110101101001;
        x_t[58] = 26'b00000000001101010100010001;
        x_t[59] = 26'b00000000001100010010011101;
        x_t[60] = 26'b00000000100001101110110010;
        x_t[61] = 26'b00000000011100011010011010;
        x_t[62] = 26'b00000000010110110110010110;
        x_t[63] = 26'b00000000011001100110001001;
        
        h_t_prev[0] = 26'b00000000000001011111110000;
        h_t_prev[1] = 26'b00000000000100011100010001;
        h_t_prev[2] = 26'b00000000000001000000110110;
        h_t_prev[3] = 26'b11111111111110101000110101;
        h_t_prev[4] = 26'b11111111111100011101110111;
        h_t_prev[5] = 26'b11111111110110011110100000;
        h_t_prev[6] = 26'b11111111110101101011111001;
        h_t_prev[7] = 26'b00000000001101101101101010;
        h_t_prev[8] = 26'b00000000001100101011000100;
        h_t_prev[9] = 26'b00000000001010001000110011;
        h_t_prev[10] = 26'b00000000001010011011101101;
        h_t_prev[11] = 26'b00000000000100011001111110;
        h_t_prev[12] = 26'b11111111111111000110110010;
        h_t_prev[13] = 26'b11111111110010000100110001;
        h_t_prev[14] = 26'b00000000010010011111010111;
        h_t_prev[15] = 26'b00000000010010111010101111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 41 timeout!");
                $fdisplay(fd_cycles, "Test Vector  41: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  41: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 41");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 42
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001000100101100100;
        x_t[1] = 26'b00000000001110100010010101;
        x_t[2] = 26'b00000000001011010101001111;
        x_t[3] = 26'b00000000001001100000111100;
        x_t[4] = 26'b00000000000101100111111001;
        x_t[5] = 26'b11111111111101011010010001;
        x_t[6] = 26'b11111111110111101000010111;
        x_t[7] = 26'b00000000011001001010100100;
        x_t[8] = 26'b00000000010110000001010100;
        x_t[9] = 26'b00000000010011100010001000;
        x_t[10] = 26'b00000000010001001010001111;
        x_t[11] = 26'b00000000001011011010011010;
        x_t[12] = 26'b00000000000011001000010101;
        x_t[13] = 26'b11111111110001101001100001;
        x_t[14] = 26'b00000000011110000001101001;
        x_t[15] = 26'b00000000011010001110100110;
        x_t[16] = 26'b00000000010110011001010001;
        x_t[17] = 26'b00000000010000010001111101;
        x_t[18] = 26'b00000000001110101011001110;
        x_t[19] = 26'b00000000001001001111111100;
        x_t[20] = 26'b00000000000000100000000111;
        x_t[21] = 26'b11111111111100101101011001;
        x_t[22] = 26'b11111111111000000100100001;
        x_t[23] = 26'b11111111111001110001110001;
        x_t[24] = 26'b11111111111110111110100000;
        x_t[25] = 26'b00000000000000000001000001;
        x_t[26] = 26'b11111111111101000011110011;
        x_t[27] = 26'b11111111111101001001110010;
        x_t[28] = 26'b11111111111001001000101100;
        x_t[29] = 26'b00000000000111000100010001;
        x_t[30] = 26'b11111111111111110111010110;
        x_t[31] = 26'b00000000001010110001001111;
        x_t[32] = 26'b00000000001001100001111010;
        x_t[33] = 26'b00000000000101100101011000;
        x_t[34] = 26'b00000000000001101100101000;
        x_t[35] = 26'b11111111111110101001011001;
        x_t[36] = 26'b11111111111010111100010111;
        x_t[37] = 26'b11111111110000000000001010;
        x_t[38] = 26'b00000000001010010110111001;
        x_t[39] = 26'b11111111110101010100110110;
        x_t[40] = 26'b00000000001001101100100101;
        x_t[41] = 26'b11111111110011100001000011;
        x_t[42] = 26'b00000000001111011101100111;
        x_t[43] = 26'b11111111111000111011001101;
        x_t[44] = 26'b00000000001110001101001111;
        x_t[45] = 26'b00000000000000011101001001;
        x_t[46] = 26'b00000000011011101001001010;
        x_t[47] = 26'b00000000011101111100111100;
        x_t[48] = 26'b00000000011011010001100101;
        x_t[49] = 26'b00000000100000001010010100;
        x_t[50] = 26'b00000000011001011100010110;
        x_t[51] = 26'b00000000010011011101101011;
        x_t[52] = 26'b00000000010000110001011001;
        x_t[53] = 26'b00000000001000010000000101;
        x_t[54] = 26'b00000000001000100011100001;
        x_t[55] = 26'b00000000100001100011000011;
        x_t[56] = 26'b00000000100010111111000000;
        x_t[57] = 26'b00000000100000101000100110;
        x_t[58] = 26'b00000000010001011001111111;
        x_t[59] = 26'b00000000010000001111000101;
        x_t[60] = 26'b00000000100001101110110010;
        x_t[61] = 26'b00000000011100001001110110;
        x_t[62] = 26'b00000000010111110001100001;
        x_t[63] = 26'b00000000011001110111101111;
        
        h_t_prev[0] = 26'b00000000001000100101100100;
        h_t_prev[1] = 26'b00000000001110100010010101;
        h_t_prev[2] = 26'b00000000001011010101001111;
        h_t_prev[3] = 26'b00000000001001100000111100;
        h_t_prev[4] = 26'b00000000000101100111111001;
        h_t_prev[5] = 26'b11111111111101011010010001;
        h_t_prev[6] = 26'b11111111110111101000010111;
        h_t_prev[7] = 26'b00000000011001001010100100;
        h_t_prev[8] = 26'b00000000010110000001010100;
        h_t_prev[9] = 26'b00000000010011100010001000;
        h_t_prev[10] = 26'b00000000010001001010001111;
        h_t_prev[11] = 26'b00000000001011011010011010;
        h_t_prev[12] = 26'b00000000000011001000010101;
        h_t_prev[13] = 26'b11111111110001101001100001;
        h_t_prev[14] = 26'b00000000011110000001101001;
        h_t_prev[15] = 26'b00000000011010001110100110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 42 timeout!");
                $fdisplay(fd_cycles, "Test Vector  42: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  42: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 42");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 43
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001011000011011010;
        x_t[1] = 26'b00000000001101100111100110;
        x_t[2] = 26'b00000000001010101110011000;
        x_t[3] = 26'b00000000001010011010111100;
        x_t[4] = 26'b00000000000110111000101110;
        x_t[5] = 26'b00000000000000100001111101;
        x_t[6] = 26'b11111111111110001111100100;
        x_t[7] = 26'b00000000010011011100000111;
        x_t[8] = 26'b00000000010001100000100000;
        x_t[9] = 26'b00000000010000000101101001;
        x_t[10] = 26'b00000000001111010100110100;
        x_t[11] = 26'b00000000001100101011111100;
        x_t[12] = 26'b00000000000110011011000010;
        x_t[13] = 26'b11111111111011110111101100;
        x_t[14] = 26'b00000000010110000111011001;
        x_t[15] = 26'b00000000010100100000011101;
        x_t[16] = 26'b00000000010011010010111111;
        x_t[17] = 26'b00000000001110011011100001;
        x_t[18] = 26'b00000000010000010100101001;
        x_t[19] = 26'b00000000001110000011011110;
        x_t[20] = 26'b00000000001001000110101110;
        x_t[21] = 26'b11111111111010111110111000;
        x_t[22] = 26'b11111111110101111000111010;
        x_t[23] = 26'b11111111111000110111110001;
        x_t[24] = 26'b11111111111100101100010110;
        x_t[25] = 26'b11111111111101011111011010;
        x_t[26] = 26'b11111111111001101000001001;
        x_t[27] = 26'b11111111111011101011011100;
        x_t[28] = 26'b11111111111000100010111010;
        x_t[29] = 26'b00000000000110110011101000;
        x_t[30] = 26'b11111111111110101001010011;
        x_t[31] = 26'b00000000000111101110000101;
        x_t[32] = 26'b00000000000011100100010011;
        x_t[33] = 26'b00000000000000111101010110;
        x_t[34] = 26'b11111111111110001000000000;
        x_t[35] = 26'b11111111111010111100100010;
        x_t[36] = 26'b11111111111001101100110110;
        x_t[37] = 26'b11111111110000010000011110;
        x_t[38] = 26'b00000000001101110100110000;
        x_t[39] = 26'b11111111111011110000011001;
        x_t[40] = 26'b00000000010100100100001110;
        x_t[41] = 26'b00000000001101100110001001;
        x_t[42] = 26'b00000000010110100000001110;
        x_t[43] = 26'b11111111111010010010111111;
        x_t[44] = 26'b00000000001110111001111011;
        x_t[45] = 26'b00000000000110010000100100;
        x_t[46] = 26'b00000000010110001000111000;
        x_t[47] = 26'b00000000010110011111100000;
        x_t[48] = 26'b00000000010011001111000000;
        x_t[49] = 26'b00000000011010010111101001;
        x_t[50] = 26'b00000000010011110011001111;
        x_t[51] = 26'b00000000010001000011001000;
        x_t[52] = 26'b00000000010000011100111011;
        x_t[53] = 26'b00000000001010101011111110;
        x_t[54] = 26'b00000000001010110011010110;
        x_t[55] = 26'b00000000011001111111101011;
        x_t[56] = 26'b00000000011100010001010101;
        x_t[57] = 26'b00000000011011100100100110;
        x_t[58] = 26'b00000000010000010100001100;
        x_t[59] = 26'b00000000010000001111000101;
        x_t[60] = 26'b00000000100001000000110010;
        x_t[61] = 26'b00000000011100011010011010;
        x_t[62] = 26'b00000000011000101100101101;
        x_t[63] = 26'b00000000011010101100100011;
        
        h_t_prev[0] = 26'b00000000001011000011011010;
        h_t_prev[1] = 26'b00000000001101100111100110;
        h_t_prev[2] = 26'b00000000001010101110011000;
        h_t_prev[3] = 26'b00000000001010011010111100;
        h_t_prev[4] = 26'b00000000000110111000101110;
        h_t_prev[5] = 26'b00000000000000100001111101;
        h_t_prev[6] = 26'b11111111111110001111100100;
        h_t_prev[7] = 26'b00000000010011011100000111;
        h_t_prev[8] = 26'b00000000010001100000100000;
        h_t_prev[9] = 26'b00000000010000000101101001;
        h_t_prev[10] = 26'b00000000001111010100110100;
        h_t_prev[11] = 26'b00000000001100101011111100;
        h_t_prev[12] = 26'b00000000000110011011000010;
        h_t_prev[13] = 26'b11111111111011110111101100;
        h_t_prev[14] = 26'b00000000010110000111011001;
        h_t_prev[15] = 26'b00000000010100100000011101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 43 timeout!");
                $fdisplay(fd_cycles, "Test Vector  43: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  43: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 43");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 44
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001010001000001110;
        x_t[1] = 26'b00000000001010010000001111;
        x_t[2] = 26'b00000000000111000101010011;
        x_t[3] = 26'b00000000000111101100111011;
        x_t[4] = 26'b00000000000100101011010001;
        x_t[5] = 26'b11111111111111110101100101;
        x_t[6] = 26'b00000000000100000100111110;
        x_t[7] = 26'b00000000001110111111000110;
        x_t[8] = 26'b00000000001100111111101100;
        x_t[9] = 26'b00000000001011011000111110;
        x_t[10] = 26'b00000000001100100100101100;
        x_t[11] = 26'b00000000001101000000010101;
        x_t[12] = 26'b00000000001000111110111011;
        x_t[13] = 26'b00000000000110100001000111;
        x_t[14] = 26'b00000000001111100001100001;
        x_t[15] = 26'b00000000001111101111010101;
        x_t[16] = 26'b00000000001110111101011010;
        x_t[17] = 26'b00000000001100100101000101;
        x_t[18] = 26'b00000000010000010100101001;
        x_t[19] = 26'b00000000010000000111010001;
        x_t[20] = 26'b00000000010000111011010010;
        x_t[21] = 26'b11111111111100111000011100;
        x_t[22] = 26'b11111111110111110111110101;
        x_t[23] = 26'b11111111111001110001110001;
        x_t[24] = 26'b11111111111111010110110110;
        x_t[25] = 26'b00000000000000000001000001;
        x_t[26] = 26'b11111111111100100010000000;
        x_t[27] = 26'b11111111111101001001110010;
        x_t[28] = 26'b11111111111001001000101100;
        x_t[29] = 26'b00000000001001111011010010;
        x_t[30] = 26'b00000000000001100100101000;
        x_t[31] = 26'b00000000001010001101110000;
        x_t[32] = 26'b00000000000111010000100010;
        x_t[33] = 26'b00000000000100101101111000;
        x_t[34] = 26'b00000000000001011001100101;
        x_t[35] = 26'b11111111111111100100100110;
        x_t[36] = 26'b11111111111110000011001010;
        x_t[37] = 26'b11111111110100100101101100;
        x_t[38] = 26'b00000000001110110001010001;
        x_t[39] = 26'b00000000000100111100010101;
        x_t[40] = 26'b00000000010010001100000011;
        x_t[41] = 26'b00000000010101011010110111;
        x_t[42] = 26'b00000000010110100000001110;
        x_t[43] = 26'b00000000000011001101100000;
        x_t[44] = 26'b00000000001000111110000101;
        x_t[45] = 26'b00000000001101100000110110;
        x_t[46] = 26'b00000000010011100011000110;
        x_t[47] = 26'b00000000010100111100000010;
        x_t[48] = 26'b00000000010010010101110100;
        x_t[49] = 26'b00000000011001100000000011;
        x_t[50] = 26'b00000000010100011001010000;
        x_t[51] = 26'b00000000010010110111000011;
        x_t[52] = 26'b00000000010100010010011110;
        x_t[53] = 26'b00000000010000100110100011;
        x_t[54] = 26'b00000000010001100010110101;
        x_t[55] = 26'b00000000010111010011000010;
        x_t[56] = 26'b00000000011001010100010010;
        x_t[57] = 26'b00000000011001111110010010;
        x_t[58] = 26'b00000000010010011111110001;
        x_t[59] = 26'b00000000010011001100100011;
        x_t[60] = 26'b00000000011101011010110000;
        x_t[61] = 26'b00000000011010010101111110;
        x_t[62] = 26'b00000000011001011001000110;
        x_t[63] = 26'b00000000010111111100100001;
        
        h_t_prev[0] = 26'b00000000001010001000001110;
        h_t_prev[1] = 26'b00000000001010010000001111;
        h_t_prev[2] = 26'b00000000000111000101010011;
        h_t_prev[3] = 26'b00000000000111101100111011;
        h_t_prev[4] = 26'b00000000000100101011010001;
        h_t_prev[5] = 26'b11111111111111110101100101;
        h_t_prev[6] = 26'b00000000000100000100111110;
        h_t_prev[7] = 26'b00000000001110111111000110;
        h_t_prev[8] = 26'b00000000001100111111101100;
        h_t_prev[9] = 26'b00000000001011011000111110;
        h_t_prev[10] = 26'b00000000001100100100101100;
        h_t_prev[11] = 26'b00000000001101000000010101;
        h_t_prev[12] = 26'b00000000001000111110111011;
        h_t_prev[13] = 26'b00000000000110100001000111;
        h_t_prev[14] = 26'b00000000001111100001100001;
        h_t_prev[15] = 26'b00000000001111101111010101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 44 timeout!");
                $fdisplay(fd_cycles, "Test Vector  44: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  44: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 44");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 45
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001110001000101110;
        x_t[1] = 26'b00000000001111110000101000;
        x_t[2] = 26'b00000000001110000100000010;
        x_t[3] = 26'b00000000001100110101101000;
        x_t[4] = 26'b00000000001001101110100110;
        x_t[5] = 26'b00000000000110000100111110;
        x_t[6] = 26'b00000000001001001000100110;
        x_t[7] = 26'b00000000010100011001001100;
        x_t[8] = 26'b00000000010010110011000001;
        x_t[9] = 26'b00000000010000011001101100;
        x_t[10] = 26'b00000000010000100011000110;
        x_t[11] = 26'b00000000001111100011011001;
        x_t[12] = 26'b00000000001110000110101101;
        x_t[13] = 26'b00000000001000001110001001;
        x_t[14] = 26'b00000000010011110011101111;
        x_t[15] = 26'b00000000010001111101101110;
        x_t[16] = 26'b00000000010000100000100011;
        x_t[17] = 26'b00000000001110011011100001;
        x_t[18] = 26'b00000000010000111110110100;
        x_t[19] = 26'b00000000010000110011001101;
        x_t[20] = 26'b00000000010010000110010111;
        x_t[21] = 26'b11111111111101100100101001;
        x_t[22] = 26'b11111111110111011110011100;
        x_t[23] = 26'b11111111111000101100001010;
        x_t[24] = 26'b11111111111110111110100000;
        x_t[25] = 26'b00000000000000011001111000;
        x_t[26] = 26'b11111111111110000111011000;
        x_t[27] = 26'b11111111111110101000000111;
        x_t[28] = 26'b11111111111000101111100000;
        x_t[29] = 26'b00000000000111100101100010;
        x_t[30] = 26'b00000000000010110010101011;
        x_t[31] = 26'b00000000001101010000111011;
        x_t[32] = 26'b00000000001001001111101111;
        x_t[33] = 26'b00000000000101100101011000;
        x_t[34] = 26'b00000000000010111000110110;
        x_t[35] = 26'b00000000000000110011100011;
        x_t[36] = 26'b00000000000001001001111101;
        x_t[37] = 26'b11111111111001011011100010;
        x_t[38] = 26'b00000000010000111110011101;
        x_t[39] = 26'b00000000000011100100001001;
        x_t[40] = 26'b00000000010101001111101101;
        x_t[41] = 26'b00000000001010100011011010;
        x_t[42] = 26'b00000000001101111110110000;
        x_t[43] = 26'b00000000001010110000001111;
        x_t[44] = 26'b00000000001000100111101111;
        x_t[45] = 26'b00000000001101111111110011;
        x_t[46] = 26'b00000000010001100110110000;
        x_t[47] = 26'b00000000010001100001001110;
        x_t[48] = 26'b00000000001110110001000111;
        x_t[49] = 26'b00000000010100010010011100;
        x_t[50] = 26'b00000000001111111100001011;
        x_t[51] = 26'b00000000001110000001111101;
        x_t[52] = 26'b00000000001110110110100111;
        x_t[53] = 26'b00000000001011101110110001;
        x_t[54] = 26'b00000000001100101011001101;
        x_t[55] = 26'b00000000010000100011011101;
        x_t[56] = 26'b00000000010010100110100111;
        x_t[57] = 26'b00000000010001011100100111;
        x_t[58] = 26'b00000000001011111101000010;
        x_t[59] = 26'b00000000001010010100001001;
        x_t[60] = 26'b00000000010101000010000010;
        x_t[61] = 26'b00000000001111011110101110;
        x_t[62] = 26'b00000000010010001110011100;
        x_t[63] = 26'b00000000001011010010110011;
        
        h_t_prev[0] = 26'b00000000001110001000101110;
        h_t_prev[1] = 26'b00000000001111110000101000;
        h_t_prev[2] = 26'b00000000001110000100000010;
        h_t_prev[3] = 26'b00000000001100110101101000;
        h_t_prev[4] = 26'b00000000001001101110100110;
        h_t_prev[5] = 26'b00000000000110000100111110;
        h_t_prev[6] = 26'b00000000001001001000100110;
        h_t_prev[7] = 26'b00000000010100011001001100;
        h_t_prev[8] = 26'b00000000010010110011000001;
        h_t_prev[9] = 26'b00000000010000011001101100;
        h_t_prev[10] = 26'b00000000010000100011000110;
        h_t_prev[11] = 26'b00000000001111100011011001;
        h_t_prev[12] = 26'b00000000001110000110101101;
        h_t_prev[13] = 26'b00000000001000001110001001;
        h_t_prev[14] = 26'b00000000010011110011101111;
        h_t_prev[15] = 26'b00000000010001111101101110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 45 timeout!");
                $fdisplay(fd_cycles, "Test Vector  45: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  45: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 45");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 46
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001101001101100010;
        x_t[1] = 26'b00000000010000010111110010;
        x_t[2] = 26'b00000000001101001001110001;
        x_t[3] = 26'b00000000001011101000010010;
        x_t[4] = 26'b00000000000111110101010110;
        x_t[5] = 26'b00000000000101000010011010;
        x_t[6] = 26'b00000000000110110011001111;
        x_t[7] = 26'b00000000010110100111101101;
        x_t[8] = 26'b00000000010011011100010010;
        x_t[9] = 26'b00000000010001010101110100;
        x_t[10] = 26'b00000000010001011101110100;
        x_t[11] = 26'b00000000001101101001000110;
        x_t[12] = 26'b00000000001101000000011110;
        x_t[13] = 26'b00000000000110000101110111;
        x_t[14] = 26'b00000000010111110000110111;
        x_t[15] = 26'b00000000010011110111110001;
        x_t[16] = 26'b00000000010001011100000010;
        x_t[17] = 26'b00000000001111000011000000;
        x_t[18] = 26'b00000000010000111110110100;
        x_t[19] = 26'b00000000010000011101001111;
        x_t[20] = 26'b00000000010000100010010000;
        x_t[21] = 26'b11111111111101100100101001;
        x_t[22] = 26'b11111111111000010001001110;
        x_t[23] = 26'b11111111110111111101110000;
        x_t[24] = 26'b11111111111111001010101011;
        x_t[25] = 26'b00000000000000011001111000;
        x_t[26] = 26'b11111111111110011000010010;
        x_t[27] = 26'b11111111111111100111000000;
        x_t[28] = 26'b11111111111001010101010010;
        x_t[29] = 26'b00000000000110110011101000;
        x_t[30] = 26'b00000000000101101110000000;
        x_t[31] = 26'b00000000001101100010101011;
        x_t[32] = 26'b00000000001011001110111100;
        x_t[33] = 26'b00000000000110011100111001;
        x_t[34] = 26'b00000000000010111000110110;
        x_t[35] = 26'b00000000000001101110110001;
        x_t[36] = 26'b00000000000000001110010100;
        x_t[37] = 26'b11111111111010011100110001;
        x_t[38] = 26'b00000000010100011100010100;
        x_t[39] = 26'b00000000000010101001010110;
        x_t[40] = 26'b00000000010010100001110010;
        x_t[41] = 26'b00000000000110001101001111;
        x_t[42] = 26'b00000000001111011101100111;
        x_t[43] = 26'b00000000010001100111000110;
        x_t[44] = 26'b00000000001011000100001001;
        x_t[45] = 26'b00000000010101010000000101;
        x_t[46] = 26'b00000000010100110101111111;
        x_t[47] = 26'b00000000010101001111111100;
        x_t[48] = 26'b00000000010010000010110001;
        x_t[49] = 26'b00000000010111110000110110;
        x_t[50] = 26'b00000000010100101100010000;
        x_t[51] = 26'b00000000010011110001000000;
        x_t[52] = 26'b00000000010100100110111100;
        x_t[53] = 26'b00000000010001010011000101;
        x_t[54] = 26'b00000000010011110010101011;
        x_t[55] = 26'b00000000010001101000100000;
        x_t[56] = 26'b00000000010100001101101111;
        x_t[57] = 26'b00000000010100111010010010;
        x_t[58] = 26'b00000000010001101011011011;
        x_t[59] = 26'b00000000010000001111000101;
        x_t[60] = 26'b00000000010000000000000000;
        x_t[61] = 26'b00000000001001010001011011;
        x_t[62] = 26'b00000000001110000100001001;
        x_t[63] = 26'b00000000000110100111100011;
        
        h_t_prev[0] = 26'b00000000001101001101100010;
        h_t_prev[1] = 26'b00000000010000010111110010;
        h_t_prev[2] = 26'b00000000001101001001110001;
        h_t_prev[3] = 26'b00000000001011101000010010;
        h_t_prev[4] = 26'b00000000000111110101010110;
        h_t_prev[5] = 26'b00000000000101000010011010;
        h_t_prev[6] = 26'b00000000000110110011001111;
        h_t_prev[7] = 26'b00000000010110100111101101;
        h_t_prev[8] = 26'b00000000010011011100010010;
        h_t_prev[9] = 26'b00000000010001010101110100;
        h_t_prev[10] = 26'b00000000010001011101110100;
        h_t_prev[11] = 26'b00000000001101101001000110;
        h_t_prev[12] = 26'b00000000001101000000011110;
        h_t_prev[13] = 26'b00000000000110000101110111;
        h_t_prev[14] = 26'b00000000010111110000110111;
        h_t_prev[15] = 26'b00000000010011110111110001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 46 timeout!");
                $fdisplay(fd_cycles, "Test Vector  46: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  46: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 46");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 47
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000010010110000101100;
        x_t[1] = 26'b00000000010101111000001011;
        x_t[2] = 26'b00000000010001101101000111;
        x_t[3] = 26'b00000000010001111110010110;
        x_t[4] = 26'b00000000001101001100111000;
        x_t[5] = 26'b00000000000111000111100010;
        x_t[6] = 26'b00000000000110011010010110;
        x_t[7] = 26'b00000000011010000111101001;
        x_t[8] = 26'b00000000010110101010100100;
        x_t[9] = 26'b00000000011000100010110110;
        x_t[10] = 26'b00000000011000001100010110;
        x_t[11] = 26'b00000000010101010010010011;
        x_t[12] = 26'b00000000010001000010000000;
        x_t[13] = 26'b00000000001000101001011001;
        x_t[14] = 26'b00000000010101011101001101;
        x_t[15] = 26'b00000000010110011010100000;
        x_t[16] = 26'b00000000010110101101000110;
        x_t[17] = 26'b00000000010101001101110011;
        x_t[18] = 26'b00000000010111111001100101;
        x_t[19] = 26'b00000000010110010010101100;
        x_t[20] = 26'b00000000010011010001011100;
        x_t[21] = 26'b11111111111101011001100110;
        x_t[22] = 26'b11111111111001011101011000;
        x_t[23] = 26'b11111111111001100110001011;
        x_t[24] = 26'b11111111111111001010101011;
        x_t[25] = 26'b00000000000000011001111000;
        x_t[26] = 26'b00000000000000110000010110;
        x_t[27] = 26'b00000000000000000110011100;
        x_t[28] = 26'b11111111111010100000110111;
        x_t[29] = 26'b00000000001011101111110000;
        x_t[30] = 26'b00000000000001100100101000;
        x_t[31] = 26'b00000000001100111111001100;
        x_t[32] = 26'b00000000001011110011010010;
        x_t[33] = 26'b00000000001000001011111010;
        x_t[34] = 26'b00000000000100000101000011;
        x_t[35] = 26'b00000000000000110011100011;
        x_t[36] = 26'b11111111111110010111000010;
        x_t[37] = 26'b11111111110111001000110001;
        x_t[38] = 26'b00000000001101100000100101;
        x_t[39] = 26'b00000000000001101110100011;
        x_t[40] = 26'b00000000000100100110100000;
        x_t[41] = 26'b00000000001010000111100110;
        x_t[42] = 26'b00000000010111001111101010;
        x_t[43] = 26'b00000000010000001111010101;
        x_t[44] = 26'b00000000001000111110000101;
        x_t[45] = 26'b00000000010010110101010100;
        x_t[46] = 26'b00000000010000010011111000;
        x_t[47] = 26'b00000000010001001101010101;
        x_t[48] = 26'b00000000001111101010010010;
        x_t[49] = 26'b00000000010100100100111110;
        x_t[50] = 26'b00000000010011110011001111;
        x_t[51] = 26'b00000000010100101010111101;
        x_t[52] = 26'b00000000010100010010011110;
        x_t[53] = 26'b00000000010000010000010010;
        x_t[54] = 26'b00000000010000110010111001;
        x_t[55] = 26'b00000000001101100101100011;
        x_t[56] = 26'b00000000010001110011000011;
        x_t[57] = 26'b00000000010011110110000101;
        x_t[58] = 26'b00000000010010011111110001;
        x_t[59] = 26'b00000000010000101110101010;
        x_t[60] = 26'b00000000001101110110000000;
        x_t[61] = 26'b00000000001001010001011011;
        x_t[62] = 26'b00000000001111001110000111;
        x_t[63] = 26'b00000000001001101001001100;
        
        h_t_prev[0] = 26'b00000000010010110000101100;
        h_t_prev[1] = 26'b00000000010101111000001011;
        h_t_prev[2] = 26'b00000000010001101101000111;
        h_t_prev[3] = 26'b00000000010001111110010110;
        h_t_prev[4] = 26'b00000000001101001100111000;
        h_t_prev[5] = 26'b00000000000111000111100010;
        h_t_prev[6] = 26'b00000000000110011010010110;
        h_t_prev[7] = 26'b00000000011010000111101001;
        h_t_prev[8] = 26'b00000000010110101010100100;
        h_t_prev[9] = 26'b00000000011000100010110110;
        h_t_prev[10] = 26'b00000000011000001100010110;
        h_t_prev[11] = 26'b00000000010101010010010011;
        h_t_prev[12] = 26'b00000000010001000010000000;
        h_t_prev[13] = 26'b00000000001000101001011001;
        h_t_prev[14] = 26'b00000000010101011101001101;
        h_t_prev[15] = 26'b00000000010110011010100000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 47 timeout!");
                $fdisplay(fd_cycles, "Test Vector  47: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  47: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 47");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 48
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001010101111101011;
        x_t[1] = 26'b00000000001101111011001011;
        x_t[2] = 26'b00000000001100100010111011;
        x_t[3] = 26'b00000000001111110110111111;
        x_t[4] = 26'b00000000001100010000010000;
        x_t[5] = 26'b00000000000110000100111110;
        x_t[6] = 26'b00000000000111100101000001;
        x_t[7] = 26'b00000000001011011111001001;
        x_t[8] = 26'b00000000001111111001010111;
        x_t[9] = 26'b00000000010001111101111010;
        x_t[10] = 26'b00000000010010111111101010;
        x_t[11] = 26'b00000000010001001001010100;
        x_t[12] = 26'b00000000010000010011001011;
        x_t[13] = 26'b00000000001000001110001001;
        x_t[14] = 26'b00000000001110100010001111;
        x_t[15] = 26'b00000000010001000000101100;
        x_t[16] = 26'b00000000010010000011101100;
        x_t[17] = 26'b00000000010000100101101101;
        x_t[18] = 26'b00000000010101100101111111;
        x_t[19] = 26'b00000000010100001110111000;
        x_t[20] = 26'b00000000010001010100010011;
        x_t[21] = 26'b11111111111100111000011100;
        x_t[22] = 26'b11111111111001000011111111;
        x_t[23] = 26'b11111111111001011010100100;
        x_t[24] = 26'b11111111111110001101110010;
        x_t[25] = 26'b11111111111111001111010010;
        x_t[26] = 26'b11111111111111101100110001;
        x_t[27] = 26'b11111111111111110110101110;
        x_t[28] = 26'b11111111111010000111101010;
        x_t[29] = 26'b00000000001001101010101001;
        x_t[30] = 26'b11111111111111011000001000;
        x_t[31] = 26'b00000000001100101101011100;
        x_t[32] = 26'b00000000001000000111000011;
        x_t[33] = 26'b00000000000101100101011000;
        x_t[34] = 26'b00000000000011001011111001;
        x_t[35] = 26'b11111111111111010000110111;
        x_t[36] = 26'b11111111111111100110100011;
        x_t[37] = 26'b11111111111001111100001010;
        x_t[38] = 26'b00000000001011100111100100;
        x_t[39] = 26'b00000000000100000001100010;
        x_t[40] = 26'b00000000001110000111001100;
        x_t[41] = 26'b00000000001111110001001111;
        x_t[42] = 26'b00000000011000010110110100;
        x_t[43] = 26'b11111111111010010010111111;
        x_t[44] = 26'b00000000001101001010001101;
        x_t[45] = 26'b00000000010011010100010001;
        x_t[46] = 26'b00000000001101011001010111;
        x_t[47] = 26'b00000000010001001101010101;
        x_t[48] = 26'b00000000001111010111001111;
        x_t[49] = 26'b00000000010100110111100000;
        x_t[50] = 26'b00000000010100101100010000;
        x_t[51] = 26'b00000000010111101100001001;
        x_t[52] = 26'b00000000010110100001101110;
        x_t[53] = 26'b00000000010011011000101101;
        x_t[54] = 26'b00000000010011110010101011;
        x_t[55] = 26'b00000000001110101010100111;
        x_t[56] = 26'b00000000010011101011010111;
        x_t[57] = 26'b00000000010111110101110111;
        x_t[58] = 26'b00000000010111111100101110;
        x_t[59] = 26'b00000000010110011001110011;
        x_t[60] = 26'b00000000001111000010101011;
        x_t[61] = 26'b00000000001110011100100000;
        x_t[62] = 26'b00000000010101011101100101;
        x_t[63] = 26'b00000000010001010110000100;
        
        h_t_prev[0] = 26'b00000000001010101111101011;
        h_t_prev[1] = 26'b00000000001101111011001011;
        h_t_prev[2] = 26'b00000000001100100010111011;
        h_t_prev[3] = 26'b00000000001111110110111111;
        h_t_prev[4] = 26'b00000000001100010000010000;
        h_t_prev[5] = 26'b00000000000110000100111110;
        h_t_prev[6] = 26'b00000000000111100101000001;
        h_t_prev[7] = 26'b00000000001011011111001001;
        h_t_prev[8] = 26'b00000000001111111001010111;
        h_t_prev[9] = 26'b00000000010001111101111010;
        h_t_prev[10] = 26'b00000000010010111111101010;
        h_t_prev[11] = 26'b00000000010001001001010100;
        h_t_prev[12] = 26'b00000000010000010011001011;
        h_t_prev[13] = 26'b00000000001000001110001001;
        h_t_prev[14] = 26'b00000000001110100010001111;
        h_t_prev[15] = 26'b00000000010001000000101100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 48 timeout!");
                $fdisplay(fd_cycles, "Test Vector  48: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  48: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 48");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 49
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111110011100111110111;
        x_t[1] = 26'b11111111101011111110000110;
        x_t[2] = 26'b11111111100011010001011000;
        x_t[3] = 26'b11111111011011111001001011;
        x_t[4] = 26'b11111111011110001001111001;
        x_t[5] = 26'b11111111011100001000001100;
        x_t[6] = 26'b11111111100011000000111110;
        x_t[7] = 26'b11111111110111011100100011;
        x_t[8] = 26'b11111111100011000101111010;
        x_t[9] = 26'b11111111100000110010111011;
        x_t[10] = 26'b11111111011110011001101010;
        x_t[11] = 26'b11111111011010101011101111;
        x_t[12] = 26'b11111111100000000000101101;
        x_t[13] = 26'b11111111011011100000001001;
        x_t[14] = 26'b11111111101000111101100001;
        x_t[15] = 26'b11111111100110000110100101;
        x_t[16] = 26'b11111111100010000010011100;
        x_t[17] = 26'b11111111011111110110110011;
        x_t[18] = 26'b11111111100101011111110000;
        x_t[19] = 26'b11111111100111010001001100;
        x_t[20] = 26'b11111111100101100001001101;
        x_t[21] = 26'b11111111110101010010001100;
        x_t[22] = 26'b11111111101100111101101111;
        x_t[23] = 26'b11111111101100101110011101;
        x_t[24] = 26'b11111111111100100000001010;
        x_t[25] = 26'b11111111111011101111100001;
        x_t[26] = 26'b11111111100000110011110110;
        x_t[27] = 26'b11111111011111011011011100;
        x_t[28] = 26'b11111111101001110010010001;
        x_t[29] = 26'b11111111110110111100101101;
        x_t[30] = 26'b11111111110010011100110001;
        x_t[31] = 26'b11111111011110011010011010;
        x_t[32] = 26'b11111111100000101001001001;
        x_t[33] = 26'b11111111011100100010000001;
        x_t[34] = 26'b11111111011010111111110110;
        x_t[35] = 26'b11111111100000000111010111;
        x_t[36] = 26'b11111111011101000111111100;
        x_t[37] = 26'b11111111110100000101000101;
        x_t[38] = 26'b11111111101110111100001000;
        x_t[39] = 26'b11111111011010101011110110;
        x_t[40] = 26'b11111111100110101101011111;
        x_t[41] = 26'b11111111011011001011010000;
        x_t[42] = 26'b11111111101010110001101100;
        x_t[43] = 26'b11111111110001011000011110;
        x_t[44] = 26'b11111111101101000010100111;
        x_t[45] = 26'b11111111110000011111101110;
        x_t[46] = 26'b11111111101100010111101011;
        x_t[47] = 26'b11111111101010101010100110;
        x_t[48] = 26'b11111111101000111100101010;
        x_t[49] = 26'b11111111100111101100010010;
        x_t[50] = 26'b11111111100100010010011010;
        x_t[51] = 26'b11111111101101001000010000;
        x_t[52] = 26'b11111111110000001010001101;
        x_t[53] = 26'b11111111110101000111010000;
        x_t[54] = 26'b11111111101111110101011000;
        x_t[55] = 26'b11111111111001111001010101;
        x_t[56] = 26'b11111111110001000010010001;
        x_t[57] = 26'b11111111110010100010100011;
        x_t[58] = 26'b11111111111001001001001010;
        x_t[59] = 26'b11111111111001110010010001;
        x_t[60] = 26'b00000000000011010011010001;
        x_t[61] = 26'b11111111111011000010111110;
        x_t[62] = 26'b00000000000001110100000000;
        x_t[63] = 26'b00000000000100101100010101;
        
        h_t_prev[0] = 26'b11111111110011100111110111;
        h_t_prev[1] = 26'b11111111101011111110000110;
        h_t_prev[2] = 26'b11111111100011010001011000;
        h_t_prev[3] = 26'b11111111011011111001001011;
        h_t_prev[4] = 26'b11111111011110001001111001;
        h_t_prev[5] = 26'b11111111011100001000001100;
        h_t_prev[6] = 26'b11111111100011000000111110;
        h_t_prev[7] = 26'b11111111110111011100100011;
        h_t_prev[8] = 26'b11111111100011000101111010;
        h_t_prev[9] = 26'b11111111100000110010111011;
        h_t_prev[10] = 26'b11111111011110011001101010;
        h_t_prev[11] = 26'b11111111011010101011101111;
        h_t_prev[12] = 26'b11111111100000000000101101;
        h_t_prev[13] = 26'b11111111011011100000001001;
        h_t_prev[14] = 26'b11111111101000111101100001;
        h_t_prev[15] = 26'b11111111100110000110100101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 49 timeout!");
                $fdisplay(fd_cycles, "Test Vector  49: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  49: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 49");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 50
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111101011100110110111;
        x_t[1] = 26'b11111111100100111011110100;
        x_t[2] = 26'b11111111011010011110000111;
        x_t[3] = 26'b11111111010010001110011011;
        x_t[4] = 26'b11111111010001110101110010;
        x_t[5] = 26'b11111111001101111010011111;
        x_t[6] = 26'b11111111011001010010100111;
        x_t[7] = 26'b11111111101111110011111100;
        x_t[8] = 26'b11111111011100101001010101;
        x_t[9] = 26'b11111111011001111001111100;
        x_t[10] = 26'b11111111010111000011111111;
        x_t[11] = 26'b11111111010100010100000100;
        x_t[12] = 26'b11111111010100010011100000;
        x_t[13] = 26'b11111111010101100010100011;
        x_t[14] = 26'b11111111100100101011010011;
        x_t[15] = 26'b11111111100000011000011100;
        x_t[16] = 26'b11111111011100110001011000;
        x_t[17] = 26'b11111111011011001110101101;
        x_t[18] = 26'b11111111011110111010000100;
        x_t[19] = 26'b11111111011111010111111100;
        x_t[20] = 26'b11111111011110110111101111;
        x_t[21] = 26'b11111111110011000010100010;
        x_t[22] = 26'b11111111101011011000001100;
        x_t[23] = 26'b11111111101011101000110110;
        x_t[24] = 26'b11111111111011101111011100;
        x_t[25] = 26'b11111111111010111101110011;
        x_t[26] = 26'b11111111011100010100100110;
        x_t[27] = 26'b11111111011011011111111001;
        x_t[28] = 26'b11111111101000110011010011;
        x_t[29] = 26'b11111111110111001101010110;
        x_t[30] = 26'b11111111110001111101100011;
        x_t[31] = 26'b11111111011001011011000011;
        x_t[32] = 26'b11111111011100000110011001;
        x_t[33] = 26'b11111111010111000010011101;
        x_t[34] = 26'b11111111010101010101110110;
        x_t[35] = 26'b11111111011010100100000101;
        x_t[36] = 26'b11111111011000001001111000;
        x_t[37] = 26'b11111111110010010010111011;
        x_t[38] = 26'b11111111101111111000101000;
        x_t[39] = 26'b11111111011000011000110111;
        x_t[40] = 26'b11111111101000101111111011;
        x_t[41] = 26'b11111111010011110010010101;
        x_t[42] = 26'b11111111110111000000010101;
        x_t[43] = 26'b11111111100001100111000110;
        x_t[44] = 26'b11111111110001111011011011;
        x_t[45] = 26'b11111111101110100011111011;
        x_t[46] = 26'b11111111110000111001110011;
        x_t[47] = 26'b11111111101100100001111101;
        x_t[48] = 26'b11111111101010011011111101;
        x_t[49] = 26'b11111111101010100101100111;
        x_t[50] = 26'b11111111100111100011011101;
        x_t[51] = 26'b11111111101111100010110011;
        x_t[52] = 26'b11111111110000110011001000;
        x_t[53] = 26'b11111111110101000111010000;
        x_t[54] = 26'b11111111110001101101001111;
        x_t[55] = 26'b11111111111011100000111010;
        x_t[56] = 26'b11111111110010111010100101;
        x_t[57] = 26'b11111111110111110111100101;
        x_t[58] = 26'b11111111111001101100000011;
        x_t[59] = 26'b11111111111001000010111010;
        x_t[60] = 26'b11111111111110000001111010;
        x_t[61] = 26'b11111111110111101011110010;
        x_t[62] = 26'b11111111111100010000111011;
        x_t[63] = 26'b11111111111001101100001110;
        
        h_t_prev[0] = 26'b11111111101011100110110111;
        h_t_prev[1] = 26'b11111111100100111011110100;
        h_t_prev[2] = 26'b11111111011010011110000111;
        h_t_prev[3] = 26'b11111111010010001110011011;
        h_t_prev[4] = 26'b11111111010001110101110010;
        h_t_prev[5] = 26'b11111111001101111010011111;
        h_t_prev[6] = 26'b11111111011001010010100111;
        h_t_prev[7] = 26'b11111111101111110011111100;
        h_t_prev[8] = 26'b11111111011100101001010101;
        h_t_prev[9] = 26'b11111111011001111001111100;
        h_t_prev[10] = 26'b11111111010111000011111111;
        h_t_prev[11] = 26'b11111111010100010100000100;
        h_t_prev[12] = 26'b11111111010100010011100000;
        h_t_prev[13] = 26'b11111111010101100010100011;
        h_t_prev[14] = 26'b11111111100100101011010011;
        h_t_prev[15] = 26'b11111111100000011000011100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 50 timeout!");
                $fdisplay(fd_cycles, "Test Vector  50: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  50: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 50");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 51
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111101100100010000011;
        x_t[1] = 26'b11111111100100010100101010;
        x_t[2] = 26'b11111111011100100110000101;
        x_t[3] = 26'b11111111010100111100011100;
        x_t[4] = 26'b11111111010100101011101001;
        x_t[5] = 26'b11111111010011000111010011;
        x_t[6] = 26'b11111111011101001011100100;
        x_t[7] = 26'b11111111110010010110110100;
        x_t[8] = 26'b11111111100001110011011001;
        x_t[9] = 26'b11111111011111100010110000;
        x_t[10] = 26'b11111111011101110010100001;
        x_t[11] = 26'b11111111011011010100100000;
        x_t[12] = 26'b11111111010111111101101000;
        x_t[13] = 26'b11111111011000111100100110;
        x_t[14] = 26'b11111111101011111011010111;
        x_t[15] = 26'b11111111100111101100010010;
        x_t[16] = 26'b11111111100100110100111001;
        x_t[17] = 26'b11111111100010111100001101;
        x_t[18] = 26'b11111111100110001001111010;
        x_t[19] = 26'b11111111100101100011010111;
        x_t[20] = 26'b11111111100010011000111111;
        x_t[21] = 26'b11111111110100111100000110;
        x_t[22] = 26'b11111111101101010111000111;
        x_t[23] = 26'b11111111101101101000011110;
        x_t[24] = 26'b11111111111110001101110010;
        x_t[25] = 26'b11111111111101101011110101;
        x_t[26] = 26'b11111111100000110011110110;
        x_t[27] = 26'b11111111011111011011011100;
        x_t[28] = 26'b11111111101010100100101010;
        x_t[29] = 26'b11111111111010110110010001;
        x_t[30] = 26'b11111111110110010110100010;
        x_t[31] = 26'b11111111100000101000010110;
        x_t[32] = 26'b11111111100010000100000000;
        x_t[33] = 26'b11111111011100100010000001;
        x_t[34] = 26'b11111111011011111001000000;
        x_t[35] = 26'b11111111100001010110010100;
        x_t[36] = 26'b11111111011110010111011101;
        x_t[37] = 26'b11111111111001011011100010;
        x_t[38] = 26'b11111111111001010101101110;
        x_t[39] = 26'b11111111100011011010011000;
        x_t[40] = 26'b11111111111011011011100011;
        x_t[41] = 26'b11111111100000011001000100;
        x_t[42] = 26'b11111111111010101101100000;
        x_t[43] = 26'b11111111100110011010010011;
        x_t[44] = 26'b11111111111011101101000010;
        x_t[45] = 26'b11111111111010001010110001;
        x_t[46] = 26'b11111111111000111111110111;
        x_t[47] = 26'b11111111110101001110111101;
        x_t[48] = 26'b11111111110011010111101101;
        x_t[49] = 26'b11111111110101000000110100;
        x_t[50] = 26'b11111111110011011011101011;
        x_t[51] = 26'b11111111111000111001101010;
        x_t[52] = 26'b11111111111001000111001010;
        x_t[53] = 26'b11111111111011101110011000;
        x_t[54] = 26'b11111111111001001100101011;
        x_t[55] = 26'b11111111111100110111001110;
        x_t[56] = 26'b11111111110110111100011000;
        x_t[57] = 26'b00000000000000001000001101;
        x_t[58] = 26'b11111111111110010100101010;
        x_t[59] = 26'b11111111111010010001110110;
        x_t[60] = 26'b11111111111100000111001110;
        x_t[61] = 26'b11111111111000011101011100;
        x_t[62] = 26'b11111111111100101110100001;
        x_t[63] = 26'b11111111110111011111011010;
        
        h_t_prev[0] = 26'b11111111101100100010000011;
        h_t_prev[1] = 26'b11111111100100010100101010;
        h_t_prev[2] = 26'b11111111011100100110000101;
        h_t_prev[3] = 26'b11111111010100111100011100;
        h_t_prev[4] = 26'b11111111010100101011101001;
        h_t_prev[5] = 26'b11111111010011000111010011;
        h_t_prev[6] = 26'b11111111011101001011100100;
        h_t_prev[7] = 26'b11111111110010010110110100;
        h_t_prev[8] = 26'b11111111100001110011011001;
        h_t_prev[9] = 26'b11111111011111100010110000;
        h_t_prev[10] = 26'b11111111011101110010100001;
        h_t_prev[11] = 26'b11111111011011010100100000;
        h_t_prev[12] = 26'b11111111010111111101101000;
        h_t_prev[13] = 26'b11111111011000111100100110;
        h_t_prev[14] = 26'b11111111101011111011010111;
        h_t_prev[15] = 26'b11111111100111101100010010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 51 timeout!");
                $fdisplay(fd_cycles, "Test Vector  51: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  51: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 51");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 52
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111110110101101001011;
        x_t[1] = 26'b11111111110000100011110000;
        x_t[2] = 26'b11111111100111110100101111;
        x_t[3] = 26'b11111111011111110100100011;
        x_t[4] = 26'b11111111100000000011001001;
        x_t[5] = 26'b11111111011111001111111001;
        x_t[6] = 26'b11111111101011001011110000;
        x_t[7] = 26'b00000000000011001101110100;
        x_t[8] = 26'b11111111101111010101110100;
        x_t[9] = 26'b11111111101110111000111011;
        x_t[10] = 26'b11111111101101000101000000;
        x_t[11] = 26'b11111111100110001001100010;
        x_t[12] = 26'b11111111100101011111111001;
        x_t[13] = 26'b11111111100100011100100011;
        x_t[14] = 26'b11111111111011000101101100;
        x_t[15] = 26'b11111111110101101011010100;
        x_t[16] = 26'b11111111110010011101010011;
        x_t[17] = 26'b11111111110001011011111110;
        x_t[18] = 26'b11111111110010010110000001;
        x_t[19] = 26'b11111111110000111000010001;
        x_t[20] = 26'b11111111101011011000101000;
        x_t[21] = 26'b11111111111000001110000100;
        x_t[22] = 26'b11111111110000111011100101;
        x_t[23] = 26'b11111111110000100010000110;
        x_t[24] = 26'b00000000000001101001000000;
        x_t[25] = 26'b00000000000001001011100111;
        x_t[26] = 26'b11111111100101000010001100;
        x_t[27] = 26'b11111111100011110110011011;
        x_t[28] = 26'b11111111101101101110001011;
        x_t[29] = 26'b11111111111111100001110000;
        x_t[30] = 26'b11111111111010011111111011;
        x_t[31] = 26'b11111111100101010101111111;
        x_t[32] = 26'b11111111101001011100011110;
        x_t[33] = 26'b11111111100100000011000101;
        x_t[34] = 26'b11111111100010101111001101;
        x_t[35] = 26'b11111111101000011100010001;
        x_t[36] = 26'b11111111100111000100000101;
        x_t[37] = 26'b11111111111110110001111111;
        x_t[38] = 26'b00000000000000111001110011;
        x_t[39] = 26'b11111111101010110000101110;
        x_t[40] = 26'b11111111111100000111000010;
        x_t[41] = 26'b11111111110000000010100001;
        x_t[42] = 26'b11111111111011011100111011;
        x_t[43] = 26'b11111111111111110010000100;
        x_t[44] = 26'b11111111111110110110001000;
        x_t[45] = 26'b11111111111100000110100101;
        x_t[46] = 26'b11111111110110101110110011;
        x_t[47] = 26'b11111111110111000110010100;
        x_t[48] = 26'b11111111110110010110010011;
        x_t[49] = 26'b11111111111000001100101100;
        x_t[50] = 26'b11111111111001101010110010;
        x_t[51] = 26'b11111111111100001110001010;
        x_t[52] = 26'b11111111111011010110011001;
        x_t[53] = 26'b11111111111100000100101001;
        x_t[54] = 26'b11111111110111101100110010;
        x_t[55] = 26'b11111111111010001010100110;
        x_t[56] = 26'b11111111110101010101010000;
        x_t[57] = 26'b00000000000000101010010100;
        x_t[58] = 26'b11111111111100101011111110;
        x_t[59] = 26'b11111111110101000110010010;
        x_t[60] = 26'b11111111111010101011001110;
        x_t[61] = 26'b11111111111000101101111111;
        x_t[62] = 26'b11111111111101101001101100;
        x_t[63] = 26'b11111111110110111100001100;
        
        h_t_prev[0] = 26'b11111111110110101101001011;
        h_t_prev[1] = 26'b11111111110000100011110000;
        h_t_prev[2] = 26'b11111111100111110100101111;
        h_t_prev[3] = 26'b11111111011111110100100011;
        h_t_prev[4] = 26'b11111111100000000011001001;
        h_t_prev[5] = 26'b11111111011111001111111001;
        h_t_prev[6] = 26'b11111111101011001011110000;
        h_t_prev[7] = 26'b00000000000011001101110100;
        h_t_prev[8] = 26'b11111111101111010101110100;
        h_t_prev[9] = 26'b11111111101110111000111011;
        h_t_prev[10] = 26'b11111111101101000101000000;
        h_t_prev[11] = 26'b11111111100110001001100010;
        h_t_prev[12] = 26'b11111111100101011111111001;
        h_t_prev[13] = 26'b11111111100100011100100011;
        h_t_prev[14] = 26'b11111111111011000101101100;
        h_t_prev[15] = 26'b11111111110101101011010100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 52 timeout!");
                $fdisplay(fd_cycles, "Test Vector  52: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  52: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 52");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 53
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111111110101110001011;
        x_t[1] = 26'b11111111111000001101001011;
        x_t[2] = 26'b11111111110000101000000000;
        x_t[3] = 26'b11111111101010111111111111;
        x_t[4] = 26'b11111111101010110010001101;
        x_t[5] = 26'b11111111101000111101001010;
        x_t[6] = 26'b11111111110100100001001101;
        x_t[7] = 26'b00000000000110011001011010;
        x_t[8] = 26'b11111111110011001101010111;
        x_t[9] = 26'b11111111110101110001111010;
        x_t[10] = 26'b11111111110101111100100010;
        x_t[11] = 26'b11111111101101011110010111;
        x_t[12] = 26'b11111111101110010001110011;
        x_t[13] = 26'b11111111101100100010011011;
        x_t[14] = 26'b11111111110111001000100100;
        x_t[15] = 26'b11111111110110010100000000;
        x_t[16] = 26'b11111111110110011111000011;
        x_t[17] = 26'b11111111110101110000010101;
        x_t[18] = 26'b11111111110110101000000111;
        x_t[19] = 26'b11111111110100101001111010;
        x_t[20] = 26'b11111111101111010010111001;
        x_t[21] = 26'b11111111111001111100100101;
        x_t[22] = 26'b11111111110011111001111110;
        x_t[23] = 26'b11111111110100010101101110;
        x_t[24] = 26'b00000000000010111110010001;
        x_t[25] = 26'b00000000000010101111000100;
        x_t[26] = 26'b11111111101001110010010101;
        x_t[27] = 26'b11111111101001100000000010;
        x_t[28] = 26'b11111111110010101001000011;
        x_t[29] = 26'b00000000000000110100111101;
        x_t[30] = 26'b11111111111110111000111010;
        x_t[31] = 26'b11111111101100010001100011;
        x_t[32] = 26'b11111111101101111111001110;
        x_t[33] = 26'b11111111101001110101001000;
        x_t[34] = 26'b11111111101000101100010000;
        x_t[35] = 26'b11111111101101111111100011;
        x_t[36] = 26'b11111111101101111001011011;
        x_t[37] = 26'b00000000000011010111100010;
        x_t[38] = 26'b00000000000000010001011101;
        x_t[39] = 26'b11111111110000010001011111;
        x_t[40] = 26'b11111111111001101110110111;
        x_t[41] = 26'b11111111101110101111000100;
        x_t[42] = 26'b00000000000111010011110111;
        x_t[43] = 26'b11111111111101101110011010;
        x_t[44] = 26'b00000000000010010101100011;
        x_t[45] = 26'b11111111110111010001000011;
        x_t[46] = 26'b11111111110110011010000101;
        x_t[47] = 26'b11111111110100111011000100;
        x_t[48] = 26'b11111111110100100011111100;
        x_t[49] = 26'b11111111110111000010100011;
        x_t[50] = 26'b11111111111001101010110010;
        x_t[51] = 26'b11111111111011000000111001;
        x_t[52] = 26'b11111111111001011011101000;
        x_t[53] = 26'b11111111111001010010011111;
        x_t[54] = 26'b11111111110000001101010110;
        x_t[55] = 26'b11111111110101110110011000;
        x_t[56] = 26'b11111111110001010011011101;
        x_t[57] = 26'b11111111111101001100101000;
        x_t[58] = 26'b11111111110110011010101100;
        x_t[59] = 26'b11111111101110111011100011;
        x_t[60] = 26'b11111111110110100110100010;
        x_t[61] = 26'b11111111110100010100100101;
        x_t[62] = 26'b11111111111000010101011010;
        x_t[63] = 26'b11111111110011010111010111;
        
        h_t_prev[0] = 26'b11111111111110101110001011;
        h_t_prev[1] = 26'b11111111111000001101001011;
        h_t_prev[2] = 26'b11111111110000101000000000;
        h_t_prev[3] = 26'b11111111101010111111111111;
        h_t_prev[4] = 26'b11111111101010110010001101;
        h_t_prev[5] = 26'b11111111101000111101001010;
        h_t_prev[6] = 26'b11111111110100100001001101;
        h_t_prev[7] = 26'b00000000000110011001011010;
        h_t_prev[8] = 26'b11111111110011001101010111;
        h_t_prev[9] = 26'b11111111110101110001111010;
        h_t_prev[10] = 26'b11111111110101111100100010;
        h_t_prev[11] = 26'b11111111101101011110010111;
        h_t_prev[12] = 26'b11111111101110010001110011;
        h_t_prev[13] = 26'b11111111101100100010011011;
        h_t_prev[14] = 26'b11111111110111001000100100;
        h_t_prev[15] = 26'b11111111110110010100000000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 53 timeout!");
                $fdisplay(fd_cycles, "Test Vector  53: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  53: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 53");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 54
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111111101011111010000;
        x_t[1] = 26'b11111111110111100110000010;
        x_t[2] = 26'b11111111110001001110110110;
        x_t[3] = 26'b11111111101100110100000000;
        x_t[4] = 26'b11111111101100010111010000;
        x_t[5] = 26'b11111111101001111111101110;
        x_t[6] = 26'b11111111110010111101101000;
        x_t[7] = 26'b00000000000011110110100010;
        x_t[8] = 26'b11111111110001111010110110;
        x_t[9] = 26'b11111111110011111001101001;
        x_t[10] = 26'b11111111110011001100011010;
        x_t[11] = 26'b11111111101010111011010011;
        x_t[12] = 26'b11111111101101100010111110;
        x_t[13] = 26'b11111111101110001111011101;
        x_t[14] = 26'b11111111110110011110011000;
        x_t[15] = 26'b11111111110100011001111101;
        x_t[16] = 26'b11111111110100010100010000;
        x_t[17] = 26'b11111111110010010111001100;
        x_t[18] = 26'b11111111110010101011000110;
        x_t[19] = 26'b11111111110000100010010011;
        x_t[20] = 26'b11111111101011110001101001;
        x_t[21] = 26'b11111111111010010010101011;
        x_t[22] = 26'b11111111110100100000000011;
        x_t[23] = 26'b11111111110101110010100010;
        x_t[24] = 26'b00000000000011001010011100;
        x_t[25] = 26'b00000000000010101111000100;
        x_t[26] = 26'b11111111101010000011001110;
        x_t[27] = 26'b11111111101011011101110011;
        x_t[28] = 26'b11111111110100001101110100;
        x_t[29] = 26'b00000000000001100110110111;
        x_t[30] = 26'b11111111111111011000001000;
        x_t[31] = 26'b11111111101101000110110001;
        x_t[32] = 26'b11111111101101101101000011;
        x_t[33] = 26'b11111111101000111101101000;
        x_t[34] = 26'b11111111101000101100010000;
        x_t[35] = 26'b11111111101110100111000010;
        x_t[36] = 26'b11111111101101111001011011;
        x_t[37] = 26'b00000000000110011011001110;
        x_t[38] = 26'b11111111111111010100111101;
        x_t[39] = 26'b11111111110001001100010001;
        x_t[40] = 26'b00000000000101100111101110;
        x_t[41] = 26'b11111111101100001000001001;
        x_t[42] = 26'b00000000000100101101110110;
        x_t[43] = 26'b11111111100101101110011010;
        x_t[44] = 26'b00000000001010000001000111;
        x_t[45] = 26'b11111111101100101000000111;
        x_t[46] = 26'b11111111111000101011001000;
        x_t[47] = 26'b11111111110101100010110110;
        x_t[48] = 26'b11111111110011101010110001;
        x_t[49] = 26'b11111111110011110110101100;
        x_t[50] = 26'b11111111110011011011101011;
        x_t[51] = 26'b11111111110010010000101010;
        x_t[52] = 26'b11111111110000011110101011;
        x_t[53] = 26'b11111111110000001111011111;
        x_t[54] = 26'b11111111101000010101111100;
        x_t[55] = 26'b11111111110010111000011111;
        x_t[56] = 26'b11111111101110010110011010;
        x_t[57] = 26'b11111111110110110011011000;
        x_t[58] = 26'b11111111101011110010001111;
        x_t[59] = 26'b11111111100111010010000110;
        x_t[60] = 26'b11111111110001000101110101;
        x_t[61] = 26'b11111111101100110100100001;
        x_t[62] = 26'b11111111101101011110000011;
        x_t[63] = 26'b11111111101111001111010100;
        
        h_t_prev[0] = 26'b11111111111101011111010000;
        h_t_prev[1] = 26'b11111111110111100110000010;
        h_t_prev[2] = 26'b11111111110001001110110110;
        h_t_prev[3] = 26'b11111111101100110100000000;
        h_t_prev[4] = 26'b11111111101100010111010000;
        h_t_prev[5] = 26'b11111111101001111111101110;
        h_t_prev[6] = 26'b11111111110010111101101000;
        h_t_prev[7] = 26'b00000000000011110110100010;
        h_t_prev[8] = 26'b11111111110001111010110110;
        h_t_prev[9] = 26'b11111111110011111001101001;
        h_t_prev[10] = 26'b11111111110011001100011010;
        h_t_prev[11] = 26'b11111111101010111011010011;
        h_t_prev[12] = 26'b11111111101101100010111110;
        h_t_prev[13] = 26'b11111111101110001111011101;
        h_t_prev[14] = 26'b11111111110110011110011000;
        h_t_prev[15] = 26'b11111111110100011001111101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 54 timeout!");
                $fdisplay(fd_cycles, "Test Vector  54: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  54: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 54");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 55
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111111100110111110010;
        x_t[1] = 26'b11111111110110000100001001;
        x_t[2] = 26'b11111111101101111001001100;
        x_t[3] = 26'b11111111101000010001111101;
        x_t[4] = 26'b11111111101000010000100011;
        x_t[5] = 26'b11111111100110100001110110;
        x_t[6] = 26'b11111111101110101011110011;
        x_t[7] = 26'b00000000000011100010001011;
        x_t[8] = 26'b11111111110010111000101111;
        x_t[9] = 26'b11111111110000110001001100;
        x_t[10] = 26'b11111111101101111111101110;
        x_t[11] = 26'b11111111100101001100011001;
        x_t[12] = 26'b11111111101001111000110110;
        x_t[13] = 26'b11111111100111110110100110;
        x_t[14] = 26'b11111111111100000100111110;
        x_t[15] = 26'b11111111110100000101100111;
        x_t[16] = 26'b11111111110001001101111111;
        x_t[17] = 26'b11111111101100110011111000;
        x_t[18] = 26'b11111111101101101110110110;
        x_t[19] = 26'b11111111101011101110110001;
        x_t[20] = 26'b11111111100111011110010110;
        x_t[21] = 26'b11111111111001111100100101;
        x_t[22] = 26'b11111111110011100000100110;
        x_t[23] = 26'b11111111110011010000000111;
        x_t[24] = 26'b00000000000010111110010001;
        x_t[25] = 26'b00000000000010101111000100;
        x_t[26] = 26'b11111111100111111100000011;
        x_t[27] = 26'b11111111101000100001001001;
        x_t[28] = 26'b11111111110001101010000101;
        x_t[29] = 26'b00000000000010001000001001;
        x_t[30] = 26'b11111111111101001011101000;
        x_t[31] = 26'b11111111101001001110011000;
        x_t[32] = 26'b11111111101011011011101011;
        x_t[33] = 26'b11111111100101110010000110;
        x_t[34] = 26'b11111111100101000111100111;
        x_t[35] = 26'b11111111101011100001101010;
        x_t[36] = 26'b11111111101000010011100110;
        x_t[37] = 26'b00000000000000100100001001;
        x_t[38] = 26'b00000000000100101011110101;
        x_t[39] = 26'b11111111100111000101100011;
        x_t[40] = 26'b00000000001011000011100010;
        x_t[41] = 26'b11111111010010111010101101;
        x_t[42] = 26'b00000000001000011011000000;
        x_t[43] = 26'b11111111111011101010110000;
        x_t[44] = 26'b00000000001001010100011011;
        x_t[45] = 26'b11111111110001111100100101;
        x_t[46] = 26'b11111111110111011000001111;
        x_t[47] = 26'b11111111110100100111001011;
        x_t[48] = 26'b11111111110001100101010111;
        x_t[49] = 26'b11111111101111110011001110;
        x_t[50] = 26'b11111111101110011000100101;
        x_t[51] = 26'b11111111101011111010111110;
        x_t[52] = 26'b11111111101100000000001100;
        x_t[53] = 26'b11111111101101110011100110;
        x_t[54] = 26'b11111111101011101101101100;
        x_t[55] = 26'b11111111110000111111101001;
        x_t[56] = 26'b11111111101101000000011110;
        x_t[57] = 26'b11111111110001101111011000;
        x_t[58] = 26'b11111111101000001111011010;
        x_t[59] = 26'b11111111100111010010000110;
        x_t[60] = 26'b11111111101100010011001000;
        x_t[61] = 26'b11111111100111011000111001;
        x_t[62] = 26'b11111111100100011101000011;
        x_t[63] = 26'b11111111101101000010100000;
        
        h_t_prev[0] = 26'b11111111111100110111110010;
        h_t_prev[1] = 26'b11111111110110000100001001;
        h_t_prev[2] = 26'b11111111101101111001001100;
        h_t_prev[3] = 26'b11111111101000010001111101;
        h_t_prev[4] = 26'b11111111101000010000100011;
        h_t_prev[5] = 26'b11111111100110100001110110;
        h_t_prev[6] = 26'b11111111101110101011110011;
        h_t_prev[7] = 26'b00000000000011100010001011;
        h_t_prev[8] = 26'b11111111110010111000101111;
        h_t_prev[9] = 26'b11111111110000110001001100;
        h_t_prev[10] = 26'b11111111101101111111101110;
        h_t_prev[11] = 26'b11111111100101001100011001;
        h_t_prev[12] = 26'b11111111101001111000110110;
        h_t_prev[13] = 26'b11111111100111110110100110;
        h_t_prev[14] = 26'b11111111111100000100111110;
        h_t_prev[15] = 26'b11111111110100000101100111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 55 timeout!");
                $fdisplay(fd_cycles, "Test Vector  55: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  55: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 55");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 56
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111111011101000110111;
        x_t[1] = 26'b11111111110011010011111100;
        x_t[2] = 26'b11111111101010110110111101;
        x_t[3] = 26'b11111111100110110001010010;
        x_t[4] = 26'b11111111100110010111010011;
        x_t[5] = 26'b11111111100100110010111010;
        x_t[6] = 26'b11111111101001101000001011;
        x_t[7] = 26'b00000000000000010110100110;
        x_t[8] = 26'b11111111101111111111000100;
        x_t[9] = 26'b11111111101101101000110000;
        x_t[10] = 26'b11111111101100001010010011;
        x_t[11] = 26'b11111111100100100011101000;
        x_t[12] = 26'b11111111101000000011110010;
        x_t[13] = 26'b11111111100000001011111110;
        x_t[14] = 26'b11111111111001000111001000;
        x_t[15] = 26'b11111111110001100010111000;
        x_t[16] = 26'b11111111101101110011111000;
        x_t[17] = 26'b11111111101010000010001110;
        x_t[18] = 26'b11111111101011110000010110;
        x_t[19] = 26'b11111111101010000000111011;
        x_t[20] = 26'b11111111100110101100010010;
        x_t[21] = 26'b11111111110111110111111101;
        x_t[22] = 26'b11111111110001101110010111;
        x_t[23] = 26'b11111111110001000100111001;
        x_t[24] = 26'b00000000000010000001010111;
        x_t[25] = 26'b00000000000001110000111010;
        x_t[26] = 26'b11111111100110111000011110;
        x_t[27] = 26'b11111111100110100011011000;
        x_t[28] = 26'b11111111110000101011000110;
        x_t[29] = 26'b00000000000010001000001001;
        x_t[30] = 26'b11111111111101011011010000;
        x_t[31] = 26'b11111111101000101010111001;
        x_t[32] = 26'b11111111101000100101111101;
        x_t[33] = 26'b11111111100100010101100101;
        x_t[34] = 26'b11111111100011101000010111;
        x_t[35] = 26'b11111111101001101011001110;
        x_t[36] = 26'b11111111100111000100000101;
        x_t[37] = 26'b11111111111100111111110110;
        x_t[38] = 26'b00000000000000100101101000;
        x_t[39] = 26'b11111111100101101101010111;
        x_t[40] = 26'b00000000000100010000110000;
        x_t[41] = 26'b11111111100010001000010101;
        x_t[42] = 26'b00000000000110001100101101;
        x_t[43] = 26'b11111111111010010010111111;
        x_t[44] = 26'b00000000000010101011111001;
        x_t[45] = 26'b11111111111001001100110111;
        x_t[46] = 26'b11111111111010010010101111;
        x_t[47] = 26'b11111111110100111011000100;
        x_t[48] = 26'b11111111110000111111001111;
        x_t[49] = 26'b11111111101111001110001001;
        x_t[50] = 26'b11111111101110000101100101;
        x_t[51] = 26'b11111111101101101110111000;
        x_t[52] = 26'b11111111101111100001010010;
        x_t[53] = 26'b11111111110011010111111010;
        x_t[54] = 26'b11111111110100010101000010;
        x_t[55] = 26'b11111111110001100010001010;
        x_t[56] = 26'b11111111101110000101001110;
        x_t[57] = 26'b11111111110010110011100110;
        x_t[58] = 26'b11111111110000011010110110;
        x_t[59] = 26'b11111111110010111000001011;
        x_t[60] = 26'b11111111101011010101110011;
        x_t[61] = 26'b11111111101000101011101010;
        x_t[62] = 26'b11111111100101100111000001;
        x_t[63] = 26'b11111111110001101101110000;
        
        h_t_prev[0] = 26'b11111111111011101000110111;
        h_t_prev[1] = 26'b11111111110011010011111100;
        h_t_prev[2] = 26'b11111111101010110110111101;
        h_t_prev[3] = 26'b11111111100110110001010010;
        h_t_prev[4] = 26'b11111111100110010111010011;
        h_t_prev[5] = 26'b11111111100100110010111010;
        h_t_prev[6] = 26'b11111111101001101000001011;
        h_t_prev[7] = 26'b00000000000000010110100110;
        h_t_prev[8] = 26'b11111111101111111111000100;
        h_t_prev[9] = 26'b11111111101101101000110000;
        h_t_prev[10] = 26'b11111111101100001010010011;
        h_t_prev[11] = 26'b11111111100100100011101000;
        h_t_prev[12] = 26'b11111111101000000011110010;
        h_t_prev[13] = 26'b11111111100000001011111110;
        h_t_prev[14] = 26'b11111111111001000111001000;
        h_t_prev[15] = 26'b11111111110001100010111000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 56 timeout!");
                $fdisplay(fd_cycles, "Test Vector  56: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  56: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 56");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 57
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111111011000001011010;
        x_t[1] = 26'b11111111101111101001000001;
        x_t[2] = 26'b11111111100111110100101111;
        x_t[3] = 26'b11111111100011011100100101;
        x_t[4] = 26'b11111111100100001001110110;
        x_t[5] = 26'b11111111100101001001000110;
        x_t[6] = 26'b11111111101100010110011100;
        x_t[7] = 26'b00000000000000000010001111;
        x_t[8] = 26'b11111111101101000101011010;
        x_t[9] = 26'b11111111101100000100100010;
        x_t[10] = 26'b11111111101010010100111000;
        x_t[11] = 26'b11111111100100100011101000;
        x_t[12] = 26'b11111111101001001010000001;
        x_t[13] = 26'b11111111100110001001100100;
        x_t[14] = 26'b11111111111000011100111100;
        x_t[15] = 26'b11111111110010001011100100;
        x_t[16] = 26'b11111111101110000111101101;
        x_t[17] = 26'b11111111101010010101111101;
        x_t[18] = 26'b11111111101101101110110110;
        x_t[19] = 26'b11111111101100011010101100;
        x_t[20] = 26'b11111111101001011011011111;
        x_t[21] = 26'b11111111110110001001011101;
        x_t[22] = 26'b11111111110000100010001101;
        x_t[23] = 26'b11111111101111111111010010;
        x_t[24] = 26'b00000000000000010011110000;
        x_t[25] = 26'b00000000000000001101011101;
        x_t[26] = 26'b11111111100101110100111000;
        x_t[27] = 26'b11111111100101110100001101;
        x_t[28] = 26'b11111111101111011111100010;
        x_t[29] = 26'b00000000000001010110001110;
        x_t[30] = 26'b11111111111011001110110000;
        x_t[31] = 26'b11111111100111010010001011;
        x_t[32] = 26'b11111111100110010100100101;
        x_t[33] = 26'b11111111100100000011000101;
        x_t[34] = 26'b11111111100011010101010011;
        x_t[35] = 26'b11111111101001000011110000;
        x_t[36] = 26'b11111111101001100011000111;
        x_t[37] = 26'b11111111111100101111100010;
        x_t[38] = 26'b11111111111101011011111011;
        x_t[39] = 26'b11111111101100100110010100;
        x_t[40] = 26'b11111111111110011111001101;
        x_t[41] = 26'b11111111101111100110101100;
        x_t[42] = 26'b11111111111010101101100000;
        x_t[43] = 26'b11111111101110101000111011;
        x_t[44] = 26'b00000000000000111100001100;
        x_t[45] = 26'b11111111110100010111010110;
        x_t[46] = 26'b11111111111001010100100101;
        x_t[47] = 26'b11111111111000000010000000;
        x_t[48] = 26'b11111111110011010111101101;
        x_t[49] = 26'b11111111110100011011110000;
        x_t[50] = 26'b11111111110001101001101001;
        x_t[51] = 26'b11111111110101111000011110;
        x_t[52] = 26'b11111111110111110101010100;
        x_t[53] = 26'b11111111111101011101101110;
        x_t[54] = 26'b11111111111110000100010011;
        x_t[55] = 26'b11111111111000000000011111;
        x_t[56] = 26'b11111111110100110010111000;
        x_t[57] = 26'b11111111111010010001000100;
        x_t[58] = 26'b11111111111111101011111001;
        x_t[59] = 26'b00000000000110000111101110;
        x_t[60] = 26'b11111111110001110011110101;
        x_t[61] = 26'b11111111110011000001110100;
        x_t[62] = 26'b11111111110100011001111001;
        x_t[63] = 26'b11111111111100011100010000;
        
        h_t_prev[0] = 26'b11111111111011000001011010;
        h_t_prev[1] = 26'b11111111101111101001000001;
        h_t_prev[2] = 26'b11111111100111110100101111;
        h_t_prev[3] = 26'b11111111100011011100100101;
        h_t_prev[4] = 26'b11111111100100001001110110;
        h_t_prev[5] = 26'b11111111100101001001000110;
        h_t_prev[6] = 26'b11111111101100010110011100;
        h_t_prev[7] = 26'b00000000000000000010001111;
        h_t_prev[8] = 26'b11111111101101000101011010;
        h_t_prev[9] = 26'b11111111101100000100100010;
        h_t_prev[10] = 26'b11111111101010010100111000;
        h_t_prev[11] = 26'b11111111100100100011101000;
        h_t_prev[12] = 26'b11111111101001001010000001;
        h_t_prev[13] = 26'b11111111100110001001100100;
        h_t_prev[14] = 26'b11111111111000011100111100;
        h_t_prev[15] = 26'b11111111110010001011100100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 57 timeout!");
                $fdisplay(fd_cycles, "Test Vector  57: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  57: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 57");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 58
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111110111010100101000;
        x_t[1] = 26'b11111111101101011111111110;
        x_t[2] = 26'b11111111100110010011100111;
        x_t[3] = 26'b11111111100001101000100100;
        x_t[4] = 26'b11111111100100001001110110;
        x_t[5] = 26'b11111111100100011100101110;
        x_t[6] = 26'b11111111101011111101100010;
        x_t[7] = 26'b11111111111101011111010111;
        x_t[8] = 26'b11111111101100110000110010;
        x_t[9] = 26'b11111111101100000100100010;
        x_t[10] = 26'b11111111101011100011001010;
        x_t[11] = 26'b11111111100101100000110001;
        x_t[12] = 26'b11111111101010100111101011;
        x_t[13] = 26'b11111111100111110110100110;
        x_t[14] = 26'b11111111110111110010110000;
        x_t[15] = 26'b11111111110011110001010001;
        x_t[16] = 26'b11111111110000111010001010;
        x_t[17] = 26'b11111111101011100100111010;
        x_t[18] = 26'b11111111110001010110110001;
        x_t[19] = 26'b11111111110000100010010011;
        x_t[20] = 26'b11111111101100111100101111;
        x_t[21] = 26'b11111111110100110001000011;
        x_t[22] = 26'b11111111101101110000100000;
        x_t[23] = 26'b11111111101101010001010001;
        x_t[24] = 26'b11111111111101101001001111;
        x_t[25] = 26'b11111111111101011111011010;
        x_t[26] = 26'b11111111100010101010000111;
        x_t[27] = 26'b11111111100010011000000110;
        x_t[28] = 26'b11111111101100100010100111;
        x_t[29] = 26'b11111111111011101000001100;
        x_t[30] = 26'b11111111110111000101010111;
        x_t[31] = 26'b11111111100011101011100001;
        x_t[32] = 26'b11111111100011110001000010;
        x_t[33] = 26'b11111111100000110111100011;
        x_t[34] = 26'b11111111100000111100111001;
        x_t[35] = 26'b11111111100101010110111001;
        x_t[36] = 26'b11111111100100111000111011;
        x_t[37] = 26'b11111111110111001000110001;
        x_t[38] = 26'b11111111111100110011100110;
        x_t[39] = 26'b11111111100101101101010111;
        x_t[40] = 26'b11111111111001101110110111;
        x_t[41] = 26'b11111111011011100111000100;
        x_t[42] = 26'b11111111111011110100101001;
        x_t[43] = 26'b11111111110100110011111001;
        x_t[44] = 26'b00000000000000100101110110;
        x_t[45] = 26'b11111111111101000100011110;
        x_t[46] = 26'b11111111111000111111110111;
        x_t[47] = 26'b11111111111010100001001001;
        x_t[48] = 26'b11111111111000001000101001;
        x_t[49] = 26'b11111111111001000100010010;
        x_t[50] = 26'b11111111110100111010101100;
        x_t[51] = 26'b11111111111110010101011001;
        x_t[52] = 26'b00000000000001000110101110;
        x_t[53] = 26'b00000000001000111100100111;
        x_t[54] = 26'b00000000001100101011001101;
        x_t[55] = 26'b11111111111110110000000100;
        x_t[56] = 26'b11111111111011100000100011;
        x_t[57] = 26'b00000000000001011101011110;
        x_t[58] = 26'b00000000001111011111110110;
        x_t[59] = 26'b00000000011010000110101001;
        x_t[60] = 26'b11111111111100010110100100;
        x_t[61] = 26'b00000000000011010100101100;
        x_t[62] = 26'b00000000001011110000001100;
        x_t[63] = 26'b00000000001001111010110010;
        
        h_t_prev[0] = 26'b11111111110111010100101000;
        h_t_prev[1] = 26'b11111111101101011111111110;
        h_t_prev[2] = 26'b11111111100110010011100111;
        h_t_prev[3] = 26'b11111111100001101000100100;
        h_t_prev[4] = 26'b11111111100100001001110110;
        h_t_prev[5] = 26'b11111111100100011100101110;
        h_t_prev[6] = 26'b11111111101011111101100010;
        h_t_prev[7] = 26'b11111111111101011111010111;
        h_t_prev[8] = 26'b11111111101100110000110010;
        h_t_prev[9] = 26'b11111111101100000100100010;
        h_t_prev[10] = 26'b11111111101011100011001010;
        h_t_prev[11] = 26'b11111111100101100000110001;
        h_t_prev[12] = 26'b11111111101010100111101011;
        h_t_prev[13] = 26'b11111111100111110110100110;
        h_t_prev[14] = 26'b11111111110111110010110000;
        h_t_prev[15] = 26'b11111111110011110001010001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 58 timeout!");
                $fdisplay(fd_cycles, "Test Vector  58: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  58: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 58");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 59
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111110111000000111001;
        x_t[1] = 26'b11111111101111111100100110;
        x_t[2] = 26'b11111111100110100111000010;
        x_t[3] = 26'b11111111100001010101001110;
        x_t[4] = 26'b11111111100011001101001110;
        x_t[5] = 26'b11111111100010101101110001;
        x_t[6] = 26'b11111111100110100001000001;
        x_t[7] = 26'b11111111111101001011000000;
        x_t[8] = 26'b11111111101111010101110100;
        x_t[9] = 26'b11111111101101010100101101;
        x_t[10] = 26'b11111111101100110001011100;
        x_t[11] = 26'b11111111100111000110101100;
        x_t[12] = 26'b11111111101001100001011100;
        x_t[13] = 26'b11111111100010010100010000;
        x_t[14] = 26'b11111111111001110001010100;
        x_t[15] = 26'b11111111110101111111101010;
        x_t[16] = 26'b11111111110011101100100110;
        x_t[17] = 26'b11111111101101000111100111;
        x_t[18] = 26'b11111111110011010101010001;
        x_t[19] = 26'b11111111110011010010000010;
        x_t[20] = 26'b11111111110000000100111101;
        x_t[21] = 26'b11111111110111100001110111;
        x_t[22] = 26'b11111111110000100010001101;
        x_t[23] = 26'b11111111110000010110011111;
        x_t[24] = 26'b00000000000000101100000111;
        x_t[25] = 26'b00000000000000001101011101;
        x_t[26] = 26'b11111111100110010110101011;
        x_t[27] = 26'b11111111100101100100011111;
        x_t[28] = 26'b11111111101110100000100011;
        x_t[29] = 26'b11111111111111110010011001;
        x_t[30] = 26'b11111111111010101111100010;
        x_t[31] = 26'b11111111100111110101101010;
        x_t[32] = 26'b11111111101000100101111101;
        x_t[33] = 26'b11111111100011011110000101;
        x_t[34] = 26'b11111111100011000010010000;
        x_t[35] = 26'b11111111101000110000000001;
        x_t[36] = 26'b11111111100101001100110011;
        x_t[37] = 26'b11111111110101100110111011;
        x_t[38] = 26'b00000000000001110110010011;
        x_t[39] = 26'b11111111100010111100111111;
        x_t[40] = 26'b00000000000010100100000100;
        x_t[41] = 26'b11111111011100000010111000;
        x_t[42] = 26'b00000000001010010001100101;
        x_t[43] = 26'b11111111110000101100100101;
        x_t[44] = 26'b00000000001010010111011101;
        x_t[45] = 26'b00000000001000001100011000;
        x_t[46] = 26'b00000000000001101111010111;
        x_t[47] = 26'b00000000000000101111000000;
        x_t[48] = 26'b11111111111100100110100010;
        x_t[49] = 26'b11111111111010001110011011;
        x_t[50] = 26'b11111111110101100000101101;
        x_t[51] = 26'b00000000000000101111111100;
        x_t[52] = 26'b00000000000100111100010001;
        x_t[53] = 26'b00000000001110110111001101;
        x_t[54] = 26'b00000000010100001010101001;
        x_t[55] = 26'b00000000000111101001110000;
        x_t[56] = 26'b00000000000000111000010010;
        x_t[57] = 26'b00000000000001101110100001;
        x_t[58] = 26'b00000000010100011001111010;
        x_t[59] = 26'b00000000100001110000000110;
        x_t[60] = 26'b00000000000111001000101000;
        x_t[61] = 26'b00000000001111111111110101;
        x_t[62] = 26'b00000000011110011110100101;
        x_t[63] = 26'b00000000010100010111101100;
        
        h_t_prev[0] = 26'b11111111110111000000111001;
        h_t_prev[1] = 26'b11111111101111111100100110;
        h_t_prev[2] = 26'b11111111100110100111000010;
        h_t_prev[3] = 26'b11111111100001010101001110;
        h_t_prev[4] = 26'b11111111100011001101001110;
        h_t_prev[5] = 26'b11111111100010101101110001;
        h_t_prev[6] = 26'b11111111100110100001000001;
        h_t_prev[7] = 26'b11111111111101001011000000;
        h_t_prev[8] = 26'b11111111101111010101110100;
        h_t_prev[9] = 26'b11111111101101010100101101;
        h_t_prev[10] = 26'b11111111101100110001011100;
        h_t_prev[11] = 26'b11111111100111000110101100;
        h_t_prev[12] = 26'b11111111101001100001011100;
        h_t_prev[13] = 26'b11111111100010010100010000;
        h_t_prev[14] = 26'b11111111111001110001010100;
        h_t_prev[15] = 26'b11111111110101111111101010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 59 timeout!");
                $fdisplay(fd_cycles, "Test Vector  59: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  59: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 59");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 60
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111111110101110001011;
        x_t[1] = 26'b11111111110111111001100111;
        x_t[2] = 26'b11111111101100111110111011;
        x_t[3] = 26'b11111111100111010111111101;
        x_t[4] = 26'b11111111100101101110111000;
        x_t[5] = 26'b11111111100100011100101110;
        x_t[6] = 26'b11111111101001001111010010;
        x_t[7] = 26'b00000000000100001010111001;
        x_t[8] = 26'b11111111110100110100100000;
        x_t[9] = 26'b11111111110001000101001111;
        x_t[10] = 26'b11111111101111100001100100;
        x_t[11] = 26'b11111111101000101100100111;
        x_t[12] = 26'b11111111101100011100101111;
        x_t[13] = 26'b11111111100111011011010110;
        x_t[14] = 26'b00000000000000000010000110;
        x_t[15] = 26'b11111111111000001110000011;
        x_t[16] = 26'b11111111110100010100010000;
        x_t[17] = 26'b11111111101110010110100101;
        x_t[18] = 26'b11111111110100010100100001;
        x_t[19] = 26'b11111111110110000001110001;
        x_t[20] = 26'b11111111110101001010010100;
        x_t[21] = 26'b11111111111000101111001110;
        x_t[22] = 26'b11111111110000001000110100;
        x_t[23] = 26'b11111111101111010000111000;
        x_t[24] = 26'b00000000000001110101001100;
        x_t[25] = 26'b00000000000001001011100111;
        x_t[26] = 26'b11111111100111111100000011;
        x_t[27] = 26'b11111111100100000110001010;
        x_t[28] = 26'b11111111101011110000001110;
        x_t[29] = 26'b00000000000010011000110010;
        x_t[30] = 26'b11111111111101011011010000;
        x_t[31] = 26'b11111111100111000000011100;
        x_t[32] = 26'b11111111101011011011101011;
        x_t[33] = 26'b11111111100110000100100110;
        x_t[34] = 26'b11111111100011000010010000;
        x_t[35] = 26'b11111111101001000011110000;
        x_t[36] = 26'b11111111100010000110000001;
        x_t[37] = 26'b11111111110100000101000101;
        x_t[38] = 26'b00000000000011000110111111;
        x_t[39] = 26'b11111111100011011010011000;
        x_t[40] = 26'b00000000001001010110110110;
        x_t[41] = 26'b11111111100100010011011011;
        x_t[42] = 26'b00000000001000110010101110;
        x_t[43] = 26'b11111111101111010100110100;
        x_t[44] = 26'b00000000001011000100001001;
        x_t[45] = 26'b11111111111110000010011000;
        x_t[46] = 26'b00000000000100111110100101;
        x_t[47] = 26'b00000000000001101010101011;
        x_t[48] = 26'b11111111111100000000011010;
        x_t[49] = 26'b11111111111001000100010010;
        x_t[50] = 26'b11111111110100000001101011;
        x_t[51] = 26'b00000000000000011100101000;
        x_t[52] = 26'b00000000000101100101001101;
        x_t[53] = 26'b00000000001110110111001101;
        x_t[54] = 26'b00000000010010101010110000;
        x_t[55] = 26'b00000000001010100111101010;
        x_t[56] = 26'b00000000000010001110001110;
        x_t[57] = 26'b00000000000000111011010111;
        x_t[58] = 26'b00000000010101011111101100;
        x_t[59] = 26'b00000000100011011110101000;
        x_t[60] = 26'b00000000001101100110101010;
        x_t[61] = 26'b00000000010011100111100101;
        x_t[62] = 26'b00000000100100111100110101;
        x_t[63] = 26'b00000000010101101111101101;
        
        h_t_prev[0] = 26'b11111111111110101110001011;
        h_t_prev[1] = 26'b11111111110111111001100111;
        h_t_prev[2] = 26'b11111111101100111110111011;
        h_t_prev[3] = 26'b11111111100111010111111101;
        h_t_prev[4] = 26'b11111111100101101110111000;
        h_t_prev[5] = 26'b11111111100100011100101110;
        h_t_prev[6] = 26'b11111111101001001111010010;
        h_t_prev[7] = 26'b00000000000100001010111001;
        h_t_prev[8] = 26'b11111111110100110100100000;
        h_t_prev[9] = 26'b11111111110001000101001111;
        h_t_prev[10] = 26'b11111111101111100001100100;
        h_t_prev[11] = 26'b11111111101000101100100111;
        h_t_prev[12] = 26'b11111111101100011100101111;
        h_t_prev[13] = 26'b11111111100111011011010110;
        h_t_prev[14] = 26'b00000000000000000010000110;
        h_t_prev[15] = 26'b11111111111000001110000011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 60 timeout!");
                $fdisplay(fd_cycles, "Test Vector  60: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  60: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 60");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 61
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111111110011010011100;
        x_t[1] = 26'b11111111110101011100111111;
        x_t[2] = 26'b11111111101011011101110011;
        x_t[3] = 26'b11111111100100111101010000;
        x_t[4] = 26'b11111111100010100100110011;
        x_t[5] = 26'b11111111100000111110110101;
        x_t[6] = 26'b11111111100100001011101010;
        x_t[7] = 26'b00000000000011001101110100;
        x_t[8] = 26'b11111111110010111000101111;
        x_t[9] = 26'b11111111101111110101000100;
        x_t[10] = 26'b11111111101111100001100100;
        x_t[11] = 26'b11111111100110011101111011;
        x_t[12] = 26'b11111111101011101101111010;
        x_t[13] = 26'b11111111100111110110100110;
        x_t[14] = 26'b00000000000000010111001100;
        x_t[15] = 26'b11111111110110101000010110;
        x_t[16] = 26'b11111111110100000000011011;
        x_t[17] = 26'b11111111101111100101100010;
        x_t[18] = 26'b11111111110110010011000001;
        x_t[19] = 26'b11111111111000000101100101;
        x_t[20] = 26'b11111111110111111001100000;
        x_t[21] = 26'b11111111110100001111111001;
        x_t[22] = 26'b11111111101010110010000111;
        x_t[23] = 26'b11111111101010000000011100;
        x_t[24] = 26'b11111111111110011001111101;
        x_t[25] = 26'b11111111111101101011110101;
        x_t[26] = 26'b11111111100010101010000111;
        x_t[27] = 26'b11111111011101011101101010;
        x_t[28] = 26'b11111111100111000001111100;
        x_t[29] = 26'b00000000000100111111001010;
        x_t[30] = 26'b11111111111001000010010000;
        x_t[31] = 26'b11111111100011101011100001;
        x_t[32] = 26'b11111111100111101111011100;
        x_t[33] = 26'b11111111100001101111000100;
        x_t[34] = 26'b11111111011101101011010100;
        x_t[35] = 26'b11111111100011001100101111;
        x_t[36] = 26'b11111111011110000011100101;
        x_t[37] = 26'b11111111110011010100001010;
        x_t[38] = 26'b00000000000101111100100001;
        x_t[39] = 26'b11111111011111101111001101;
        x_t[40] = 26'b00000000001010011000000100;
        x_t[41] = 26'b11111111100010111111111110;
        x_t[42] = 26'b00000000000110111100001001;
        x_t[43] = 26'b00000000001000000000101101;
        x_t[44] = 26'b00000000001111111100111101;
        x_t[45] = 26'b00000000000111001110011110;
        x_t[46] = 26'b00000000001101011001010111;
        x_t[47] = 26'b00000000001001001000000111;
        x_t[48] = 26'b00000000000001111101100110;
        x_t[49] = 26'b11111111111111011100000001;
        x_t[50] = 26'b11111111111011001001110100;
        x_t[51] = 26'b00000000000111011000111100;
        x_t[52] = 26'b00000000001011111110011101;
        x_t[53] = 26'b00000000010101110100100101;
        x_t[54] = 26'b00000000011001011010001111;
        x_t[55] = 26'b00000000010100010101001001;
        x_t[56] = 26'b00000000001010110100001100;
        x_t[57] = 26'b00000000000111010100101000;
        x_t[58] = 26'b00000000011010011001110000;
        x_t[59] = 26'b00000000100101011100111100;
        x_t[60] = 26'b00000000010011000111010111;
        x_t[61] = 26'b00000000010100001000101100;
        x_t[62] = 26'b00000000100100010000011101;
        x_t[63] = 26'b00000000010110100100100001;
        
        h_t_prev[0] = 26'b11111111111110011010011100;
        h_t_prev[1] = 26'b11111111110101011100111111;
        h_t_prev[2] = 26'b11111111101011011101110011;
        h_t_prev[3] = 26'b11111111100100111101010000;
        h_t_prev[4] = 26'b11111111100010100100110011;
        h_t_prev[5] = 26'b11111111100000111110110101;
        h_t_prev[6] = 26'b11111111100100001011101010;
        h_t_prev[7] = 26'b00000000000011001101110100;
        h_t_prev[8] = 26'b11111111110010111000101111;
        h_t_prev[9] = 26'b11111111101111110101000100;
        h_t_prev[10] = 26'b11111111101111100001100100;
        h_t_prev[11] = 26'b11111111100110011101111011;
        h_t_prev[12] = 26'b11111111101011101101111010;
        h_t_prev[13] = 26'b11111111100111110110100110;
        h_t_prev[14] = 26'b00000000000000010111001100;
        h_t_prev[15] = 26'b11111111110110101000010110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 61 timeout!");
                $fdisplay(fd_cycles, "Test Vector  61: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  61: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 61");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 62
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000010011010111100;
        x_t[1] = 26'b11111111111001000111111010;
        x_t[2] = 26'b11111111101101111001001100;
        x_t[3] = 26'b11111111100010110101111010;
        x_t[4] = 26'b11111111100001111100011001;
        x_t[5] = 26'b11111111100000111110110101;
        x_t[6] = 26'b11111111100111010010110100;
        x_t[7] = 26'b00000000001010100010000100;
        x_t[8] = 26'b11111111111001101001111100;
        x_t[9] = 26'b11111111110110011010000000;
        x_t[10] = 26'b11111111110101000001110100;
        x_t[11] = 26'b11111111101001111110001001;
        x_t[12] = 26'b11111111101101100010111110;
        x_t[13] = 26'b11111111101110101010101101;
        x_t[14] = 26'b00000000001001100101110100;
        x_t[15] = 26'b00000000000000110011010001;
        x_t[16] = 26'b11111111111100111111011011;
        x_t[17] = 26'b11111111110110111111010010;
        x_t[18] = 26'b11111111111100111000101101;
        x_t[19] = 26'b11111111111101111011000001;
        x_t[20] = 26'b11111111111110111100000000;
        x_t[21] = 26'b11111111110101011101010000;
        x_t[22] = 26'b11111111101011111110010001;
        x_t[23] = 26'b11111111101100000000000011;
        x_t[24] = 26'b11111111111111100011000010;
        x_t[25] = 26'b11111111111110101010000000;
        x_t[26] = 26'b11111111100010111011000001;
        x_t[27] = 26'b11111111011110001100110101;
        x_t[28] = 26'b11111111101001100101101011;
        x_t[29] = 26'b00000000000100011101111000;
        x_t[30] = 26'b11111111111010111111001001;
        x_t[31] = 26'b11111111100011011001110010;
        x_t[32] = 26'b11111111101001001010010011;
        x_t[33] = 26'b11111111100001001010000011;
        x_t[34] = 26'b11111111011101000101001101;
        x_t[35] = 26'b11111111100011001100101111;
        x_t[36] = 26'b11111111011111111010110111;
        x_t[37] = 26'b11111111110111111001101100;
        x_t[38] = 26'b00000000001000011101111000;
        x_t[39] = 26'b11111111100100010101001011;
        x_t[40] = 26'b00000000000111101010001001;
        x_t[41] = 26'b11111111100100101111001111;
        x_t[42] = 26'b00000000010010000011101000;
        x_t[43] = 26'b11111111111010111110111000;
        x_t[44] = 26'b00000000011011000111111100;
        x_t[45] = 26'b00000000001101100000110110;
        x_t[46] = 26'b00000000011010101010111111;
        x_t[47] = 26'b00000000010000111001011011;
        x_t[48] = 26'b00000000000111100111101101;
        x_t[49] = 26'b00000000000100111100001010;
        x_t[50] = 26'b11111111111111010011111000;
        x_t[51] = 26'b00000000001000010010111001;
        x_t[52] = 26'b00000000001011000001000100;
        x_t[53] = 26'b00000000010100000101001111;
        x_t[54] = 26'b00000000010111001010011010;
        x_t[55] = 26'b00000000011100001001110001;
        x_t[56] = 26'b00000000010000101110010011;
        x_t[57] = 26'b00000000001010010000001100;
        x_t[58] = 26'b00000000010111011001110101;
        x_t[59] = 26'b00000000100000010001010111;
        x_t[60] = 26'b00000000011001000110101111;
        x_t[61] = 26'b00000000010101011011011101;
        x_t[62] = 26'b00000000100001101101101101;
        x_t[63] = 26'b00000000011011110010111101;
        
        h_t_prev[0] = 26'b00000000000010011010111100;
        h_t_prev[1] = 26'b11111111111001000111111010;
        h_t_prev[2] = 26'b11111111101101111001001100;
        h_t_prev[3] = 26'b11111111100010110101111010;
        h_t_prev[4] = 26'b11111111100001111100011001;
        h_t_prev[5] = 26'b11111111100000111110110101;
        h_t_prev[6] = 26'b11111111100111010010110100;
        h_t_prev[7] = 26'b00000000001010100010000100;
        h_t_prev[8] = 26'b11111111111001101001111100;
        h_t_prev[9] = 26'b11111111110110011010000000;
        h_t_prev[10] = 26'b11111111110101000001110100;
        h_t_prev[11] = 26'b11111111101001111110001001;
        h_t_prev[12] = 26'b11111111101101100010111110;
        h_t_prev[13] = 26'b11111111101110101010101101;
        h_t_prev[14] = 26'b00000000001001100101110100;
        h_t_prev[15] = 26'b00000000000000110011010001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 62 timeout!");
                $fdisplay(fd_cycles, "Test Vector  62: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  62: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 62");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 63
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000000010000110101;
        x_t[1] = 26'b11111111111011010000111101;
        x_t[2] = 26'b11111111110000010100100101;
        x_t[3] = 26'b11111111100101010000100110;
        x_t[4] = 26'b11111111100000010111010110;
        x_t[5] = 26'b11111111011100110100100101;
        x_t[6] = 26'b11111111100100111101011100;
        x_t[7] = 26'b00000000001010001101101101;
        x_t[8] = 26'b11111111111010100111110101;
        x_t[9] = 26'b11111111111001001110011001;
        x_t[10] = 26'b11111111110101010101011001;
        x_t[11] = 26'b11111111100110001001100010;
        x_t[12] = 26'b11111111100101011111111001;
        x_t[13] = 26'b11111111100111110110100110;
        x_t[14] = 26'b00000000001101111000000011;
        x_t[15] = 26'b00000000000010101101010100;
        x_t[16] = 26'b11111111111110001110101111;
        x_t[17] = 26'b11111111110111100110110001;
        x_t[18] = 26'b11111111111010100101000111;
        x_t[19] = 26'b11111111111000011011100011;
        x_t[20] = 26'b11111111110110101110011011;
        x_t[21] = 26'b11111111110111100001110111;
        x_t[22] = 26'b11111111101110001001111001;
        x_t[23] = 26'b11111111101101101000011110;
        x_t[24] = 26'b00000000000001110101001100;
        x_t[25] = 26'b00000000000000111111001011;
        x_t[26] = 26'b11111111100101000010001100;
        x_t[27] = 26'b11111111011110111011111111;
        x_t[28] = 26'b11111111100111011011001000;
        x_t[29] = 26'b00000000000111010100111001;
        x_t[30] = 26'b11111111111101001011101000;
        x_t[31] = 26'b11111111100101000100001111;
        x_t[32] = 26'b11111111101100100100010111;
        x_t[33] = 26'b11111111100100111010100101;
        x_t[34] = 26'b11111111100000000011101111;
        x_t[35] = 26'b11111111100101010110111001;
        x_t[36] = 26'b11111111100000100010100111;
        x_t[37] = 26'b11111111111000001010000000;
        x_t[38] = 26'b00000000001001000110001101;
        x_t[39] = 26'b11111111100101001111111110;
        x_t[40] = 26'b00000000001101011011101101;
        x_t[41] = 26'b11111111101101110111011011;
        x_t[42] = 26'b00000000010101110000110011;
        x_t[43] = 26'b11111111110101011111110010;
        x_t[44] = 26'b00000000011011000111111100;
        x_t[45] = 26'b00000000000010011000111101;
        x_t[46] = 26'b00000000011000000101001101;
        x_t[47] = 26'b00000000010000100101100010;
        x_t[48] = 26'b00000000000110101110100010;
        x_t[49] = 26'b00000000000100101001101000;
        x_t[50] = 26'b11111111111101100001110110;
        x_t[51] = 26'b00000000000011011101110011;
        x_t[52] = 26'b00000000000101010000101111;
        x_t[53] = 26'b00000000001011011000100000;
        x_t[54] = 26'b00000000001110001011000110;
        x_t[55] = 26'b00000000011011010101111111;
        x_t[56] = 26'b00000000001111111010110000;
        x_t[57] = 26'b00000000001000011000110101;
        x_t[58] = 26'b00000000001111001110011010;
        x_t[59] = 26'b00000000010001011110000001;
        x_t[60] = 26'b00000000011010110010000101;
        x_t[61] = 26'b00000000010001010010100110;
        x_t[62] = 26'b00000000011001110110101011;
        x_t[63] = 26'b00000000011001110111101111;
        
        h_t_prev[0] = 26'b00000000000000010000110101;
        h_t_prev[1] = 26'b11111111111011010000111101;
        h_t_prev[2] = 26'b11111111110000010100100101;
        h_t_prev[3] = 26'b11111111100101010000100110;
        h_t_prev[4] = 26'b11111111100000010111010110;
        h_t_prev[5] = 26'b11111111011100110100100101;
        h_t_prev[6] = 26'b11111111100100111101011100;
        h_t_prev[7] = 26'b00000000001010001101101101;
        h_t_prev[8] = 26'b11111111111010100111110101;
        h_t_prev[9] = 26'b11111111111001001110011001;
        h_t_prev[10] = 26'b11111111110101010101011001;
        h_t_prev[11] = 26'b11111111100110001001100010;
        h_t_prev[12] = 26'b11111111100101011111111001;
        h_t_prev[13] = 26'b11111111100111110110100110;
        h_t_prev[14] = 26'b00000000001101111000000011;
        h_t_prev[15] = 26'b00000000000010101101010100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 63 timeout!");
                $fdisplay(fd_cycles, "Test Vector  63: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  63: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 63");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 64
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000011101001110111;
        x_t[1] = 26'b11111111111101011010000000;
        x_t[2] = 26'b11111111110001110101101100;
        x_t[3] = 26'b11111111100111010111111101;
        x_t[4] = 26'b11111111100011100001011011;
        x_t[5] = 26'b11111111011110100011100001;
        x_t[6] = 26'b11111111100101101111001111;
        x_t[7] = 26'b00000000001011011111001001;
        x_t[8] = 26'b11111111111010111100011110;
        x_t[9] = 26'b11111111111000010010010001;
        x_t[10] = 26'b11111111110010100101010001;
        x_t[11] = 26'b11111111100110001001100010;
        x_t[12] = 26'b11111111100011010011011011;
        x_t[13] = 26'b11111111100111110110100110;
        x_t[14] = 26'b00000000001011100100011001;
        x_t[15] = 26'b00000000000001011011111101;
        x_t[16] = 26'b11111111111100101011100110;
        x_t[17] = 26'b11111111110110101011100011;
        x_t[18] = 26'b11111111111000010001100010;
        x_t[19] = 26'b11111111110100101001111010;
        x_t[20] = 26'b11111111110010011011000111;
        x_t[21] = 26'b11111111111010010010101011;
        x_t[22] = 26'b11111111110001101110010111;
        x_t[23] = 26'b11111111110001011100000110;
        x_t[24] = 26'b00000000000100000111010101;
        x_t[25] = 26'b00000000000011010100010111;
        x_t[26] = 26'b11111111101000011101110110;
        x_t[27] = 26'b11111111100011100110101101;
        x_t[28] = 26'b11111111101110010011111101;
        x_t[29] = 26'b00000000001010001011111011;
        x_t[30] = 26'b11111111111101101010110111;
        x_t[31] = 26'b11111111101010000011100111;
        x_t[32] = 26'b11111111101100110110100010;
        x_t[33] = 26'b11111111100110101001100110;
        x_t[34] = 26'b11111111100011010101010011;
        x_t[35] = 26'b11111111101000001000100010;
        x_t[36] = 26'b11111111100011101001011010;
        x_t[37] = 26'b11111111111001111100001010;
        x_t[38] = 26'b00000000001100001111111010;
        x_t[39] = 26'b11111111101010010011010101;
        x_t[40] = 26'b00000000010100111001111101;
        x_t[41] = 26'b11111111110101101100001001;
        x_t[42] = 26'b00000000010110110111111100;
        x_t[43] = 26'b11111111110010000100010111;
        x_t[44] = 26'b00000000011010110001100110;
        x_t[45] = 26'b11111111111111000000010010;
        x_t[46] = 26'b00000000010100110101111111;
        x_t[47] = 26'b00000000001101011110100111;
        x_t[48] = 26'b00000000000101001111001111;
        x_t[49] = 26'b00000000000100000100100100;
        x_t[50] = 26'b11111111111110101101111000;
        x_t[51] = 26'b00000000000010100011110110;
        x_t[52] = 26'b00000000000011000001100000;
        x_t[53] = 26'b00000000000110001010011101;
        x_t[54] = 26'b00000000000110010011101100;
        x_t[55] = 26'b00000000011000000110110101;
        x_t[56] = 26'b00000000001101100000000100;
        x_t[57] = 26'b00000000001000000111110010;
        x_t[58] = 26'b00000000001010110111001111;
        x_t[59] = 26'b00000000001000010101110101;
        x_t[60] = 26'b00000000010111011011011001;
        x_t[61] = 26'b00000000001011000101010100;
        x_t[62] = 26'b00000000010001000100011110;
        x_t[63] = 26'b00000000010101101111101101;
        
        h_t_prev[0] = 26'b00000000000011101001110111;
        h_t_prev[1] = 26'b11111111111101011010000000;
        h_t_prev[2] = 26'b11111111110001110101101100;
        h_t_prev[3] = 26'b11111111100111010111111101;
        h_t_prev[4] = 26'b11111111100011100001011011;
        h_t_prev[5] = 26'b11111111011110100011100001;
        h_t_prev[6] = 26'b11111111100101101111001111;
        h_t_prev[7] = 26'b00000000001011011111001001;
        h_t_prev[8] = 26'b11111111111010111100011110;
        h_t_prev[9] = 26'b11111111111000010010010001;
        h_t_prev[10] = 26'b11111111110010100101010001;
        h_t_prev[11] = 26'b11111111100110001001100010;
        h_t_prev[12] = 26'b11111111100011010011011011;
        h_t_prev[13] = 26'b11111111100111110110100110;
        h_t_prev[14] = 26'b00000000001011100100011001;
        h_t_prev[15] = 26'b00000000000001011011111101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 64 timeout!");
                $fdisplay(fd_cycles, "Test Vector  64: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  64: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 64");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 65
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111100100110100110001;
        x_t[1] = 26'b11111111101111000001110111;
        x_t[2] = 26'b11111111110000101000000000;
        x_t[3] = 26'b11111111111010011010001000;
        x_t[4] = 26'b11111111111100011101110111;
        x_t[5] = 26'b11111111111100000001100001;
        x_t[6] = 26'b11111111110100001000010100;
        x_t[7] = 26'b11111111101101100101011100;
        x_t[8] = 26'b11111111110110000111000010;
        x_t[9] = 26'b11111111111001100010011100;
        x_t[10] = 26'b11111111111101100101110001;
        x_t[11] = 26'b11111111111111111100100111;
        x_t[12] = 26'b00000000000001101010101011;
        x_t[13] = 26'b11111111111100101110001101;
        x_t[14] = 26'b11111111110110001001010010;
        x_t[15] = 26'b11111111111010001000000110;
        x_t[16] = 26'b11111111111011110000000111;
        x_t[17] = 26'b00000000000001110010001100;
        x_t[18] = 26'b00000000000010011111001000;
        x_t[19] = 26'b00000000000100011100011001;
        x_t[20] = 26'b00000000000101111110100000;
        x_t[21] = 26'b11111111100101111010101010;
        x_t[22] = 26'b11111111100100101000101001;
        x_t[23] = 26'b11111111101001000110011011;
        x_t[24] = 26'b11111111100100001001001101;
        x_t[25] = 26'b11111111100100011011101110;
        x_t[26] = 26'b11111111101011000110110100;
        x_t[27] = 26'b11111111101100011100101100;
        x_t[28] = 26'b11111111101010111101110110;
        x_t[29] = 26'b11111111100010011010010011;
        x_t[30] = 26'b11111111101001011011001011;
        x_t[31] = 26'b11111111101101101010010001;
        x_t[32] = 26'b11111111101110100011100100;
        x_t[33] = 26'b11111111110001101000101101;
        x_t[34] = 26'b11111111110101001100011100;
        x_t[35] = 26'b11111111110100011110000011;
        x_t[36] = 26'b11111111110011110011001001;
        x_t[37] = 26'b11111111110100110110000000;
        x_t[38] = 26'b11111111100101001010110111;
        x_t[39] = 26'b11111111110101010100110110;
        x_t[40] = 26'b11111111100111000011001110;
        x_t[41] = 26'b00000000000000000111110010;
        x_t[42] = 26'b11111111011110111010110001;
        x_t[43] = 26'b00000000000011001101100000;
        x_t[44] = 26'b11111111110000100010000011;
        x_t[45] = 26'b11111111111110000010011000;
        x_t[46] = 26'b11111111111110100000001001;
        x_t[47] = 26'b11111111111101111011111101;
        x_t[48] = 26'b00000000000001010111011110;
        x_t[49] = 26'b00000000000010010101010111;
        x_t[50] = 26'b00000000000010110111111100;
        x_t[51] = 26'b00000000001000111001100010;
        x_t[52] = 26'b00000000000101100101001101;
        x_t[53] = 26'b00000000001000010000000101;
        x_t[54] = 26'b00000000000101100011101111;
        x_t[55] = 26'b00000000000110010011011100;
        x_t[56] = 26'b00000000000110100001001101;
        x_t[57] = 26'b00000000001101111110111011;
        x_t[58] = 26'b00000000001101110111001010;
        x_t[59] = 26'b00000000001011000011100000;
        x_t[60] = 26'b00000000001110010100101011;
        x_t[61] = 26'b00000000010011010111000010;
        x_t[62] = 26'b00000000000101101111100001;
        x_t[63] = 26'b00000000001101001110000001;
        
        h_t_prev[0] = 26'b11111111100100110100110001;
        h_t_prev[1] = 26'b11111111101111000001110111;
        h_t_prev[2] = 26'b11111111110000101000000000;
        h_t_prev[3] = 26'b11111111111010011010001000;
        h_t_prev[4] = 26'b11111111111100011101110111;
        h_t_prev[5] = 26'b11111111111100000001100001;
        h_t_prev[6] = 26'b11111111110100001000010100;
        h_t_prev[7] = 26'b11111111101101100101011100;
        h_t_prev[8] = 26'b11111111110110000111000010;
        h_t_prev[9] = 26'b11111111111001100010011100;
        h_t_prev[10] = 26'b11111111111101100101110001;
        h_t_prev[11] = 26'b11111111111111111100100111;
        h_t_prev[12] = 26'b00000000000001101010101011;
        h_t_prev[13] = 26'b11111111111100101110001101;
        h_t_prev[14] = 26'b11111111110110001001010010;
        h_t_prev[15] = 26'b11111111111010001000000110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 65 timeout!");
                $fdisplay(fd_cycles, "Test Vector  65: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  65: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 65");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 66
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111100110111110111001;
        x_t[1] = 26'b11111111110010000101101001;
        x_t[2] = 26'b11111111110011101010001111;
        x_t[3] = 26'b11111111111010101101011101;
        x_t[4] = 26'b11111111111101011010011111;
        x_t[5] = 26'b11111111111111001001001101;
        x_t[6] = 26'b11111111111011111010001101;
        x_t[7] = 26'b11111111110001000101011000;
        x_t[8] = 26'b11111111111000101100000100;
        x_t[9] = 26'b11111111111010001010100010;
        x_t[10] = 26'b11111111111010110101101001;
        x_t[11] = 26'b11111111111111101000001110;
        x_t[12] = 26'b00000000000010011001100000;
        x_t[13] = 26'b00000000000010101011110011;
        x_t[14] = 26'b11111111110101011111000110;
        x_t[15] = 26'b11111111111001011111011011;
        x_t[16] = 26'b11111111111010110100101000;
        x_t[17] = 26'b11111111111101110001100100;
        x_t[18] = 26'b11111111111011111001011101;
        x_t[19] = 26'b11111111111111010010111001;
        x_t[20] = 26'b00000000000010011101010000;
        x_t[21] = 26'b11111111100100101101010011;
        x_t[22] = 26'b11111111100101110100110011;
        x_t[23] = 26'b11111111101011010001101001;
        x_t[24] = 26'b11111111100011100100101011;
        x_t[25] = 26'b11111111100100001111010010;
        x_t[26] = 26'b11111111101011101000100111;
        x_t[27] = 26'b11111111101111101001000101;
        x_t[28] = 26'b11111111101110101101001010;
        x_t[29] = 26'b11111111100011011100110110;
        x_t[30] = 26'b11111111101100010110100000;
        x_t[31] = 26'b11111111101111100110011101;
        x_t[32] = 26'b11111111101110100011100100;
        x_t[33] = 26'b11111111110001111011001101;
        x_t[34] = 26'b11111111110110000101100110;
        x_t[35] = 26'b11111111110101101101000000;
        x_t[36] = 26'b11111111111000110001001101;
        x_t[37] = 26'b11111111111000001010000000;
        x_t[38] = 26'b11111111100101110011001101;
        x_t[39] = 26'b11111111111110000011011000;
        x_t[40] = 26'b11111111101000000100011100;
        x_t[41] = 26'b00000000010100100011001110;
        x_t[42] = 26'b11111111011111101010001101;
        x_t[43] = 26'b11111111101111010100110100;
        x_t[44] = 26'b11111111101011111111100101;
        x_t[45] = 26'b11111111110101010101010000;
        x_t[46] = 26'b11111111111001101001010011;
        x_t[47] = 26'b11111111111100101100011001;
        x_t[48] = 26'b00000000000001101010100010;
        x_t[49] = 26'b00000000000000010011101000;
        x_t[50] = 26'b11111111111111000000111000;
        x_t[51] = 26'b00000000000011110001001000;
        x_t[52] = 26'b00000000000001000110101110;
        x_t[53] = 26'b00000000000101011101111011;
        x_t[54] = 26'b00000000000010111011111100;
        x_t[55] = 26'b00000000000101110000111010;
        x_t[56] = 26'b00000000000101011100011101;
        x_t[57] = 26'b00000000001100011000100111;
        x_t[58] = 26'b00000000001100001110011111;
        x_t[59] = 26'b00000000001010010100001001;
        x_t[60] = 26'b00000000001100011001111111;
        x_t[61] = 26'b00000000010001010010100110;
        x_t[62] = 26'b00000000000010101111001100;
        x_t[63] = 26'b00000000001011100100011010;
        
        h_t_prev[0] = 26'b11111111100110111110111001;
        h_t_prev[1] = 26'b11111111110010000101101001;
        h_t_prev[2] = 26'b11111111110011101010001111;
        h_t_prev[3] = 26'b11111111111010101101011101;
        h_t_prev[4] = 26'b11111111111101011010011111;
        h_t_prev[5] = 26'b11111111111111001001001101;
        h_t_prev[6] = 26'b11111111111011111010001101;
        h_t_prev[7] = 26'b11111111110001000101011000;
        h_t_prev[8] = 26'b11111111111000101100000100;
        h_t_prev[9] = 26'b11111111111010001010100010;
        h_t_prev[10] = 26'b11111111111010110101101001;
        h_t_prev[11] = 26'b11111111111111101000001110;
        h_t_prev[12] = 26'b00000000000010011001100000;
        h_t_prev[13] = 26'b00000000000010101011110011;
        h_t_prev[14] = 26'b11111111110101011111000110;
        h_t_prev[15] = 26'b11111111111001011111011011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 66 timeout!");
                $fdisplay(fd_cycles, "Test Vector  66: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  66: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 66");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 67
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111101010010111111100;
        x_t[1] = 26'b11111111110101011100111111;
        x_t[2] = 26'b11111111110101011110110001;
        x_t[3] = 26'b11111111111010000110110010;
        x_t[4] = 26'b11111111111100011101110111;
        x_t[5] = 26'b11111111111111001001001101;
        x_t[6] = 26'b00000000000000001100000010;
        x_t[7] = 26'b11111111110101100010011001;
        x_t[8] = 26'b11111111111011010001000110;
        x_t[9] = 26'b11111111111000111010010110;
        x_t[10] = 26'b11111111110111011110011000;
        x_t[11] = 26'b11111111111100001000000000;
        x_t[12] = 26'b00000000000000111011110110;
        x_t[13] = 26'b00000000000101001111010110;
        x_t[14] = 26'b11111111110111110010110000;
        x_t[15] = 26'b11111111111011101101110100;
        x_t[16] = 26'b11111111111010001100111110;
        x_t[17] = 26'b11111111111011111011001000;
        x_t[18] = 26'b11111111110111111100011100;
        x_t[19] = 26'b11111111111011110111001110;
        x_t[20] = 26'b00000000000010110110010010;
        x_t[21] = 26'b11111111101000010101011000;
        x_t[22] = 26'b11111111101000011001110011;
        x_t[23] = 26'b11111111101100111010000100;
        x_t[24] = 26'b11111111100111011000010000;
        x_t[25] = 26'b11111111100111100010101000;
        x_t[26] = 26'b11111111101101011110111001;
        x_t[27] = 26'b11111111110000011000001111;
        x_t[28] = 26'b11111111101110101101001010;
        x_t[29] = 26'b11111111101000101001100111;
        x_t[30] = 26'b11111111101100110101101110;
        x_t[31] = 26'b11111111110001100010101010;
        x_t[32] = 26'b11111111110001101011011101;
        x_t[33] = 26'b11111111110011101010001110;
        x_t[34] = 26'b11111111110110111110110000;
        x_t[35] = 26'b11111111110111001111101100;
        x_t[36] = 26'b11111111111000110001001101;
        x_t[37] = 26'b11111111110111001000110001;
        x_t[38] = 26'b11111111101101101011011100;
        x_t[39] = 26'b11111111111100001101110010;
        x_t[40] = 26'b11111111110000001110001011;
        x_t[41] = 26'b00000000001001101011110010;
        x_t[42] = 26'b11111111011101110011101000;
        x_t[43] = 26'b00000000000011001101100000;
        x_t[44] = 26'b11111111110001111011011011;
        x_t[45] = 26'b11111111111100000110100101;
        x_t[46] = 26'b11111111111111011110010011;
        x_t[47] = 26'b00000000000000011011000111;
        x_t[48] = 26'b00000000000100101001000111;
        x_t[49] = 26'b00000000000001110000010011;
        x_t[50] = 26'b11111111111111100110111001;
        x_t[51] = 26'b00000000000010100011110110;
        x_t[52] = 26'b00000000000000001001010101;
        x_t[53] = 26'b00000000000111001101010001;
        x_t[54] = 26'b00000000000111110011100100;
        x_t[55] = 26'b00000000000110110101111110;
        x_t[56] = 26'b00000000000110010000000001;
        x_t[57] = 26'b00000000001100101001101011;
        x_t[58] = 26'b00000000001101010100010001;
        x_t[59] = 26'b00000000001100010010011101;
        x_t[60] = 26'b00000000001011011100101001;
        x_t[61] = 26'b00000000010000100000111100;
        x_t[62] = 26'b00000000000010101111001100;
        x_t[63] = 26'b00000000001011110110000000;
        
        h_t_prev[0] = 26'b11111111101010010111111100;
        h_t_prev[1] = 26'b11111111110101011100111111;
        h_t_prev[2] = 26'b11111111110101011110110001;
        h_t_prev[3] = 26'b11111111111010000110110010;
        h_t_prev[4] = 26'b11111111111100011101110111;
        h_t_prev[5] = 26'b11111111111111001001001101;
        h_t_prev[6] = 26'b00000000000000001100000010;
        h_t_prev[7] = 26'b11111111110101100010011001;
        h_t_prev[8] = 26'b11111111111011010001000110;
        h_t_prev[9] = 26'b11111111111000111010010110;
        h_t_prev[10] = 26'b11111111110111011110011000;
        h_t_prev[11] = 26'b11111111111100001000000000;
        h_t_prev[12] = 26'b00000000000000111011110110;
        h_t_prev[13] = 26'b00000000000101001111010110;
        h_t_prev[14] = 26'b11111111110111110010110000;
        h_t_prev[15] = 26'b11111111111011101101110100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 67 timeout!");
                $fdisplay(fd_cycles, "Test Vector  67: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  67: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 67");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 68
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111110000110110010010;
        x_t[1] = 26'b11111111111001000111111010;
        x_t[2] = 26'b11111111110111100110101111;
        x_t[3] = 26'b11111111111010011010001000;
        x_t[4] = 26'b11111111111011110101011100;
        x_t[5] = 26'b11111111111101000100000101;
        x_t[6] = 26'b11111111111011111010001101;
        x_t[7] = 26'b11111111111010101000001001;
        x_t[8] = 26'b11111111111101100001100000;
        x_t[9] = 26'b11111111111010011110100101;
        x_t[10] = 26'b11111111111001111010111100;
        x_t[11] = 26'b11111111111001111001010100;
        x_t[12] = 26'b11111111111011110100000100;
        x_t[13] = 26'b11111111111001010100001001;
        x_t[14] = 26'b11111111111100011010000100;
        x_t[15] = 26'b11111111111100111111001011;
        x_t[16] = 26'b11111111111100000011111100;
        x_t[17] = 26'b11111111111100001110111000;
        x_t[18] = 26'b11111111110101101000110111;
        x_t[19] = 26'b11111111110111101111100111;
        x_t[20] = 26'b11111111111100001100110100;
        x_t[21] = 26'b11111111101000010101011000;
        x_t[22] = 26'b11111111100111110011101110;
        x_t[23] = 26'b11111111101100010111010000;
        x_t[24] = 26'b11111111100111111100110011;
        x_t[25] = 26'b11111111101000100000110010;
        x_t[26] = 26'b11111111101110000000101011;
        x_t[27] = 26'b11111111110000011000001111;
        x_t[28] = 26'b11111111101110101101001010;
        x_t[29] = 26'b11111111101001111100110011;
        x_t[30] = 26'b11111111101111100001011100;
        x_t[31] = 26'b11111111110000111111001011;
        x_t[32] = 26'b11111111110001111101101000;
        x_t[33] = 26'b11111111110011101010001110;
        x_t[34] = 26'b11111111110111010001110011;
        x_t[35] = 26'b11111111111000001010111001;
        x_t[36] = 26'b11111111110101111110010011;
        x_t[37] = 26'b11111111110110010111110110;
        x_t[38] = 26'b11111111101011110010011011;
        x_t[39] = 26'b11111111110010100100011110;
        x_t[40] = 26'b11111111101011011101110101;
        x_t[41] = 26'b11111111101000001101110010;
        x_t[42] = 26'b11111111100001111000100000;
        x_t[43] = 26'b11111111110011011100001000;
        x_t[44] = 26'b11111111110000100010000011;
        x_t[45] = 26'b11111111110101110100001100;
        x_t[46] = 26'b11111111111010111100001100;
        x_t[47] = 26'b11111111111011001000111011;
        x_t[48] = 26'b11111111111110101011111100;
        x_t[49] = 26'b11111111111101101100110101;
        x_t[50] = 26'b11111111111110000111110111;
        x_t[51] = 26'b11111111111111001111010110;
        x_t[52] = 26'b11111111111100010011110010;
        x_t[53] = 26'b00000000000000111100011011;
        x_t[54] = 26'b00000000000001011100000011;
        x_t[55] = 26'b11111111111100010100101100;
        x_t[56] = 26'b11111111111101011000110111;
        x_t[57] = 26'b00000000000110110010100001;
        x_t[58] = 26'b00000000000111000010111111;
        x_t[59] = 26'b00000000000110010111100001;
        x_t[60] = 26'b00000000000110001011010010;
        x_t[61] = 26'b00000000001011010101110111;
        x_t[62] = 26'b11111111111110110011101011;
        x_t[63] = 26'b00000000000101110010110000;
        
        h_t_prev[0] = 26'b11111111110000110110010010;
        h_t_prev[1] = 26'b11111111111001000111111010;
        h_t_prev[2] = 26'b11111111110111100110101111;
        h_t_prev[3] = 26'b11111111111010011010001000;
        h_t_prev[4] = 26'b11111111111011110101011100;
        h_t_prev[5] = 26'b11111111111101000100000101;
        h_t_prev[6] = 26'b11111111111011111010001101;
        h_t_prev[7] = 26'b11111111111010101000001001;
        h_t_prev[8] = 26'b11111111111101100001100000;
        h_t_prev[9] = 26'b11111111111010011110100101;
        h_t_prev[10] = 26'b11111111111001111010111100;
        h_t_prev[11] = 26'b11111111111001111001010100;
        h_t_prev[12] = 26'b11111111111011110100000100;
        h_t_prev[13] = 26'b11111111111001010100001001;
        h_t_prev[14] = 26'b11111111111100011010000100;
        h_t_prev[15] = 26'b11111111111100111111001011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 68 timeout!");
                $fdisplay(fd_cycles, "Test Vector  68: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  68: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 68");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 69
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111101111100111010111;
        x_t[1] = 26'b11111111110111100110000010;
        x_t[2] = 26'b11111111110110111111111000;
        x_t[3] = 26'b11111111111010011010001000;
        x_t[4] = 26'b11111111111011100001001111;
        x_t[5] = 26'b11111111111011101011010101;
        x_t[6] = 26'b11111111110110110110100101;
        x_t[7] = 26'b11111111110110001011000111;
        x_t[8] = 26'b11111111111011100101101110;
        x_t[9] = 26'b11111111111011011010101101;
        x_t[10] = 26'b11111111111100101011000100;
        x_t[11] = 26'b11111111111110000010010011;
        x_t[12] = 26'b11111111111011000101010000;
        x_t[13] = 26'b11111111110111100111000111;
        x_t[14] = 26'b11111111110100110100111010;
        x_t[15] = 26'b11111111111001011111011011;
        x_t[16] = 26'b11111111111100101011100110;
        x_t[17] = 26'b11111111111110000101010100;
        x_t[18] = 26'b11111111111010100101000111;
        x_t[19] = 26'b11111111111011001011010010;
        x_t[20] = 26'b11111111111110001001111101;
        x_t[21] = 26'b11111111100101101111100111;
        x_t[22] = 26'b11111111100100011011111101;
        x_t[23] = 26'b11111111101000011000000001;
        x_t[24] = 26'b11111111100100010101011001;
        x_t[25] = 26'b11111111100101011001111000;
        x_t[26] = 26'b11111111101100011011010011;
        x_t[27] = 26'b11111111101101101011010011;
        x_t[28] = 26'b11111111101011100011101000;
        x_t[29] = 26'b11111111100110110101001001;
        x_t[30] = 26'b11111111110010111011111111;
        x_t[31] = 26'b11111111110010000110001001;
        x_t[32] = 26'b11111111110001101011011101;
        x_t[33] = 26'b11111111110011111100101110;
        x_t[34] = 26'b11111111110111100100110111;
        x_t[35] = 26'b11111111110111001111101100;
        x_t[36] = 26'b11111111110011110011001001;
        x_t[37] = 26'b11111111111000001010000000;
        x_t[38] = 26'b11111111101101000011000110;
        x_t[39] = 26'b11111111110111001010011011;
        x_t[40] = 26'b11111111110010100110010110;
        x_t[41] = 26'b00000000001000011000010100;
        x_t[42] = 26'b11111111100001100000110010;
        x_t[43] = 26'b11111111110100001000000001;
        x_t[44] = 26'b11111111110001001110101111;
        x_t[45] = 26'b11111111111001101011110100;
        x_t[46] = 26'b11111111110110101110110011;
        x_t[47] = 26'b11111111111000101001110010;
        x_t[48] = 26'b11111111111111111000001011;
        x_t[49] = 26'b00000000000000100110001010;
        x_t[50] = 26'b00000000000011001010111101;
        x_t[51] = 26'b00000000000110011110111111;
        x_t[52] = 26'b00000000000100111100010001;
        x_t[53] = 26'b00000000000111001101010001;
        x_t[54] = 26'b00000000000111000011101000;
        x_t[55] = 26'b11111111111010001010100110;
        x_t[56] = 26'b11111111111101000111101011;
        x_t[57] = 26'b00000000001000101001111000;
        x_t[58] = 26'b00000000001011011010001001;
        x_t[59] = 26'b00000000001010010100001001;
        x_t[60] = 26'b00000000000000001011111011;
        x_t[61] = 26'b00000000000110001010110010;
        x_t[62] = 26'b11111111111100010000111011;
        x_t[63] = 26'b11111111111110111010101011;
        
        h_t_prev[0] = 26'b11111111101111100111010111;
        h_t_prev[1] = 26'b11111111110111100110000010;
        h_t_prev[2] = 26'b11111111110110111111111000;
        h_t_prev[3] = 26'b11111111111010011010001000;
        h_t_prev[4] = 26'b11111111111011100001001111;
        h_t_prev[5] = 26'b11111111111011101011010101;
        h_t_prev[6] = 26'b11111111110110110110100101;
        h_t_prev[7] = 26'b11111111110110001011000111;
        h_t_prev[8] = 26'b11111111111011100101101110;
        h_t_prev[9] = 26'b11111111111011011010101101;
        h_t_prev[10] = 26'b11111111111100101011000100;
        h_t_prev[11] = 26'b11111111111110000010010011;
        h_t_prev[12] = 26'b11111111111011000101010000;
        h_t_prev[13] = 26'b11111111110111100111000111;
        h_t_prev[14] = 26'b11111111110100110100111010;
        h_t_prev[15] = 26'b11111111111001011111011011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 69 timeout!");
                $fdisplay(fd_cycles, "Test Vector  69: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  69: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 69");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 70
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111101111111011000110;
        x_t[1] = 26'b11111111111000001101001011;
        x_t[2] = 26'b11111111111010000010000111;
        x_t[3] = 26'b11111111111111001111100000;
        x_t[4] = 26'b00000000000001001100111111;
        x_t[5] = 26'b00000000000001111010101110;
        x_t[6] = 26'b11111111111110101000011101;
        x_t[7] = 26'b11111111111001000010010110;
        x_t[8] = 26'b11111111111110001010110000;
        x_t[9] = 26'b11111111111110110111001100;
        x_t[10] = 26'b00000000000000000010010101;
        x_t[11] = 26'b00000000000010001011010010;
        x_t[12] = 26'b00000000000011110111001001;
        x_t[13] = 26'b00000000000010010000100010;
        x_t[14] = 26'b11111111110011110101101000;
        x_t[15] = 26'b11111111111010110000110010;
        x_t[16] = 26'b11111111111110100010100100;
        x_t[17] = 26'b00000000000010000101111011;
        x_t[18] = 26'b00000000000010011111001000;
        x_t[19] = 26'b00000000000011000100100001;
        x_t[20] = 26'b00000000000010110110010010;
        x_t[21] = 26'b11111111100110111100111101;
        x_t[22] = 26'b11111111100111011010010110;
        x_t[23] = 26'b11111111101011000110000011;
        x_t[24] = 26'b11111111100101011110011110;
        x_t[25] = 26'b11111111100110001011100111;
        x_t[26] = 26'b11111111101110000000101011;
        x_t[27] = 26'b11111111101111101001000101;
        x_t[28] = 26'b11111111101100111011110011;
        x_t[29] = 26'b11111111101010011110000101;
        x_t[30] = 26'b11111111101111100001011100;
        x_t[31] = 26'b11111111110001100010101010;
        x_t[32] = 26'b11111111110001111101101000;
        x_t[33] = 26'b11111111110100001111001110;
        x_t[34] = 26'b11111111111000110001000100;
        x_t[35] = 26'b11111111110111001111101100;
        x_t[36] = 26'b11111111110101010110100010;
        x_t[37] = 26'b11111111111001011011100010;
        x_t[38] = 26'b11111111101100000110100110;
        x_t[39] = 26'b11111111110110101101000010;
        x_t[40] = 26'b11111111101000000100011100;
        x_t[41] = 26'b11111111110011000101001111;
        x_t[42] = 26'b11111111011110100011000011;
        x_t[43] = 26'b00000000000001110101101110;
        x_t[44] = 26'b11111111101101101111010011;
        x_t[45] = 26'b11111111110011011001011100;
        x_t[46] = 26'b11111111110011001010110110;
        x_t[47] = 26'b11111111110011111111011001;
        x_t[48] = 26'b11111111111011011010010011;
        x_t[49] = 26'b11111111111011111101101000;
        x_t[50] = 26'b00000000000000001100111001;
        x_t[51] = 26'b00000000000110001011101011;
        x_t[52] = 26'b00000000000011111110111001;
        x_t[53] = 26'b00000000000100011011000111;
        x_t[54] = 26'b00000000000010111011111100;
        x_t[55] = 26'b11111111110110111011011011;
        x_t[56] = 26'b11111111111001101000010000;
        x_t[57] = 26'b00000000000101011101010000;
        x_t[58] = 26'b00000000001000001000110001;
        x_t[59] = 26'b00000000000110010111100001;
        x_t[60] = 26'b11111111111011101000100100;
        x_t[61] = 26'b00000000000010010010011111;
        x_t[62] = 26'b11111111111010101001010111;
        x_t[63] = 26'b11111111111001001001000001;
        
        h_t_prev[0] = 26'b11111111101111111011000110;
        h_t_prev[1] = 26'b11111111111000001101001011;
        h_t_prev[2] = 26'b11111111111010000010000111;
        h_t_prev[3] = 26'b11111111111111001111100000;
        h_t_prev[4] = 26'b00000000000001001100111111;
        h_t_prev[5] = 26'b00000000000001111010101110;
        h_t_prev[6] = 26'b11111111111110101000011101;
        h_t_prev[7] = 26'b11111111111001000010010110;
        h_t_prev[8] = 26'b11111111111110001010110000;
        h_t_prev[9] = 26'b11111111111110110111001100;
        h_t_prev[10] = 26'b00000000000000000010010101;
        h_t_prev[11] = 26'b00000000000010001011010010;
        h_t_prev[12] = 26'b00000000000011110111001001;
        h_t_prev[13] = 26'b00000000000010010000100010;
        h_t_prev[14] = 26'b11111111110011110101101000;
        h_t_prev[15] = 26'b11111111111010110000110010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 70 timeout!");
                $fdisplay(fd_cycles, "Test Vector  70: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  70: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 70");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 71
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111101000100001100011;
        x_t[1] = 26'b11111111110001110010000100;
        x_t[2] = 26'b11111111110011010110110011;
        x_t[3] = 26'b11111111111011010100001000;
        x_t[4] = 26'b11111111111101101110101100;
        x_t[5] = 26'b11111111111101110000011101;
        x_t[6] = 26'b11111111111000110011000011;
        x_t[7] = 26'b11111111101111011111100101;
        x_t[8] = 26'b11111111110111000100111010;
        x_t[9] = 26'b11111111110111010110001000;
        x_t[10] = 26'b11111111111001111010111100;
        x_t[11] = 26'b11111111111111010011110101;
        x_t[12] = 26'b00000000000010011001100000;
        x_t[13] = 26'b11111111111100010010111100;
        x_t[14] = 26'b11111111101111100011011010;
        x_t[15] = 26'b11111111110011110001010001;
        x_t[16] = 26'b11111111111000010110000001;
        x_t[17] = 26'b11111111111110000101010100;
        x_t[18] = 26'b00000000000000110101101101;
        x_t[19] = 26'b00000000000011000100100001;
        x_t[20] = 26'b00000000000000111001001001;
        x_t[21] = 26'b11111111100100111000010110;
        x_t[22] = 26'b11111111100101110100110011;
        x_t[23] = 26'b11111111101010111010011100;
        x_t[24] = 26'b11111111100011111101000010;
        x_t[25] = 26'b11111111100100011011101110;
        x_t[26] = 26'b11111111101011101000100111;
        x_t[27] = 26'b11111111101111101001000101;
        x_t[28] = 26'b11111111101101100001100101;
        x_t[29] = 26'b11111111100111000101110010;
        x_t[30] = 26'b11111111101111000010001110;
        x_t[31] = 26'b11111111110000001001111100;
        x_t[32] = 26'b11111111101110110101101111;
        x_t[33] = 26'b11111111110001101000101101;
        x_t[34] = 26'b11111111110111010001110011;
        x_t[35] = 26'b11111111110110111011111100;
        x_t[36] = 26'b11111111110111001101110100;
        x_t[37] = 26'b11111111111001001011001111;
        x_t[38] = 26'b11111111100101110011001101;
        x_t[39] = 26'b11111111111001011101011010;
        x_t[40] = 26'b11111111100010101000100111;
        x_t[41] = 26'b11111111110011100001000011;
        x_t[42] = 26'b11111111100001001001000100;
        x_t[43] = 26'b11111111111101101110011010;
        x_t[44] = 26'b11111111101110000101101001;
        x_t[45] = 26'b11111111111000101101111010;
        x_t[46] = 26'b11111111110110101110110011;
        x_t[47] = 26'b11111111110110011110100010;
        x_t[48] = 26'b11111111111100000000011010;
        x_t[49] = 26'b11111111111101000111110000;
        x_t[50] = 26'b00000000000011001010111101;
        x_t[51] = 26'b00000000001010101101011101;
        x_t[52] = 26'b00000000001000011101010111;
        x_t[53] = 26'b00000000001001010010111001;
        x_t[54] = 26'b00000000000111011011100110;
        x_t[55] = 26'b11111111111100010100101100;
        x_t[56] = 26'b11111111111110001100011011;
        x_t[57] = 26'b00000000001010110010010011;
        x_t[58] = 26'b00000000001100001110011111;
        x_t[59] = 26'b00000000001010000100010110;
        x_t[60] = 26'b11111111111100000111001110;
        x_t[61] = 26'b00000000000010010010011111;
        x_t[62] = 26'b11111111111011010101110000;
        x_t[63] = 26'b11111111111000010100001101;
        
        h_t_prev[0] = 26'b11111111101000100001100011;
        h_t_prev[1] = 26'b11111111110001110010000100;
        h_t_prev[2] = 26'b11111111110011010110110011;
        h_t_prev[3] = 26'b11111111111011010100001000;
        h_t_prev[4] = 26'b11111111111101101110101100;
        h_t_prev[5] = 26'b11111111111101110000011101;
        h_t_prev[6] = 26'b11111111111000110011000011;
        h_t_prev[7] = 26'b11111111101111011111100101;
        h_t_prev[8] = 26'b11111111110111000100111010;
        h_t_prev[9] = 26'b11111111110111010110001000;
        h_t_prev[10] = 26'b11111111111001111010111100;
        h_t_prev[11] = 26'b11111111111111010011110101;
        h_t_prev[12] = 26'b00000000000010011001100000;
        h_t_prev[13] = 26'b11111111111100010010111100;
        h_t_prev[14] = 26'b11111111101111100011011010;
        h_t_prev[15] = 26'b11111111110011110001010001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 71 timeout!");
                $fdisplay(fd_cycles, "Test Vector  71: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  71: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 71");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 72
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111101010101011101010;
        x_t[1] = 26'b11111111110100110101110101;
        x_t[2] = 26'b11111111110100110111111011;
        x_t[3] = 26'b11111111111101011011011111;
        x_t[4] = 26'b00000000000001110101011001;
        x_t[5] = 26'b00000000000100010110000010;
        x_t[6] = 26'b11111111111101000100111000;
        x_t[7] = 26'b11111111110101100010011001;
        x_t[8] = 26'b11111111111001000000101100;
        x_t[9] = 26'b11111111111001110110011111;
        x_t[10] = 26'b11111111111101111001010110;
        x_t[11] = 26'b00000000000101010111001000;
        x_t[12] = 26'b00000000001001101101110000;
        x_t[13] = 26'b00000000000100011000110101;
        x_t[14] = 26'b11111111110011110101101000;
        x_t[15] = 26'b11111111110101010110111110;
        x_t[16] = 26'b11111111111010100000110011;
        x_t[17] = 26'b00000000000001110010001100;
        x_t[18] = 26'b00000000001000011010101000;
        x_t[19] = 26'b00000000001010010001110101;
        x_t[20] = 26'b00000000001001011111110000;
        x_t[21] = 26'b11111111101000101011011110;
        x_t[22] = 26'b11111111101001110010101001;
        x_t[23] = 26'b11111111101101000101101010;
        x_t[24] = 26'b11111111100111001100000101;
        x_t[25] = 26'b11111111100111010110001100;
        x_t[26] = 26'b11111111110000000111110110;
        x_t[27] = 26'b11111111110011010100111010;
        x_t[28] = 26'b11111111101111101100001000;
        x_t[29] = 26'b11111111101001111100110011;
        x_t[30] = 26'b11111111110100111000111000;
        x_t[31] = 26'b11111111110101101100110011;
        x_t[32] = 26'b11111111110001111101101000;
        x_t[33] = 26'b11111111110101000110101111;
        x_t[34] = 26'b11111111111011011100100010;
        x_t[35] = 26'b11111111111011010000010001;
        x_t[36] = 26'b11111111111011100100001000;
        x_t[37] = 26'b11111111111000111010111011;
        x_t[38] = 26'b11111111101110010011110010;
        x_t[39] = 26'b11111111111101100101111111;
        x_t[40] = 26'b11111111110011111101010011;
        x_t[41] = 26'b11111111111010011110001001;
        x_t[42] = 26'b11111111100011101111000101;
        x_t[43] = 26'b00000000000010100001100111;
        x_t[44] = 26'b11111111110010101000000111;
        x_t[45] = 26'b00000000000000011101001001;
        x_t[46] = 26'b11111111111010111100001100;
        x_t[47] = 26'b11111111111001100101011101;
        x_t[48] = 26'b11111111111101001100101001;
        x_t[49] = 26'b00000000000000111000101100;
        x_t[50] = 26'b00000000000111000010000001;
        x_t[51] = 26'b00000000001110111011111010;
        x_t[52] = 26'b00000000001011111110011101;
        x_t[53] = 26'b00000000001101000111110110;
        x_t[54] = 26'b00000000001010110011010110;
        x_t[55] = 26'b00000000000000101000111010;
        x_t[56] = 26'b00000000000001011010101010;
        x_t[57] = 26'b00000000001101011100110101;
        x_t[58] = 26'b00000000001110111100111101;
        x_t[59] = 26'b00000000001100100010001111;
        x_t[60] = 26'b00000000000001001001010000;
        x_t[61] = 26'b00000000001000011111110001;
        x_t[62] = 26'b00000000000001000111100111;
        x_t[63] = 26'b11111111111110111010101011;
        
        h_t_prev[0] = 26'b11111111101010101011101010;
        h_t_prev[1] = 26'b11111111110100110101110101;
        h_t_prev[2] = 26'b11111111110100110111111011;
        h_t_prev[3] = 26'b11111111111101011011011111;
        h_t_prev[4] = 26'b00000000000001110101011001;
        h_t_prev[5] = 26'b00000000000100010110000010;
        h_t_prev[6] = 26'b11111111111101000100111000;
        h_t_prev[7] = 26'b11111111110101100010011001;
        h_t_prev[8] = 26'b11111111111001000000101100;
        h_t_prev[9] = 26'b11111111111001110110011111;
        h_t_prev[10] = 26'b11111111111101111001010110;
        h_t_prev[11] = 26'b00000000000101010111001000;
        h_t_prev[12] = 26'b00000000001001101101110000;
        h_t_prev[13] = 26'b00000000000100011000110101;
        h_t_prev[14] = 26'b11111111110011110101101000;
        h_t_prev[15] = 26'b11111111110101010110111110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 72 timeout!");
                $fdisplay(fd_cycles, "Test Vector  72: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  72: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 72");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 73
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111110001110001011110;
        x_t[1] = 26'b11111111111000110100010101;
        x_t[2] = 26'b11111111111000001101100101;
        x_t[3] = 26'b00000000000000001001100001;
        x_t[4] = 26'b00000000000011000110001110;
        x_t[5] = 26'b00000000000011101001101010;
        x_t[6] = 26'b11111111111101110110101011;
        x_t[7] = 26'b11111111110110110011110101;
        x_t[8] = 26'b11111111111001000000101100;
        x_t[9] = 26'b11111111111011011010101101;
        x_t[10] = 26'b11111111111111011011001100;
        x_t[11] = 26'b00000000000100011001111110;
        x_t[12] = 26'b00000000000110110010011101;
        x_t[13] = 26'b00000000000000100011100001;
        x_t[14] = 26'b11111111110000100010101100;
        x_t[15] = 26'b11111111110101000010101001;
        x_t[16] = 26'b11111111111011110000000111;
        x_t[17] = 26'b00000000000010011001101011;
        x_t[18] = 26'b00000000000110011100001000;
        x_t[19] = 26'b00000000000110110110001010;
        x_t[20] = 26'b00000000000101001100011101;
        x_t[21] = 26'b11111111101011111101011100;
        x_t[22] = 26'b11111111101100100100010110;
        x_t[23] = 26'b11111111101110101110000101;
        x_t[24] = 26'b11111111101010011011001000;
        x_t[25] = 26'b11111111101010110101111110;
        x_t[26] = 26'b11111111110011000001101110;
        x_t[27] = 26'b11111111110011100100101000;
        x_t[28] = 26'b11111111101110101101001010;
        x_t[29] = 26'b11111111101101010101000110;
        x_t[30] = 26'b11111111111001010001110111;
        x_t[31] = 26'b11111111110101011011000011;
        x_t[32] = 26'b11111111110101010111101101;
        x_t[33] = 26'b11111111110110110101110000;
        x_t[34] = 26'b11111111111011101111100101;
        x_t[35] = 26'b11111111111100001011011111;
        x_t[36] = 26'b11111111111000011101010101;
        x_t[37] = 26'b11111111111000111010111011;
        x_t[38] = 26'b11111111110010101110001010;
        x_t[39] = 26'b11111111111001011101011010;
        x_t[40] = 26'b11111111101111001100111101;
        x_t[41] = 26'b00000000000101010101100110;
        x_t[42] = 26'b11111111100010111111101001;
        x_t[43] = 26'b11111111110110110111100011;
        x_t[44] = 26'b11111111110011101011001000;
        x_t[45] = 26'b11111111110100010111010110;
        x_t[46] = 26'b11111111111100001111000101;
        x_t[47] = 26'b11111111111000101001110010;
        x_t[48] = 26'b11111111111100111001100110;
        x_t[49] = 26'b11111111111110100100011011;
        x_t[50] = 26'b00000000000011011101111101;
        x_t[51] = 26'b00000000000110001011101011;
        x_t[52] = 26'b00000000000010101101000010;
        x_t[53] = 26'b00000000000010010101100000;
        x_t[54] = 26'b11111111111110000100010011;
        x_t[55] = 26'b11111111111110011110110011;
        x_t[56] = 26'b11111111111110111111111111;
        x_t[57] = 26'b00000000000110110010100001;
        x_t[58] = 26'b00000000000100100101111101;
        x_t[59] = 26'b00000000000000111100001010;
        x_t[60] = 26'b00000000000011010011010001;
        x_t[61] = 26'b00000000000111111110101010;
        x_t[62] = 26'b11111111111111101110110110;
        x_t[63] = 26'b11111111111101100010101010;
        
        h_t_prev[0] = 26'b11111111110001110001011110;
        h_t_prev[1] = 26'b11111111111000110100010101;
        h_t_prev[2] = 26'b11111111111000001101100101;
        h_t_prev[3] = 26'b00000000000000001001100001;
        h_t_prev[4] = 26'b00000000000011000110001110;
        h_t_prev[5] = 26'b00000000000011101001101010;
        h_t_prev[6] = 26'b11111111111101110110101011;
        h_t_prev[7] = 26'b11111111110110110011110101;
        h_t_prev[8] = 26'b11111111111001000000101100;
        h_t_prev[9] = 26'b11111111111011011010101101;
        h_t_prev[10] = 26'b11111111111111011011001100;
        h_t_prev[11] = 26'b00000000000100011001111110;
        h_t_prev[12] = 26'b00000000000110110010011101;
        h_t_prev[13] = 26'b00000000000000100011100001;
        h_t_prev[14] = 26'b11111111110000100010101100;
        h_t_prev[15] = 26'b11111111110101000010101001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 73 timeout!");
                $fdisplay(fd_cycles, "Test Vector  73: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  73: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 73");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 74
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111110011010100001000;
        x_t[1] = 26'b11111111111011111000000111;
        x_t[2] = 26'b11111111111001101110101100;
        x_t[3] = 26'b00000000000001000011100001;
        x_t[4] = 26'b00000000000001001100111111;
        x_t[5] = 26'b00000000000000100001111101;
        x_t[6] = 26'b11111111111011111010001101;
        x_t[7] = 26'b11111111111001101011000100;
        x_t[8] = 26'b11111111111011100101101110;
        x_t[9] = 26'b11111111111101111011000100;
        x_t[10] = 26'b00000000000000111101000011;
        x_t[11] = 26'b00000000000100011001111110;
        x_t[12] = 26'b00000000000100100101111110;
        x_t[13] = 26'b11111111111111010001101111;
        x_t[14] = 26'b11111111110101110100001100;
        x_t[15] = 26'b11111111111010001000000110;
        x_t[16] = 26'b11111111111110110110011001;
        x_t[17] = 26'b00000000000100010000000111;
        x_t[18] = 26'b00000000000011001001010011;
        x_t[19] = 26'b00000000000011000100100001;
        x_t[20] = 26'b00000000000010011101010000;
        x_t[21] = 26'b11111111101101001010110011;
        x_t[22] = 26'b11111111101101001010011011;
        x_t[23] = 26'b11111111110000001010111001;
        x_t[24] = 26'b11111111101011110000011000;
        x_t[25] = 26'b11111111101100001100111111;
        x_t[26] = 26'b11111111110101001000111001;
        x_t[27] = 26'b11111111110101000010111101;
        x_t[28] = 26'b11111111110001000100010011;
        x_t[29] = 26'b11111111101100110011110100;
        x_t[30] = 26'b11111111111001110001000101;
        x_t[31] = 26'b11111111110111010111010000;
        x_t[32] = 26'b11111111110111010110111010;
        x_t[33] = 26'b11111111111000110111010001;
        x_t[34] = 26'b11111111111101001110110110;
        x_t[35] = 26'b11111111111101000110101101;
        x_t[36] = 26'b11111111111010000000101110;
        x_t[37] = 26'b11111111111101110000110001;
        x_t[38] = 26'b11111111101101010111010001;
        x_t[39] = 26'b11111111111101100101111111;
        x_t[40] = 26'b11111111101100011111000011;
        x_t[41] = 26'b00000000001011110110110111;
        x_t[42] = 26'b11111111100111011100010000;
        x_t[43] = 26'b11111111110011011100001000;
        x_t[44] = 26'b11111111110110000111100010;
        x_t[45] = 26'b11111111111001001100110111;
        x_t[46] = 26'b11111111111110110100110111;
        x_t[47] = 26'b11111111111111011111011011;
        x_t[48] = 26'b00000000000100101001000111;
        x_t[49] = 26'b00000000000100000100100100;
        x_t[50] = 26'b00000000000110001001000000;
        x_t[51] = 26'b00000000000110011110111111;
        x_t[52] = 26'b00000000000011010101111101;
        x_t[53] = 26'b00000000000011101110100101;
        x_t[54] = 26'b00000000000010100011111110;
        x_t[55] = 26'b00000000000110010011011100;
        x_t[56] = 26'b00000000000101011100011101;
        x_t[57] = 26'b00000000001010010000001100;
        x_t[58] = 26'b00000000000100010100100000;
        x_t[59] = 26'b00000000000010101010101011;
        x_t[60] = 26'b00000000000101111011111101;
        x_t[61] = 26'b00000000000101111010001111;
        x_t[62] = 26'b11111111111100010000111011;
        x_t[63] = 26'b11111111111100111111011101;
        
        h_t_prev[0] = 26'b11111111110011010100001000;
        h_t_prev[1] = 26'b11111111111011111000000111;
        h_t_prev[2] = 26'b11111111111001101110101100;
        h_t_prev[3] = 26'b00000000000001000011100001;
        h_t_prev[4] = 26'b00000000000001001100111111;
        h_t_prev[5] = 26'b00000000000000100001111101;
        h_t_prev[6] = 26'b11111111111011111010001101;
        h_t_prev[7] = 26'b11111111111001101011000100;
        h_t_prev[8] = 26'b11111111111011100101101110;
        h_t_prev[9] = 26'b11111111111101111011000100;
        h_t_prev[10] = 26'b00000000000000111101000011;
        h_t_prev[11] = 26'b00000000000100011001111110;
        h_t_prev[12] = 26'b00000000000100100101111110;
        h_t_prev[13] = 26'b11111111111111010001101111;
        h_t_prev[14] = 26'b11111111110101110100001100;
        h_t_prev[15] = 26'b11111111111010001000000110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 74 timeout!");
                $fdisplay(fd_cycles, "Test Vector  74: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  74: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 74");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 75
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111110010000101001101;
        x_t[1] = 26'b11111111111101000110011011;
        x_t[2] = 26'b11111111111010000010000111;
        x_t[3] = 26'b00000000000000110000001100;
        x_t[4] = 26'b00000000000000100100100100;
        x_t[5] = 26'b00000000000001111010101110;
        x_t[6] = 26'b11111111111101000100111000;
        x_t[7] = 26'b11111111111101110011101110;
        x_t[8] = 26'b00000000000000000110100010;
        x_t[9] = 26'b11111111111111001011001111;
        x_t[10] = 26'b11111111111111011011001100;
        x_t[11] = 26'b00000000000100011001111110;
        x_t[12] = 26'b00000000000011001000010101;
        x_t[13] = 26'b00000000000000100011100001;
        x_t[14] = 26'b11111111111011101111111000;
        x_t[15] = 26'b11111111111110010000100010;
        x_t[16] = 26'b00000000000000000101101100;
        x_t[17] = 26'b00000000000010000101111011;
        x_t[18] = 26'b11111111111111110110011101;
        x_t[19] = 26'b11111111111111010010111001;
        x_t[20] = 26'b00000000000000111001001001;
        x_t[21] = 26'b11111111101101101011111101;
        x_t[22] = 26'b11111111101110100011010001;
        x_t[23] = 26'b11111111110000111001010011;
        x_t[24] = 26'b11111111101010100111010011;
        x_t[25] = 26'b11111111101011000010011001;
        x_t[26] = 26'b11111111110100111000000000;
        x_t[27] = 26'b11111111110101100010011010;
        x_t[28] = 26'b11111111110010011100011101;
        x_t[29] = 26'b11111111101010111111010111;
        x_t[30] = 26'b11111111110101110111010100;
        x_t[31] = 26'b11111111110100110111100100;
        x_t[32] = 26'b11111111110100100001001100;
        x_t[33] = 26'b11111111110101111110001111;
        x_t[34] = 26'b11111111111010010000010101;
        x_t[35] = 26'b11111111111001011001110110;
        x_t[36] = 26'b11111111111000011101010101;
        x_t[37] = 26'b11111111111010011100110001;
        x_t[38] = 26'b11111111101111100100011101;
        x_t[39] = 26'b11111111110111100111110101;
        x_t[40] = 26'b11111111110011100111100100;
        x_t[41] = 26'b11111111110110000111111110;
        x_t[42] = 26'b11111111101011100001001000;
        x_t[43] = 26'b11111111101101010001001010;
        x_t[44] = 26'b11111111110110110100001110;
        x_t[45] = 26'b11111111110001111100100101;
        x_t[46] = 26'b11111111111110110100110111;
        x_t[47] = 26'b11111111111110001111110111;
        x_t[48] = 26'b00000000000001101010100010;
        x_t[49] = 26'b11111111111110100100011011;
        x_t[50] = 26'b11111111111100111011110110;
        x_t[51] = 26'b11111111111100110100110011;
        x_t[52] = 26'b11111111111000011110001111;
        x_t[53] = 26'b11111111111011101110011000;
        x_t[54] = 26'b11111111111011000100100010;
        x_t[55] = 26'b00000000000011010101100011;
        x_t[56] = 26'b00000000000001101011110110;
        x_t[57] = 26'b00000000000010010000101000;
        x_t[58] = 26'b11111111111011100110001100;
        x_t[59] = 26'b11111111111110001110011110;
        x_t[60] = 26'b00000000000110101001111101;
        x_t[61] = 26'b00000000000011100101010000;
        x_t[62] = 26'b11111111111010011010100100;
        x_t[63] = 26'b11111111111110010111011110;
        
        h_t_prev[0] = 26'b11111111110010000101001101;
        h_t_prev[1] = 26'b11111111111101000110011011;
        h_t_prev[2] = 26'b11111111111010000010000111;
        h_t_prev[3] = 26'b00000000000000110000001100;
        h_t_prev[4] = 26'b00000000000000100100100100;
        h_t_prev[5] = 26'b00000000000001111010101110;
        h_t_prev[6] = 26'b11111111111101000100111000;
        h_t_prev[7] = 26'b11111111111101110011101110;
        h_t_prev[8] = 26'b00000000000000000110100010;
        h_t_prev[9] = 26'b11111111111111001011001111;
        h_t_prev[10] = 26'b11111111111111011011001100;
        h_t_prev[11] = 26'b00000000000100011001111110;
        h_t_prev[12] = 26'b00000000000011001000010101;
        h_t_prev[13] = 26'b00000000000000100011100001;
        h_t_prev[14] = 26'b11111111111011101111111000;
        h_t_prev[15] = 26'b11111111111110010000100010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 75 timeout!");
                $fdisplay(fd_cycles, "Test Vector  75: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  75: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 75");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 76
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111101110101100001010;
        x_t[1] = 26'b11111111110011111011000110;
        x_t[2] = 26'b11111111110011010110110011;
        x_t[3] = 26'b11111111111011100111011110;
        x_t[4] = 26'b11111111111010111000110100;
        x_t[5] = 26'b11111111111001010000000000;
        x_t[6] = 26'b11111111110101010011000000;
        x_t[7] = 26'b11111111110110001011000111;
        x_t[8] = 26'b11111111111000010111011011;
        x_t[9] = 26'b11111111110111000010000101;
        x_t[10] = 26'b11111111110111011110011000;
        x_t[11] = 26'b11111111111101000101001010;
        x_t[12] = 26'b11111111111001100111100110;
        x_t[13] = 26'b11111111110100101000010100;
        x_t[14] = 26'b11111111110111001000100100;
        x_t[15] = 26'b11111111110111111001101101;
        x_t[16] = 26'b11111111111000101001110110;
        x_t[17] = 26'b11111111111000100001111111;
        x_t[18] = 26'b11111111110110010011000001;
        x_t[19] = 26'b11111111110111000011101011;
        x_t[20] = 26'b11111111110111111001100000;
        x_t[21] = 26'b11111111101101010101110110;
        x_t[22] = 26'b11111111101110001001111001;
        x_t[23] = 26'b11111111110000101101101100;
        x_t[24] = 26'b11111111101010110011011111;
        x_t[25] = 26'b11111111101011000010011001;
        x_t[26] = 26'b11111111110100111000000000;
        x_t[27] = 26'b11111111110011110100010110;
        x_t[28] = 26'b11111111110001000100010011;
        x_t[29] = 26'b11111111101100100011001100;
        x_t[30] = 26'b11111111110110000110111011;
        x_t[31] = 26'b11111111110010111011011000;
        x_t[32] = 26'b11111111110101000101100010;
        x_t[33] = 26'b11111111110111011010110000;
        x_t[34] = 26'b11111111111010110110011011;
        x_t[35] = 26'b11111111111001011001110110;
        x_t[36] = 26'b11111111110101111110010011;
        x_t[37] = 26'b11111111111000011010010100;
        x_t[38] = 26'b11111111110110100000001100;
        x_t[39] = 26'b11111111110100110111011100;
        x_t[40] = 26'b11111111111010000100100110;
        x_t[41] = 26'b11111111110000111010001001;
        x_t[42] = 26'b11111111110100110010000010;
        x_t[43] = 26'b11111111110011011100001000;
        x_t[44] = 26'b11111111110111110111010000;
        x_t[45] = 26'b11111111110101110100001100;
        x_t[46] = 26'b00000000000000011100011110;
        x_t[47] = 26'b11111111111111001011100010;
        x_t[48] = 26'b00000000000001000100011010;
        x_t[49] = 26'b11111111111100110101001110;
        x_t[50] = 26'b11111111111010110110110011;
        x_t[51] = 26'b11111111111011000000111001;
        x_t[52] = 26'b11111111111000110010101101;
        x_t[53] = 26'b11111111111110100000100010;
        x_t[54] = 26'b11111111111111111100001010;
        x_t[55] = 26'b00000000000101110000111010;
        x_t[56] = 26'b00000000000011110101010110;
        x_t[57] = 26'b00000000000001111111100101;
        x_t[58] = 26'b11111111111101001110111000;
        x_t[59] = 26'b00000000000010111010011110;
        x_t[60] = 26'b00000000000101111011111101;
        x_t[61] = 26'b00000000000011000100001001;
        x_t[62] = 26'b11111111111011100100100010;
        x_t[63] = 26'b00000000000011100101111011;
        
        h_t_prev[0] = 26'b11111111101110101100001010;
        h_t_prev[1] = 26'b11111111110011111011000110;
        h_t_prev[2] = 26'b11111111110011010110110011;
        h_t_prev[3] = 26'b11111111111011100111011110;
        h_t_prev[4] = 26'b11111111111010111000110100;
        h_t_prev[5] = 26'b11111111111001010000000000;
        h_t_prev[6] = 26'b11111111110101010011000000;
        h_t_prev[7] = 26'b11111111110110001011000111;
        h_t_prev[8] = 26'b11111111111000010111011011;
        h_t_prev[9] = 26'b11111111110111000010000101;
        h_t_prev[10] = 26'b11111111110111011110011000;
        h_t_prev[11] = 26'b11111111111101000101001010;
        h_t_prev[12] = 26'b11111111111001100111100110;
        h_t_prev[13] = 26'b11111111110100101000010100;
        h_t_prev[14] = 26'b11111111110111001000100100;
        h_t_prev[15] = 26'b11111111110111111001101101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 76 timeout!");
                $fdisplay(fd_cycles, "Test Vector  76: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  76: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 76");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 77
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111111000100011100011;
        x_t[1] = 26'b11111111111101011010000000;
        x_t[2] = 26'b11111111111100001010000101;
        x_t[3] = 26'b00000000000011011110001101;
        x_t[4] = 26'b00000000000011000110001110;
        x_t[5] = 26'b00000000000000100001111101;
        x_t[6] = 26'b11111111111010101111100001;
        x_t[7] = 26'b00000000000101011100010101;
        x_t[8] = 26'b00000000000011000000001100;
        x_t[9] = 26'b00000000000000000111011000;
        x_t[10] = 26'b00000000000000101001011110;
        x_t[11] = 26'b00000000000110101000101010;
        x_t[12] = 26'b00000000000010000010000101;
        x_t[13] = 26'b11111111111100101110001101;
        x_t[14] = 26'b00000000000001010110011110;
        x_t[15] = 26'b00000000000010011000111111;
        x_t[16] = 26'b00000000000001000001001011;
        x_t[17] = 26'b00000000000001001010101101;
        x_t[18] = 26'b11111111111110001101000010;
        x_t[19] = 26'b11111111111111010010111001;
        x_t[20] = 26'b00000000000010000100001110;
        x_t[21] = 26'b11111111110001101010001000;
        x_t[22] = 26'b11111111110010010100011100;
        x_t[23] = 26'b11111111110011100111010100;
        x_t[24] = 26'b11111111110001000101011010;
        x_t[25] = 26'b11111111110001000011110010;
        x_t[26] = 26'b11111111111010101011101110;
        x_t[27] = 26'b11111111111000111110100000;
        x_t[28] = 26'b11111111110011011011011100;
        x_t[29] = 26'b11111111110100010110010101;
        x_t[30] = 26'b00000000000000000110111101;
        x_t[31] = 26'b11111111111010111101111010;
        x_t[32] = 26'b11111111111011100111011111;
        x_t[33] = 26'b11111111111100111010010011;
        x_t[34] = 26'b00000000000001011001100101;
        x_t[35] = 26'b11111111111111100100100110;
        x_t[36] = 26'b11111111111011100100001000;
        x_t[37] = 26'b11111111111100101111100010;
        x_t[38] = 26'b11111111111110000100010001;
        x_t[39] = 26'b11111111110110101101000010;
        x_t[40] = 26'b00000000000000110111011000;
        x_t[41] = 26'b11111111110111110111001111;
        x_t[42] = 26'b11111111110100000010100110;
        x_t[43] = 26'b11111111111110011010010011;
        x_t[44] = 26'b11111111111111111001001010;
        x_t[45] = 26'b11111111111001001100110111;
        x_t[46] = 26'b00000000000101010011010011;
        x_t[47] = 26'b00000000000011110101111011;
        x_t[48] = 26'b00000000000101110101010110;
        x_t[49] = 26'b00000000000000010011101000;
        x_t[50] = 26'b11111111111101001110110110;
        x_t[51] = 26'b11111111111011111010110110;
        x_t[52] = 26'b11111111111001000111001010;
        x_t[53] = 26'b11111111111101011101101110;
        x_t[54] = 26'b11111111111110011100010010;
        x_t[55] = 26'b00000000000111000111001111;
        x_t[56] = 26'b00000000000100111010000110;
        x_t[57] = 26'b00000000000000111011010111;
        x_t[58] = 26'b11111111111011000011010010;
        x_t[59] = 26'b11111111111101001111010100;
        x_t[60] = 26'b00000000000110111001010010;
        x_t[61] = 26'b00000000000101001000100100;
        x_t[62] = 26'b11111111111011010101110000;
        x_t[63] = 26'b00000000001000110100011000;
        
        h_t_prev[0] = 26'b11111111111000100011100011;
        h_t_prev[1] = 26'b11111111111101011010000000;
        h_t_prev[2] = 26'b11111111111100001010000101;
        h_t_prev[3] = 26'b00000000000011011110001101;
        h_t_prev[4] = 26'b00000000000011000110001110;
        h_t_prev[5] = 26'b00000000000000100001111101;
        h_t_prev[6] = 26'b11111111111010101111100001;
        h_t_prev[7] = 26'b00000000000101011100010101;
        h_t_prev[8] = 26'b00000000000011000000001100;
        h_t_prev[9] = 26'b00000000000000000111011000;
        h_t_prev[10] = 26'b00000000000000101001011110;
        h_t_prev[11] = 26'b00000000000110101000101010;
        h_t_prev[12] = 26'b00000000000010000010000101;
        h_t_prev[13] = 26'b11111111111100101110001101;
        h_t_prev[14] = 26'b00000000000001010110011110;
        h_t_prev[15] = 26'b00000000000010011000111111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 77 timeout!");
                $fdisplay(fd_cycles, "Test Vector  77: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  77: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 77");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 78
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111111010011001111100;
        x_t[1] = 26'b11111111111101011010000000;
        x_t[2] = 26'b11111111111010000010000111;
        x_t[3] = 26'b11111111111111100010110110;
        x_t[4] = 26'b11111111111110010111000111;
        x_t[5] = 26'b11111111111100101101111001;
        x_t[6] = 26'b11111111110111001111011110;
        x_t[7] = 26'b00000000000001111100011001;
        x_t[8] = 26'b11111111111111011101010001;
        x_t[9] = 26'b11111111111100010110110110;
        x_t[10] = 26'b11111111111011011100110010;
        x_t[11] = 26'b11111111111110101011000100;
        x_t[12] = 26'b11111111111000100001010111;
        x_t[13] = 26'b11111111110100101000010100;
        x_t[14] = 26'b11111111111010000110011010;
        x_t[15] = 26'b11111111111100000010001001;
        x_t[16] = 26'b11111111111010100000110011;
        x_t[17] = 26'b11111111111010011000011011;
        x_t[18] = 26'b11111111110101010011110001;
        x_t[19] = 26'b11111111110100101001111010;
        x_t[20] = 26'b11111111110101001010010100;
        x_t[21] = 26'b11111111101110111001010100;
        x_t[22] = 26'b11111111101111101111011011;
        x_t[23] = 26'b11111111110000001010111001;
        x_t[24] = 26'b11111111101101011110000000;
        x_t[25] = 26'b11111111101101110000011100;
        x_t[26] = 26'b11111111110100111000000000;
        x_t[27] = 26'b11111111110100010011110011;
        x_t[28] = 26'b11111111110000000101010100;
        x_t[29] = 26'b11111111101100100011001100;
        x_t[30] = 26'b11111111111110011001101100;
        x_t[31] = 26'b11111111110100000010010110;
        x_t[32] = 26'b11111111110100001111000001;
        x_t[33] = 26'b11111111110100100001101111;
        x_t[34] = 26'b11111111111001010111001011;
        x_t[35] = 26'b11111111111000001010111001;
        x_t[36] = 26'b11111111110100011010111001;
        x_t[37] = 26'b11111111110101010110100111;
        x_t[38] = 26'b11111111110001110001101001;
        x_t[39] = 26'b11111111101110111001010011;
        x_t[40] = 26'b11111111110001111010110111;
        x_t[41] = 26'b11111111110110000111111110;
        x_t[42] = 26'b11111111100101100101101010;
        x_t[43] = 26'b11111111101110101000111011;
        x_t[44] = 26'b11111111110100101110001010;
        x_t[45] = 26'b11111111100101110110110010;
        x_t[46] = 26'b11111111111000111111110111;
        x_t[47] = 26'b11111111110110110010011011;
        x_t[48] = 26'b11111111111000001000101001;
        x_t[49] = 26'b11111111110011100100001010;
        x_t[50] = 26'b11111111110001010110101000;
        x_t[51] = 26'b11111111110000001001011011;
        x_t[52] = 26'b11111111101100101001001000;
        x_t[53] = 26'b11111111101111100010111101;
        x_t[54] = 26'b11111111101101111101100001;
        x_t[55] = 26'b11111111111100100101111101;
        x_t[56] = 26'b11111111111010111110001011;
        x_t[57] = 26'b11111111110110110011011000;
        x_t[58] = 26'b11111111110001100000101000;
        x_t[59] = 26'b11111111110010011000100110;
        x_t[60] = 26'b00000000000011010011010001;
        x_t[61] = 26'b11111111111111101100111100;
        x_t[62] = 26'b11111111110011000001001000;
        x_t[63] = 26'b00000000000011000010101110;
        
        h_t_prev[0] = 26'b11111111111010011001111100;
        h_t_prev[1] = 26'b11111111111101011010000000;
        h_t_prev[2] = 26'b11111111111010000010000111;
        h_t_prev[3] = 26'b11111111111111100010110110;
        h_t_prev[4] = 26'b11111111111110010111000111;
        h_t_prev[5] = 26'b11111111111100101101111001;
        h_t_prev[6] = 26'b11111111110111001111011110;
        h_t_prev[7] = 26'b00000000000001111100011001;
        h_t_prev[8] = 26'b11111111111111011101010001;
        h_t_prev[9] = 26'b11111111111100010110110110;
        h_t_prev[10] = 26'b11111111111011011100110010;
        h_t_prev[11] = 26'b11111111111110101011000100;
        h_t_prev[12] = 26'b11111111111000100001010111;
        h_t_prev[13] = 26'b11111111110100101000010100;
        h_t_prev[14] = 26'b11111111111010000110011010;
        h_t_prev[15] = 26'b11111111111100000010001001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 78 timeout!");
                $fdisplay(fd_cycles, "Test Vector  78: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  78: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 78");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 79
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111110100100011000011;
        x_t[1] = 26'b11111111111001000111111010;
        x_t[2] = 26'b11111111110110011001000010;
        x_t[3] = 26'b11111111111010000110110010;
        x_t[4] = 26'b11111111111010100100100111;
        x_t[5] = 26'b11111111111001100110001100;
        x_t[6] = 26'b11111111110111001111011110;
        x_t[7] = 26'b11111111110111110000111010;
        x_t[8] = 26'b11111111111000010111011011;
        x_t[9] = 26'b11111111110111101010001011;
        x_t[10] = 26'b11111111110110100011101011;
        x_t[11] = 26'b11111111111011011111001111;
        x_t[12] = 26'b11111111110101111101011110;
        x_t[13] = 26'b11111111110100101000010100;
        x_t[14] = 26'b11111111110011100000100010;
        x_t[15] = 26'b11111111110100101110010011;
        x_t[16] = 26'b11111111110100111011111010;
        x_t[17] = 26'b11111111110101011100100110;
        x_t[18] = 26'b11111111110011010101010001;
        x_t[19] = 26'b11111111110011101000000000;
        x_t[20] = 26'b11111111110100011000010000;
        x_t[21] = 26'b11111111101111100101100001;
        x_t[22] = 26'b11111111101111111100001000;
        x_t[23] = 26'b11111111110000010110011111;
        x_t[24] = 26'b11111111101110110011010000;
        x_t[25] = 26'b11111111101110100010001011;
        x_t[26] = 26'b11111111110111010000000100;
        x_t[27] = 26'b11111111110101110010001000;
        x_t[28] = 26'b11111111110000000101010100;
        x_t[29] = 26'b11111111101111111011011110;
        x_t[30] = 26'b11111111111100111100000001;
        x_t[31] = 26'b11111111110101101100110011;
        x_t[32] = 26'b11111111110111111011010000;
        x_t[33] = 26'b11111111111001001001110001;
        x_t[34] = 26'b11111111111100010101101100;
        x_t[35] = 26'b11111111111010111100100010;
        x_t[36] = 26'b11111111110111100001101100;
        x_t[37] = 26'b11111111111000011010010100;
        x_t[38] = 26'b11111111110101100011101100;
        x_t[39] = 26'b11111111111001111010110100;
        x_t[40] = 26'b11111111111001101110110111;
        x_t[41] = 26'b00000000000101110001011010;
        x_t[42] = 26'b11111111101000111011000111;
        x_t[43] = 26'b11111111100111110010000100;
        x_t[44] = 26'b11111111110101011010110110;
        x_t[45] = 26'b11111111101100101000000111;
        x_t[46] = 26'b11111111111010100111011110;
        x_t[47] = 26'b11111111110111000110010100;
        x_t[48] = 26'b11111111111000011011101101;
        x_t[49] = 26'b11111111110101111000011011;
        x_t[50] = 26'b11111111110101100000101101;
        x_t[51] = 26'b11111111110111111111101101;
        x_t[52] = 26'b11111111110100101000101100;
        x_t[53] = 26'b11111111110111001100111000;
        x_t[54] = 26'b11111111110101011100111101;
        x_t[55] = 26'b11111111111110001101100010;
        x_t[56] = 26'b11111111111100100101010011;
        x_t[57] = 26'b11111111111100101010100010;
        x_t[58] = 26'b11111111111010110001110110;
        x_t[59] = 26'b11111111111010110001011011;
        x_t[60] = 26'b11111111111111011101111010;
        x_t[61] = 26'b11111111111011010011100010;
        x_t[62] = 26'b11111111101111100011001101;
        x_t[63] = 26'b11111111111101100010101010;
        
        h_t_prev[0] = 26'b11111111110100100011000011;
        h_t_prev[1] = 26'b11111111111001000111111010;
        h_t_prev[2] = 26'b11111111110110011001000010;
        h_t_prev[3] = 26'b11111111111010000110110010;
        h_t_prev[4] = 26'b11111111111010100100100111;
        h_t_prev[5] = 26'b11111111111001100110001100;
        h_t_prev[6] = 26'b11111111110111001111011110;
        h_t_prev[7] = 26'b11111111110111110000111010;
        h_t_prev[8] = 26'b11111111111000010111011011;
        h_t_prev[9] = 26'b11111111110111101010001011;
        h_t_prev[10] = 26'b11111111110110100011101011;
        h_t_prev[11] = 26'b11111111111011011111001111;
        h_t_prev[12] = 26'b11111111110101111101011110;
        h_t_prev[13] = 26'b11111111110100101000010100;
        h_t_prev[14] = 26'b11111111110011100000100010;
        h_t_prev[15] = 26'b11111111110100101110010011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 79 timeout!");
                $fdisplay(fd_cycles, "Test Vector  79: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  79: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 79");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 80
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111110101011110010000;
        x_t[1] = 26'b11111111111010111101011000;
        x_t[2] = 26'b11111111111010000010000111;
        x_t[3] = 26'b11111111111110101000110101;
        x_t[4] = 26'b11111111111111010011101111;
        x_t[5] = 26'b00000000000000001011110001;
        x_t[6] = 26'b11111111111010101111100001;
        x_t[7] = 26'b11111111111011111001100100;
        x_t[8] = 26'b11111111111010010011001101;
        x_t[9] = 26'b11111111111010001010100010;
        x_t[10] = 26'b11111111111010100010000101;
        x_t[11] = 26'b00000000000000100101011000;
        x_t[12] = 26'b11111111111101010001101110;
        x_t[13] = 26'b11111111111011110111101100;
        x_t[14] = 26'b11111111110101011111000110;
        x_t[15] = 26'b11111111110110010100000000;
        x_t[16] = 26'b11111111111000111101101011;
        x_t[17] = 26'b11111111111000110101101111;
        x_t[18] = 26'b11111111111010010000000010;
        x_t[19] = 26'b11111111111011110111001110;
        x_t[20] = 26'b11111111111100001100110100;
        x_t[21] = 26'b11111111110000000110101011;
        x_t[22] = 26'b11111111101111001001010110;
        x_t[23] = 26'b11111111110000001010111001;
        x_t[24] = 26'b11111111101110111111011011;
        x_t[25] = 26'b11111111101111010011111001;
        x_t[26] = 26'b11111111110110011101011000;
        x_t[27] = 26'b11111111110100110011001111;
        x_t[28] = 26'b11111111101111011111100010;
        x_t[29] = 26'b11111111110001101111111100;
        x_t[30] = 26'b11111111111010010000010011;
        x_t[31] = 26'b11111111110111000101100001;
        x_t[32] = 26'b11111111110111101001000101;
        x_t[33] = 26'b11111111111001011100010001;
        x_t[34] = 26'b11111111111100101000101111;
        x_t[35] = 26'b11111111111010000001010101;
        x_t[36] = 26'b11111111110110111001111011;
        x_t[37] = 26'b11111111111000101010100111;
        x_t[38] = 26'b11111111110110001100000010;
        x_t[39] = 26'b11111111111011010011000000;
        x_t[40] = 26'b11111111101101001010100001;
        x_t[41] = 26'b11111111111101000101000011;
        x_t[42] = 26'b11111111100111011100010000;
        x_t[43] = 26'b11111111111011101010110000;
        x_t[44] = 26'b11111111110100010111110100;
        x_t[45] = 26'b11111111110110010011001001;
        x_t[46] = 26'b11111111111000101011001000;
        x_t[47] = 26'b11111111110110110010011011;
        x_t[48] = 26'b11111111111000101110110001;
        x_t[49] = 26'b11111111111001010110110100;
        x_t[50] = 26'b11111111111010100011110011;
        x_t[51] = 26'b11111111111111001111010110;
        x_t[52] = 26'b11111111111100111100101101;
        x_t[53] = 26'b11111111111110110110110011;
        x_t[54] = 26'b11111111111101101100010101;
        x_t[55] = 26'b11111111111100000011011100;
        x_t[56] = 26'b11111111111010101100111111;
        x_t[57] = 26'b00000000000000101010010100;
        x_t[58] = 26'b00000000000010001000111011;
        x_t[59] = 26'b00000000000001111011010100;
        x_t[60] = 26'b11111111111110000001111010;
        x_t[61] = 26'b11111111111101000111011010;
        x_t[62] = 26'b11111111110101100011111000;
        x_t[63] = 26'b11111111111110111010101011;
        
        h_t_prev[0] = 26'b11111111110101011110010000;
        h_t_prev[1] = 26'b11111111111010111101011000;
        h_t_prev[2] = 26'b11111111111010000010000111;
        h_t_prev[3] = 26'b11111111111110101000110101;
        h_t_prev[4] = 26'b11111111111111010011101111;
        h_t_prev[5] = 26'b00000000000000001011110001;
        h_t_prev[6] = 26'b11111111111010101111100001;
        h_t_prev[7] = 26'b11111111111011111001100100;
        h_t_prev[8] = 26'b11111111111010010011001101;
        h_t_prev[9] = 26'b11111111111010001010100010;
        h_t_prev[10] = 26'b11111111111010100010000101;
        h_t_prev[11] = 26'b00000000000000100101011000;
        h_t_prev[12] = 26'b11111111111101010001101110;
        h_t_prev[13] = 26'b11111111111011110111101100;
        h_t_prev[14] = 26'b11111111110101011111000110;
        h_t_prev[15] = 26'b11111111110110010100000000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 80 timeout!");
                $fdisplay(fd_cycles, "Test Vector  80: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  80: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 80");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 81
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000111000010111010;
        x_t[1] = 26'b00000000000111001100011110;
        x_t[2] = 26'b00000000000010110101011000;
        x_t[3] = 26'b00000000000110001100001111;
        x_t[4] = 26'b00000000000111110101010110;
        x_t[5] = 26'b00000000000011101001101010;
        x_t[6] = 26'b00000000000011101100000101;
        x_t[7] = 26'b00000000000001101000000010;
        x_t[8] = 26'b00000000000100111011111110;
        x_t[9] = 26'b00000000000110000100001110;
        x_t[10] = 26'b00000000001000100110010010;
        x_t[11] = 26'b00000000000000111001110000;
        x_t[12] = 26'b00000000000101101100001101;
        x_t[13] = 26'b00000000001000001110001001;
        x_t[14] = 26'b00000000000101101000101100;
        x_t[15] = 26'b00000000000101111000101111;
        x_t[16] = 26'b00000000000110010010001111;
        x_t[17] = 26'b00000000000101011111000100;
        x_t[18] = 26'b00000000000101011100111000;
        x_t[19] = 26'b00000000000111111000000100;
        x_t[20] = 26'b00000000000100000001010111;
        x_t[21] = 26'b00000000000010001111000001;
        x_t[22] = 26'b00000000000010111110101000;
        x_t[23] = 26'b11111111111101111100100111;
        x_t[24] = 26'b11111111111101010000111000;
        x_t[25] = 26'b11111111111101111000010001;
        x_t[26] = 26'b11111111111101110110011111;
        x_t[27] = 26'b11111111111110101000000111;
        x_t[28] = 26'b00000000000001111111011110;
        x_t[29] = 26'b00000000000011001010101100;
        x_t[30] = 26'b11111111111110001010000101;
        x_t[31] = 26'b11111111111010111101111010;
        x_t[32] = 26'b11111111111110011101001101;
        x_t[33] = 26'b11111111111101011111010100;
        x_t[34] = 26'b11111111111100000010101001;
        x_t[35] = 26'b11111111111101011010011100;
        x_t[36] = 26'b11111111111101101111010010;
        x_t[37] = 26'b00000000000011111000001001;
        x_t[38] = 26'b11111111111110000100010001;
        x_t[39] = 26'b00000000000101110111000111;
        x_t[40] = 26'b11111111111111100000011011;
        x_t[41] = 26'b11111111110111110111001111;
        x_t[42] = 26'b11111111111101010011100001;
        x_t[43] = 26'b00000000001110110111100100;
        x_t[44] = 26'b11111111111000100011111100;
        x_t[45] = 26'b00000000001010100111001000;
        x_t[46] = 26'b00000000000100000000011011;
        x_t[47] = 26'b00000000000011100010000010;
        x_t[48] = 26'b00000000000100010110000100;
        x_t[49] = 26'b00000000000100000100100100;
        x_t[50] = 26'b00000000000110101111000001;
        x_t[51] = 26'b00000000000111101100010001;
        x_t[52] = 26'b00000000000110100010100101;
        x_t[53] = 26'b00000000000101011101111011;
        x_t[54] = 26'b00000000000011101011111000;
        x_t[55] = 26'b00000000000101001110011001;
        x_t[56] = 26'b00000000000011100100001010;
        x_t[57] = 26'b00000000001001001011111111;
        x_t[58] = 26'b00000000001010100101110011;
        x_t[59] = 26'b00000000001011010011010011;
        x_t[60] = 26'b00000000001011011100101001;
        x_t[61] = 26'b00000000010010010100110100;
        x_t[62] = 26'b00000000001001001101011100;
        x_t[63] = 26'b00000000000111101101111110;
        
        h_t_prev[0] = 26'b00000000000111000010111010;
        h_t_prev[1] = 26'b00000000000111001100011110;
        h_t_prev[2] = 26'b00000000000010110101011000;
        h_t_prev[3] = 26'b00000000000110001100001111;
        h_t_prev[4] = 26'b00000000000111110101010110;
        h_t_prev[5] = 26'b00000000000011101001101010;
        h_t_prev[6] = 26'b00000000000011101100000101;
        h_t_prev[7] = 26'b00000000000001101000000010;
        h_t_prev[8] = 26'b00000000000100111011111110;
        h_t_prev[9] = 26'b00000000000110000100001110;
        h_t_prev[10] = 26'b00000000001000100110010010;
        h_t_prev[11] = 26'b00000000000000111001110000;
        h_t_prev[12] = 26'b00000000000101101100001101;
        h_t_prev[13] = 26'b00000000001000001110001001;
        h_t_prev[14] = 26'b00000000000101101000101100;
        h_t_prev[15] = 26'b00000000000101111000101111;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 81 timeout!");
                $fdisplay(fd_cycles, "Test Vector  81: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  81: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 81");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 82
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000010011010111100;
        x_t[1] = 26'b00000000000011001101111110;
        x_t[2] = 26'b00000000000000011010000000;
        x_t[3] = 26'b00000000000100111110111001;
        x_t[4] = 26'b00000000000110010000010100;
        x_t[5] = 26'b00000000000000001011110001;
        x_t[6] = 26'b11111111111111000001010110;
        x_t[7] = 26'b11111111111101011111010111;
        x_t[8] = 26'b00000000000001101101101011;
        x_t[9] = 26'b00000000000100100000000000;
        x_t[10] = 26'b00000000000110011101010011;
        x_t[11] = 26'b00000000000001100010100001;
        x_t[12] = 26'b00000000000011001000010101;
        x_t[13] = 26'b00000000000011100010010100;
        x_t[14] = 26'b00000000000010111111111100;
        x_t[15] = 26'b00000000000001110000010011;
        x_t[16] = 26'b00000000000010111000001001;
        x_t[17] = 26'b00000000000011000001001001;
        x_t[18] = 26'b00000000000011110011011101;
        x_t[19] = 26'b00000000000101011110010011;
        x_t[20] = 26'b00000000000000111001001001;
        x_t[21] = 26'b00000000000011100111011011;
        x_t[22] = 26'b00000000000100010111011110;
        x_t[23] = 26'b00000000000000000111110101;
        x_t[24] = 26'b11111111111110000001100110;
        x_t[25] = 26'b11111111111110010001001000;
        x_t[26] = 26'b00000000000000001110100100;
        x_t[27] = 26'b00000000000000010110001010;
        x_t[28] = 26'b00000000000011001011000010;
        x_t[29] = 26'b00000000000001010110001110;
        x_t[30] = 26'b11111111111101111010011110;
        x_t[31] = 26'b11111111111100000100111000;
        x_t[32] = 26'b00000000000000101110100101;
        x_t[33] = 26'b00000000000000101010110110;
        x_t[34] = 26'b11111111111110011011000011;
        x_t[35] = 26'b11111111111110010101101001;
        x_t[36] = 26'b11111111111100001011111000;
        x_t[37] = 26'b00000000000010110110111010;
        x_t[38] = 26'b11111111111100011111011011;
        x_t[39] = 26'b11111111111111111000111110;
        x_t[40] = 26'b00000000000000001011111001;
        x_t[41] = 26'b11111111101100111111110010;
        x_t[42] = 26'b11111111110110101000100111;
        x_t[43] = 26'b00000000001000000000101101;
        x_t[44] = 26'b11111111110101110001001100;
        x_t[45] = 26'b00000000010000011010100100;
        x_t[46] = 26'b00000000000001101111010111;
        x_t[47] = 26'b00000000000001101010101011;
        x_t[48] = 26'b00000000000011011100111000;
        x_t[49] = 26'b00000000000100000100100100;
        x_t[50] = 26'b00000000000101100010111111;
        x_t[51] = 26'b00000000000111101100010001;
        x_t[52] = 26'b00000000000110001110001000;
        x_t[53] = 26'b00000000000101110100001100;
        x_t[54] = 26'b00000000000110101011101010;
        x_t[55] = 26'b00000000000100101011110111;
        x_t[56] = 26'b00000000000011000001110010;
        x_t[57] = 26'b00000000001000011000110101;
        x_t[58] = 26'b00000000001001001110100100;
        x_t[59] = 26'b00000000001100000010101010;
        x_t[60] = 26'b00000000001011101011111111;
        x_t[61] = 26'b00000000001111111111110101;
        x_t[62] = 26'b00000000000100110100010110;
        x_t[63] = 26'b00000000001000110100011000;
        
        h_t_prev[0] = 26'b00000000000010011010111100;
        h_t_prev[1] = 26'b00000000000011001101111110;
        h_t_prev[2] = 26'b00000000000000011010000000;
        h_t_prev[3] = 26'b00000000000100111110111001;
        h_t_prev[4] = 26'b00000000000110010000010100;
        h_t_prev[5] = 26'b00000000000000001011110001;
        h_t_prev[6] = 26'b11111111111111000001010110;
        h_t_prev[7] = 26'b11111111111101011111010111;
        h_t_prev[8] = 26'b00000000000001101101101011;
        h_t_prev[9] = 26'b00000000000100100000000000;
        h_t_prev[10] = 26'b00000000000110011101010011;
        h_t_prev[11] = 26'b00000000000001100010100001;
        h_t_prev[12] = 26'b00000000000011001000010101;
        h_t_prev[13] = 26'b00000000000011100010010100;
        h_t_prev[14] = 26'b00000000000010111111111100;
        h_t_prev[15] = 26'b00000000000001110000010011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 82 timeout!");
                $fdisplay(fd_cycles, "Test Vector  82: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  82: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 82");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 83
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111111101011111010000;
        x_t[1] = 26'b00000000000000001010001100;
        x_t[2] = 26'b00000000000000000110100101;
        x_t[3] = 26'b00000000000110001100001111;
        x_t[4] = 26'b00000000000110111000101110;
        x_t[5] = 26'b00000000000000001011110001;
        x_t[6] = 26'b11111111111101000100111000;
        x_t[7] = 26'b11111111110111011100100011;
        x_t[8] = 26'b11111111111100111000001111;
        x_t[9] = 26'b00000000000010100111101111;
        x_t[10] = 26'b00000000000111101011100101;
        x_t[11] = 26'b11111111111111111100100111;
        x_t[12] = 26'b00000000000001101010101011;
        x_t[13] = 26'b00000000000011000111000011;
        x_t[14] = 26'b11111111111011011010110010;
        x_t[15] = 26'b11111111111111001101100100;
        x_t[16] = 26'b00000000000001000001001011;
        x_t[17] = 26'b00000000000001110010001100;
        x_t[18] = 26'b00000000000001110100111101;
        x_t[19] = 26'b00000000000010101110100100;
        x_t[20] = 26'b11111111111111010101000010;
        x_t[21] = 26'b11111111111110011011111010;
        x_t[22] = 26'b11111111111110110100000101;
        x_t[23] = 26'b11111111111011110001011001;
        x_t[24] = 26'b11111111110110011010011011;
        x_t[25] = 26'b11111111110111000101001010;
        x_t[26] = 26'b11111111111010001001111011;
        x_t[27] = 26'b11111111111010101100100100;
        x_t[28] = 26'b11111111111111000010100010;
        x_t[29] = 26'b11111111111000110001001011;
        x_t[30] = 26'b11111111110100101001010001;
        x_t[31] = 26'b11111111110110110011110001;
        x_t[32] = 26'b11111111111001010110000111;
        x_t[33] = 26'b11111111111010010011110010;
        x_t[34] = 26'b11111111110111110111111010;
        x_t[35] = 26'b11111111110110111011111100;
        x_t[36] = 26'b11111111110100000111000001;
        x_t[37] = 26'b11111111111100001110111011;
        x_t[38] = 26'b11111111110011101010101011;
        x_t[39] = 26'b11111111111101001000100101;
        x_t[40] = 26'b11111111110010010000100110;
        x_t[41] = 26'b11111111110010001101100110;
        x_t[42] = 26'b11111111110001000100111000;
        x_t[43] = 26'b11111111111111000110001100;
        x_t[44] = 26'b11111111110000001011101101;
        x_t[45] = 26'b00000000001111011100101010;
        x_t[46] = 26'b11111111111011111010010111;
        x_t[47] = 26'b11111111111110001111110111;
        x_t[48] = 26'b11111111111111111000001011;
        x_t[49] = 26'b00000000000001001011001110;
        x_t[50] = 26'b00000000000001011000111011;
        x_t[51] = 26'b00000000000010010000100010;
        x_t[52] = 26'b00000000000001000110101110;
        x_t[53] = 26'b00000000000010010101100000;
        x_t[54] = 26'b00000000000110101011101010;
        x_t[55] = 26'b00000000000101001110011001;
        x_t[56] = 26'b00000000000001101011110110;
        x_t[57] = 26'b00000000000100101010000110;
        x_t[58] = 26'b00000000000101011010010011;
        x_t[59] = 26'b00000000001011110010111000;
        x_t[60] = 26'b00000000001010011111010100;
        x_t[61] = 26'b00000000001110001011111101;
        x_t[62] = 26'b00000000000001000111100111;
        x_t[63] = 26'b00000000001000100010110001;
        
        h_t_prev[0] = 26'b11111111111101011111010000;
        h_t_prev[1] = 26'b00000000000000001010001100;
        h_t_prev[2] = 26'b00000000000000000110100101;
        h_t_prev[3] = 26'b00000000000110001100001111;
        h_t_prev[4] = 26'b00000000000110111000101110;
        h_t_prev[5] = 26'b00000000000000001011110001;
        h_t_prev[6] = 26'b11111111111101000100111000;
        h_t_prev[7] = 26'b11111111110111011100100011;
        h_t_prev[8] = 26'b11111111111100111000001111;
        h_t_prev[9] = 26'b00000000000010100111101111;
        h_t_prev[10] = 26'b00000000000111101011100101;
        h_t_prev[11] = 26'b11111111111111111100100111;
        h_t_prev[12] = 26'b00000000000001101010101011;
        h_t_prev[13] = 26'b00000000000011000111000011;
        h_t_prev[14] = 26'b11111111111011011010110010;
        h_t_prev[15] = 26'b11111111111111001101100100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 83 timeout!");
                $fdisplay(fd_cycles, "Test Vector  83: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  83: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 83");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 84
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111110110101101001011;
        x_t[1] = 26'b11111111111001101111000100;
        x_t[2] = 26'b11111111111000110100011011;
        x_t[3] = 26'b11111111111110000010001010;
        x_t[4] = 26'b11111111111110111111100001;
        x_t[5] = 26'b11111111111000001101011100;
        x_t[6] = 26'b11111111110100100001001101;
        x_t[7] = 26'b11111111110000011100101010;
        x_t[8] = 26'b11111111111000000010110011;
        x_t[9] = 26'b11111111111100111110111011;
        x_t[10] = 26'b00000000000001110111110000;
        x_t[11] = 26'b11111111110111000001110111;
        x_t[12] = 26'b11111111111010010110011011;
        x_t[13] = 26'b11111111111110110110011111;
        x_t[14] = 26'b11111111111011011010110010;
        x_t[15] = 26'b11111111111110010000100010;
        x_t[16] = 26'b11111111111101100111000101;
        x_t[17] = 26'b11111111111101001010000110;
        x_t[18] = 26'b11111111111010111010001100;
        x_t[19] = 26'b11111111111011110111001110;
        x_t[20] = 26'b11111111111001011101100111;
        x_t[21] = 26'b11111111111101000011011111;
        x_t[22] = 26'b11111111111100001111000100;
        x_t[23] = 26'b11111111111000010100111101;
        x_t[24] = 26'b11111111110110001110010000;
        x_t[25] = 26'b11111111110101111010100100;
        x_t[26] = 26'b11111111110111010000000100;
        x_t[27] = 26'b11111111110110100001010010;
        x_t[28] = 26'b11111111111010101101011101;
        x_t[29] = 26'b11111111111001110011101110;
        x_t[30] = 26'b11111111110101011000000110;
        x_t[31] = 26'b11111111110010101001101000;
        x_t[32] = 26'b11111111111000001101011011;
        x_t[33] = 26'b11111111110111001000010000;
        x_t[34] = 26'b11111111110100010011010010;
        x_t[35] = 26'b11111111110101011001010000;
        x_t[36] = 26'b11111111110001000000001110;
        x_t[37] = 26'b11111111111000111010111011;
        x_t[38] = 26'b11111111110111110000111000;
        x_t[39] = 26'b00000000000001010001001010;
        x_t[40] = 26'b11111111111101011101111111;
        x_t[41] = 26'b11111111111110011000100000;
        x_t[42] = 26'b11111111111000110110111010;
        x_t[43] = 26'b11111111110110001011101011;
        x_t[44] = 26'b11111111110101000100100000;
        x_t[45] = 26'b00000000000111001110011110;
        x_t[46] = 26'b00000000000001000101111010;
        x_t[47] = 26'b00000000000000101111000000;
        x_t[48] = 26'b11111111111110000101110101;
        x_t[49] = 26'b11111111111111011100000001;
        x_t[50] = 26'b11111111111100010101110101;
        x_t[51] = 26'b11111111111011111010110110;
        x_t[52] = 26'b11111111111010000100100011;
        x_t[53] = 26'b11111111111011101110011000;
        x_t[54] = 26'b00000000000011010011111010;
        x_t[55] = 26'b00000000000110110101111110;
        x_t[56] = 26'b00000000000001001001011110;
        x_t[57] = 26'b11111111111111010101000011;
        x_t[58] = 26'b00000000000001010100100101;
        x_t[59] = 26'b00000000001100000010101010;
        x_t[60] = 26'b00000000001010011111010100;
        x_t[61] = 26'b00000000001101001001101111;
        x_t[62] = 26'b11111111111111111101101001;
        x_t[63] = 26'b00000000001000010001001011;
        
        h_t_prev[0] = 26'b11111111110110101101001011;
        h_t_prev[1] = 26'b11111111111001101111000100;
        h_t_prev[2] = 26'b11111111111000110100011011;
        h_t_prev[3] = 26'b11111111111110000010001010;
        h_t_prev[4] = 26'b11111111111110111111100001;
        h_t_prev[5] = 26'b11111111111000001101011100;
        h_t_prev[6] = 26'b11111111110100100001001101;
        h_t_prev[7] = 26'b11111111110000011100101010;
        h_t_prev[8] = 26'b11111111111000000010110011;
        h_t_prev[9] = 26'b11111111111100111110111011;
        h_t_prev[10] = 26'b00000000000001110111110000;
        h_t_prev[11] = 26'b11111111110111000001110111;
        h_t_prev[12] = 26'b11111111111010010110011011;
        h_t_prev[13] = 26'b11111111111110110110011111;
        h_t_prev[14] = 26'b11111111111011011010110010;
        h_t_prev[15] = 26'b11111111111110010000100010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 84 timeout!");
                $fdisplay(fd_cycles, "Test Vector  84: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  84: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 84");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 85
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111111010011001111100;
        x_t[1] = 26'b11111111111100110010110110;
        x_t[2] = 26'b11111111111000001101100101;
        x_t[3] = 26'b11111111111011000000110011;
        x_t[4] = 26'b11111111111011001101000010;
        x_t[5] = 26'b11111111110101011011111100;
        x_t[6] = 26'b11111111110101010011000000;
        x_t[7] = 26'b11111111110101110110110000;
        x_t[8] = 26'b11111111111010010011001101;
        x_t[9] = 26'b11111111111011101110110000;
        x_t[10] = 26'b11111111111101111001010110;
        x_t[11] = 26'b11111111110100001010011010;
        x_t[12] = 26'b11111111110101100110000011;
        x_t[13] = 26'b11111111111100101110001101;
        x_t[14] = 26'b11111111111101011001010110;
        x_t[15] = 26'b11111111111110100100111000;
        x_t[16] = 26'b11111111111011011100010010;
        x_t[17] = 26'b11111111111000100001111111;
        x_t[18] = 26'b11111111110100010100100001;
        x_t[19] = 26'b11111111110100111111111000;
        x_t[20] = 26'b11111111110010011011000111;
        x_t[21] = 26'b11111111111011001001111011;
        x_t[22] = 26'b11111111111001010000101011;
        x_t[23] = 26'b11111111110110010101010110;
        x_t[24] = 26'b11111111110011111100000110;
        x_t[25] = 26'b11111111110011111110010000;
        x_t[26] = 26'b11111111110100000101010011;
        x_t[27] = 26'b11111111110100100011100001;
        x_t[28] = 26'b11111111111001101110011110;
        x_t[29] = 26'b11111111110101101001100001;
        x_t[30] = 26'b11111111110011001011100110;
        x_t[31] = 26'b11111111110001110100011010;
        x_t[32] = 26'b11111111110110100000011001;
        x_t[33] = 26'b11111111110100001111001110;
        x_t[34] = 26'b11111111110001010100110000;
        x_t[35] = 26'b11111111110010100111100111;
        x_t[36] = 26'b11111111101111110000101101;
        x_t[37] = 26'b11111111110110111000011101;
        x_t[38] = 26'b11111111110100111011010110;
        x_t[39] = 26'b11111111111011010011000000;
        x_t[40] = 26'b11111111110110101011001101;
        x_t[41] = 26'b11111111110010001101100110;
        x_t[42] = 26'b11111111110011010011001011;
        x_t[43] = 26'b00000000001000000000101101;
        x_t[44] = 26'b11111111110101011010110110;
        x_t[45] = 26'b00000000000100010100110000;
        x_t[46] = 26'b00000000000001000101111010;
        x_t[47] = 26'b00000000000000000111001101;
        x_t[48] = 26'b11111111111100000000011010;
        x_t[49] = 26'b11111111111101011010010010;
        x_t[50] = 26'b11111111111000011110110001;
        x_t[51] = 26'b11111111110111111111101101;
        x_t[52] = 26'b11111111110110001111000000;
        x_t[53] = 26'b11111111111001111111000010;
        x_t[54] = 26'b00000000000010100011111110;
        x_t[55] = 26'b00000000000011100110110100;
        x_t[56] = 26'b11111111111110101110110011;
        x_t[57] = 26'b11111111111010110011001010;
        x_t[58] = 26'b11111111111111001001000000;
        x_t[59] = 26'b00000000001101000001110100;
        x_t[60] = 26'b00000000001001010010101001;
        x_t[61] = 26'b00000000001011100110011010;
        x_t[62] = 26'b00000000000001110100000000;
        x_t[63] = 26'b00000000001000010001001011;
        
        h_t_prev[0] = 26'b11111111111010011001111100;
        h_t_prev[1] = 26'b11111111111100110010110110;
        h_t_prev[2] = 26'b11111111111000001101100101;
        h_t_prev[3] = 26'b11111111111011000000110011;
        h_t_prev[4] = 26'b11111111111011001101000010;
        h_t_prev[5] = 26'b11111111110101011011111100;
        h_t_prev[6] = 26'b11111111110101010011000000;
        h_t_prev[7] = 26'b11111111110101110110110000;
        h_t_prev[8] = 26'b11111111111010010011001101;
        h_t_prev[9] = 26'b11111111111011101110110000;
        h_t_prev[10] = 26'b11111111111101111001010110;
        h_t_prev[11] = 26'b11111111110100001010011010;
        h_t_prev[12] = 26'b11111111110101100110000011;
        h_t_prev[13] = 26'b11111111111100101110001101;
        h_t_prev[14] = 26'b11111111111101011001010110;
        h_t_prev[15] = 26'b11111111111110100100111000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 85 timeout!");
                $fdisplay(fd_cycles, "Test Vector  85: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  85: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 85");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 86
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111111010011001111100;
        x_t[1] = 26'b11111111111101000110011011;
        x_t[2] = 26'b11111111111001011011010001;
        x_t[3] = 26'b11111111111010101101011101;
        x_t[4] = 26'b11111111111100110010000100;
        x_t[5] = 26'b11111111111000001101011100;
        x_t[6] = 26'b11111111110110011101101011;
        x_t[7] = 26'b11111111111001010110101101;
        x_t[8] = 26'b11111111111101001100110111;
        x_t[9] = 26'b11111111111101111011000100;
        x_t[10] = 26'b11111111111110110100000011;
        x_t[11] = 26'b11111111110110011001000110;
        x_t[12] = 26'b11111111110111110010100010;
        x_t[13] = 26'b11111111111100101110001101;
        x_t[14] = 26'b00000000000001000001011000;
        x_t[15] = 26'b00000000000001110000010011;
        x_t[16] = 26'b11111111111101010011010000;
        x_t[17] = 26'b11111111111010000100101100;
        x_t[18] = 26'b11111111110101111101111100;
        x_t[19] = 26'b11111111110110101101101101;
        x_t[20] = 26'b11111111110011111111001111;
        x_t[21] = 26'b11111111111101111010110000;
        x_t[22] = 26'b11111111111011001111100111;
        x_t[23] = 26'b11111111110110111000001001;
        x_t[24] = 26'b11111111110110111110111101;
        x_t[25] = 26'b11111111110110111000101110;
        x_t[26] = 26'b11111111110111010000000100;
        x_t[27] = 26'b11111111110110110001000001;
        x_t[28] = 26'b11111111111001100001111000;
        x_t[29] = 26'b11111111111010110110010001;
        x_t[30] = 26'b11111111110111010100111110;
        x_t[31] = 26'b11111111110110110011110001;
        x_t[32] = 26'b11111111111010110000111110;
        x_t[33] = 26'b11111111111000110111010001;
        x_t[34] = 26'b11111111110110101011101101;
        x_t[35] = 26'b11111111111000001010111001;
        x_t[36] = 26'b11111111110101010110100010;
        x_t[37] = 26'b11111111111001111100001010;
        x_t[38] = 26'b11111111111010010010001111;
        x_t[39] = 26'b11111111111111111000111110;
        x_t[40] = 26'b11111111111110110100111100;
        x_t[41] = 26'b11111111101111100110101100;
        x_t[42] = 26'b11111111111111001010000110;
        x_t[43] = 26'b00000000001000000000101101;
        x_t[44] = 26'b11111111111100110000000100;
        x_t[45] = 26'b00000000001001001010010010;
        x_t[46] = 26'b00000000000100010101001001;
        x_t[47] = 26'b00000000000010100110010111;
        x_t[48] = 26'b11111111111110101011111100;
        x_t[49] = 26'b11111111111110010001111001;
        x_t[50] = 26'b11111111111001000100110001;
        x_t[51] = 26'b11111111111000010011000001;
        x_t[52] = 26'b11111111110111001100011001;
        x_t[53] = 26'b11111111111011011000000111;
        x_t[54] = 26'b00000000000001000100000101;
        x_t[55] = 26'b00000000000011000100010010;
        x_t[56] = 26'b11111111111110001100011011;
        x_t[57] = 26'b11111111111001101110111101;
        x_t[58] = 26'b11111111111101110001110001;
        x_t[59] = 26'b00000000001001010100111111;
        x_t[60] = 26'b00000000000111110110101000;
        x_t[61] = 26'b00000000001000110000010101;
        x_t[62] = 26'b00000000000010010001100110;
        x_t[63] = 26'b00000000000110010101111101;
        
        h_t_prev[0] = 26'b11111111111010011001111100;
        h_t_prev[1] = 26'b11111111111101000110011011;
        h_t_prev[2] = 26'b11111111111001011011010001;
        h_t_prev[3] = 26'b11111111111010101101011101;
        h_t_prev[4] = 26'b11111111111100110010000100;
        h_t_prev[5] = 26'b11111111111000001101011100;
        h_t_prev[6] = 26'b11111111110110011101101011;
        h_t_prev[7] = 26'b11111111111001010110101101;
        h_t_prev[8] = 26'b11111111111101001100110111;
        h_t_prev[9] = 26'b11111111111101111011000100;
        h_t_prev[10] = 26'b11111111111110110100000011;
        h_t_prev[11] = 26'b11111111110110011001000110;
        h_t_prev[12] = 26'b11111111110111110010100010;
        h_t_prev[13] = 26'b11111111111100101110001101;
        h_t_prev[14] = 26'b00000000000001000001011000;
        h_t_prev[15] = 26'b00000000000001110000010011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 86 timeout!");
                $fdisplay(fd_cycles, "Test Vector  86: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  86: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 86");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 87
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000000100100100100;
        x_t[1] = 26'b00000000000001011000100000;
        x_t[2] = 26'b11111111111101000100010110;
        x_t[3] = 26'b11111111111101011011011111;
        x_t[4] = 26'b00000000000000111000110001;
        x_t[5] = 26'b11111111111110110011000001;
        x_t[6] = 26'b11111111111111011010010000;
        x_t[7] = 26'b11111111111101011111010111;
        x_t[8] = 26'b00000000000000000110100010;
        x_t[9] = 26'b00000000000001000011100000;
        x_t[10] = 26'b00000000000010001011010100;
        x_t[11] = 26'b11111111111001111001010100;
        x_t[12] = 26'b11111111111111011110001100;
        x_t[13] = 26'b00000000000100011000110101;
        x_t[14] = 26'b00000000000100101001011010;
        x_t[15] = 26'b00000000000011010110000000;
        x_t[16] = 26'b11111111111111110001111000;
        x_t[17] = 26'b11111111111100100010100111;
        x_t[18] = 26'b11111111111010111010001100;
        x_t[19] = 26'b11111111111100100011001001;
        x_t[20] = 26'b11111111111010101000101101;
        x_t[21] = 26'b00000000000011011100011000;
        x_t[22] = 26'b00000000000001100101110001;
        x_t[23] = 26'b11111111111101000010100110;
        x_t[24] = 26'b11111111111100111000100001;
        x_t[25] = 26'b11111111111100101101101011;
        x_t[26] = 26'b11111111111011001101100001;
        x_t[27] = 26'b11111111111101011001100000;
        x_t[28] = 26'b11111111111111101000010101;
        x_t[29] = 26'b00000000000010011000110010;
        x_t[30] = 26'b11111111111101101010110111;
        x_t[31] = 26'b11111111111001100101001100;
        x_t[32] = 26'b11111111111101000010010110;
        x_t[33] = 26'b11111111111010100110010010;
        x_t[34] = 26'b11111111111001101010001110;
        x_t[35] = 26'b11111111111011110111110000;
        x_t[36] = 26'b11111111111100001011111000;
        x_t[37] = 26'b11111111111111100010111011;
        x_t[38] = 26'b00000000000000100101101000;
        x_t[39] = 26'b00000000001010111010011111;
        x_t[40] = 26'b00000000000111111111111001;
        x_t[41] = 26'b00000000000010010010111000;
        x_t[42] = 26'b00000000000011100110101100;
        x_t[43] = 26'b00000000001000101100100101;
        x_t[44] = 26'b11111111111111001100011110;
        x_t[45] = 26'b00000000001100100010111100;
        x_t[46] = 26'b00000000000110010001011110;
        x_t[47] = 26'b00000000000101011001011001;
        x_t[48] = 26'b00000000000000110001010111;
        x_t[49] = 26'b11111111111111101110100100;
        x_t[50] = 26'b11111111111011011100110100;
        x_t[51] = 26'b11111111111000111001101010;
        x_t[52] = 26'b11111111111000110010101101;
        x_t[53] = 26'b11111111111101000111011101;
        x_t[54] = 26'b11111111111111100100001100;
        x_t[55] = 26'b00000000000100101011110111;
        x_t[56] = 26'b00000000000001001001011110;
        x_t[57] = 26'b11111111111010010001000100;
        x_t[58] = 26'b11111111111011000011010010;
        x_t[59] = 26'b00000000000010111010011110;
        x_t[60] = 26'b00000000000100101111010010;
        x_t[61] = 26'b00000000000010100011000010;
        x_t[62] = 26'b11111111111100010000111011;
        x_t[63] = 26'b11111111111111101111011111;
        
        h_t_prev[0] = 26'b00000000000000100100100100;
        h_t_prev[1] = 26'b00000000000001011000100000;
        h_t_prev[2] = 26'b11111111111101000100010110;
        h_t_prev[3] = 26'b11111111111101011011011111;
        h_t_prev[4] = 26'b00000000000000111000110001;
        h_t_prev[5] = 26'b11111111111110110011000001;
        h_t_prev[6] = 26'b11111111111111011010010000;
        h_t_prev[7] = 26'b11111111111101011111010111;
        h_t_prev[8] = 26'b00000000000000000110100010;
        h_t_prev[9] = 26'b00000000000001000011100000;
        h_t_prev[10] = 26'b00000000000010001011010100;
        h_t_prev[11] = 26'b11111111111001111001010100;
        h_t_prev[12] = 26'b11111111111111011110001100;
        h_t_prev[13] = 26'b00000000000100011000110101;
        h_t_prev[14] = 26'b00000000000100101001011010;
        h_t_prev[15] = 26'b00000000000011010110000000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 87 timeout!");
                $fdisplay(fd_cycles, "Test Vector  87: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  87: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 87");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 88
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000011111101100110;
        x_t[1] = 26'b00000000000100001000101100;
        x_t[2] = 26'b11111111111111011111101111;
        x_t[3] = 26'b11111111111111110110001011;
        x_t[4] = 26'b00000000000010001001100110;
        x_t[5] = 26'b00000000000000001011110001;
        x_t[6] = 26'b00000000000000001100000010;
        x_t[7] = 26'b00000000000001111100011001;
        x_t[8] = 26'b00000000000011101001011101;
        x_t[9] = 26'b00000000000100110100000011;
        x_t[10] = 26'b00000000001000010010101110;
        x_t[11] = 26'b11111111111101011001100010;
        x_t[12] = 26'b00000000000011011111101111;
        x_t[13] = 26'b00000000000110111100010111;
        x_t[14] = 26'b00000000001010010000000001;
        x_t[15] = 26'b00000000000111110010110010;
        x_t[16] = 26'b00000000000100000111011101;
        x_t[17] = 26'b00000000000001001010101101;
        x_t[18] = 26'b11111111111111001100010010;
        x_t[19] = 26'b00000000000001000000101110;
        x_t[20] = 26'b11111111111110111100000000;
        x_t[21] = 26'b11111111111111010011001010;
        x_t[22] = 26'b00000000000000001100111011;
        x_t[23] = 26'b11111111111100001000100110;
        x_t[24] = 26'b11111111111010111110101111;
        x_t[25] = 26'b11111111111010100100111011;
        x_t[26] = 26'b11111111111000100100100011;
        x_t[27] = 26'b11111111111011111011001011;
        x_t[28] = 26'b11111111111111110100111011;
        x_t[29] = 26'b00000000000000000011000010;
        x_t[30] = 26'b11111111111010010000010011;
        x_t[31] = 26'b11111111111000011110001110;
        x_t[32] = 26'b11111111111100001011110101;
        x_t[33] = 26'b11111111111000110111010001;
        x_t[34] = 26'b11111111110110011000101001;
        x_t[35] = 26'b11111111111000011110101000;
        x_t[36] = 26'b11111111110111110101100100;
        x_t[37] = 26'b11111111111000111010111011;
        x_t[38] = 26'b11111111111111111101010010;
        x_t[39] = 26'b00000000000101011001101110;
        x_t[40] = 26'b00000000001100000100110000;
        x_t[41] = 26'b11111111110110111111100110;
        x_t[42] = 26'b11111111111000011111001101;
        x_t[43] = 26'b00000000001110110111100100;
        x_t[44] = 26'b00000000000010010101100011;
        x_t[45] = 26'b00000000001101100000110110;
        x_t[46] = 26'b00000000001110010111100010;
        x_t[47] = 26'b00000000001100110110110101;
        x_t[48] = 26'b00000000000110011011011110;
        x_t[49] = 26'b00000000000110101011010111;
        x_t[50] = 26'b00000000000000110010111010;
        x_t[51] = 26'b11111111111010101101100101;
        x_t[52] = 26'b11111111111010000100100011;
        x_t[53] = 26'b11111111111101000111011101;
        x_t[54] = 26'b11111111111101101100010101;
        x_t[55] = 26'b00000000001001000000000101;
        x_t[56] = 26'b00000000001000001000010101;
        x_t[57] = 26'b11111111111100111011100101;
        x_t[58] = 26'b11111111110110101100001000;
        x_t[59] = 26'b11111111111100000000011000;
        x_t[60] = 26'b00000000000100010000100111;
        x_t[61] = 26'b11111111111100100110010011;
        x_t[62] = 26'b11111111110010010100101111;
        x_t[63] = 26'b11111111111010110010101001;
        
        h_t_prev[0] = 26'b00000000000011111101100110;
        h_t_prev[1] = 26'b00000000000100001000101100;
        h_t_prev[2] = 26'b11111111111111011111101111;
        h_t_prev[3] = 26'b11111111111111110110001011;
        h_t_prev[4] = 26'b00000000000010001001100110;
        h_t_prev[5] = 26'b00000000000000001011110001;
        h_t_prev[6] = 26'b00000000000000001100000010;
        h_t_prev[7] = 26'b00000000000001111100011001;
        h_t_prev[8] = 26'b00000000000011101001011101;
        h_t_prev[9] = 26'b00000000000100110100000011;
        h_t_prev[10] = 26'b00000000001000010010101110;
        h_t_prev[11] = 26'b11111111111101011001100010;
        h_t_prev[12] = 26'b00000000000011011111101111;
        h_t_prev[13] = 26'b00000000000110111100010111;
        h_t_prev[14] = 26'b00000000001010010000000001;
        h_t_prev[15] = 26'b00000000000111110010110010;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 88 timeout!");
                $fdisplay(fd_cycles, "Test Vector  88: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  88: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 88");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 89
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000101100000010000;
        x_t[1] = 26'b00000000000100011100010001;
        x_t[2] = 26'b00000000000000101101011011;
        x_t[3] = 26'b00000000000010110111100010;
        x_t[4] = 26'b00000000000100101011010001;
        x_t[5] = 26'b11111111111111110101100101;
        x_t[6] = 26'b11111111111010010110101000;
        x_t[7] = 26'b00000000000100001010111001;
        x_t[8] = 26'b00000000000011010100110100;
        x_t[9] = 26'b00000000000101110000001011;
        x_t[10] = 26'b00000000001010101111010001;
        x_t[11] = 26'b11111111111111111100100111;
        x_t[12] = 26'b00000000000101010100110011;
        x_t[13] = 26'b00000000000111010111101000;
        x_t[14] = 26'b00000000001011001111010011;
        x_t[15] = 26'b00000000000111011110011100;
        x_t[16] = 26'b00000000000101111110011011;
        x_t[17] = 26'b00000000000100010000000111;
        x_t[18] = 26'b00000000000000110101101101;
        x_t[19] = 26'b00000000000001101100101010;
        x_t[20] = 26'b11111111111111010101000010;
        x_t[21] = 26'b11111111111101101111101100;
        x_t[22] = 26'b11111111111110100111011000;
        x_t[23] = 26'b11111111111010010100100101;
        x_t[24] = 26'b11111111111010100110011000;
        x_t[25] = 26'b11111111111010001100000100;
        x_t[26] = 26'b11111111111001101000001001;
        x_t[27] = 26'b11111111111001111101011001;
        x_t[28] = 26'b11111111111101000100100110;
        x_t[29] = 26'b00000000000000000011000010;
        x_t[30] = 26'b11111111111001010001110111;
        x_t[31] = 26'b11111111111001000001101101;
        x_t[32] = 26'b11111111111111000001100011;
        x_t[33] = 26'b11111111111100000010110011;
        x_t[34] = 26'b11111111111000011110000001;
        x_t[35] = 26'b11111111111011100100000001;
        x_t[36] = 26'b11111111110111001101110100;
        x_t[37] = 26'b11111111110110000111100010;
        x_t[38] = 26'b00000000000010001010011110;
        x_t[39] = 26'b00000000000000010110010111;
        x_t[40] = 26'b00000000000100111100001111;
        x_t[41] = 26'b11111111101100111111110010;
        x_t[42] = 26'b11111111111001100110010110;
        x_t[43] = 26'b00000000001000000000101101;
        x_t[44] = 26'b11111111111011010110101100;
        x_t[45] = 26'b00000000000110010000100100;
        x_t[46] = 26'b00000000000100111110100101;
        x_t[47] = 26'b00000000000110111100110111;
        x_t[48] = 26'b00000000000011001001110101;
        x_t[49] = 26'b00000000000100101001101000;
        x_t[50] = 26'b11111111111111000000111000;
        x_t[51] = 26'b11111111110101010001110110;
        x_t[52] = 26'b11111111110100111101001001;
        x_t[53] = 26'b11111111110011101110001011;
        x_t[54] = 26'b11111111110010011101001011;
        x_t[55] = 26'b00000000000001011100101101;
        x_t[56] = 26'b00000000000010110000100110;
        x_t[57] = 26'b11111111110110110011011000;
        x_t[58] = 26'b11111111101010001001100011;
        x_t[59] = 26'b11111111101001010000011010;
        x_t[60] = 26'b11111111111111111100100101;
        x_t[61] = 26'b11111111110011010010010111;
        x_t[62] = 26'b11111111100011000100010010;
        x_t[63] = 26'b11111111110001011100001001;
        
        h_t_prev[0] = 26'b00000000000101100000010000;
        h_t_prev[1] = 26'b00000000000100011100010001;
        h_t_prev[2] = 26'b00000000000000101101011011;
        h_t_prev[3] = 26'b00000000000010110111100010;
        h_t_prev[4] = 26'b00000000000100101011010001;
        h_t_prev[5] = 26'b11111111111111110101100101;
        h_t_prev[6] = 26'b11111111111010010110101000;
        h_t_prev[7] = 26'b00000000000100001010111001;
        h_t_prev[8] = 26'b00000000000011010100110100;
        h_t_prev[9] = 26'b00000000000101110000001011;
        h_t_prev[10] = 26'b00000000001010101111010001;
        h_t_prev[11] = 26'b11111111111111111100100111;
        h_t_prev[12] = 26'b00000000000101010100110011;
        h_t_prev[13] = 26'b00000000000111010111101000;
        h_t_prev[14] = 26'b00000000001011001111010011;
        h_t_prev[15] = 26'b00000000000111011110011100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 89 timeout!");
                $fdisplay(fd_cycles, "Test Vector  89: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  89: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 89");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 90
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000111000010111010;
        x_t[1] = 26'b00000000000110111000111001;
        x_t[2] = 26'b00000000000100101001111011;
        x_t[3] = 26'b00000000000111101100111011;
        x_t[4] = 26'b00000000001010010111000001;
        x_t[5] = 26'b00000000000101101110110010;
        x_t[6] = 26'b00000000000000001100000010;
        x_t[7] = 26'b00000000000000000010001111;
        x_t[8] = 26'b00000000000010010110111100;
        x_t[9] = 26'b00000000000111101000011100;
        x_t[10] = 26'b00000000001101110010111110;
        x_t[11] = 26'b00000000000110010100010001;
        x_t[12] = 26'b00000000000111001001110111;
        x_t[13] = 26'b00000000000110111100010111;
        x_t[14] = 26'b00000000000010000000101010;
        x_t[15] = 26'b00000000000011101010010110;
        x_t[16] = 26'b00000000000101000010111100;
        x_t[17] = 26'b00000000000100110111100101;
        x_t[18] = 26'b00000000000001011111111000;
        x_t[19] = 26'b11111111111111101000110111;
        x_t[20] = 26'b11111111111011110011110010;
        x_t[21] = 26'b00000000000001101101111000;
        x_t[22] = 26'b00000000000010100101001111;
        x_t[23] = 26'b11111111111111000010001110;
        x_t[24] = 26'b11111111111100010011111111;
        x_t[25] = 26'b11111111111100001000011000;
        x_t[26] = 26'b00000000000000001110100100;
        x_t[27] = 26'b00000000000000110101100111;
        x_t[28] = 26'b00000000000010110001110110;
        x_t[29] = 26'b11111111111101101101010011;
        x_t[30] = 26'b11111111111100111100000001;
        x_t[31] = 26'b11111111111111011001110011;
        x_t[32] = 26'b00000000000011110110011110;
        x_t[33] = 26'b00000000000011110110010111;
        x_t[34] = 26'b00000000000000001101010111;
        x_t[35] = 26'b00000000000001101110110001;
        x_t[36] = 26'b00000000000001001001111101;
        x_t[37] = 26'b00000000000001110101101100;
        x_t[38] = 26'b11111111111111000000110010;
        x_t[39] = 26'b00000000001011110101010001;
        x_t[40] = 26'b11111111111111001010101011;
        x_t[41] = 26'b11111111110001010101111110;
        x_t[42] = 26'b11111111110011010011001011;
        x_t[43] = 26'b00000000000000011101111101;
        x_t[44] = 26'b11111111110011101011001000;
        x_t[45] = 26'b00000000000010011000111101;
        x_t[46] = 26'b11111111111001010100100101;
        x_t[47] = 26'b11111111111101000000010010;
        x_t[48] = 26'b11111111111011011010010011;
        x_t[49] = 26'b11111111111111011100000001;
        x_t[50] = 26'b11111111111100010101110101;
        x_t[51] = 26'b11111111110000011100110000;
        x_t[52] = 26'b11111111101111100001010010;
        x_t[53] = 26'b11111111101011000001011100;
        x_t[54] = 26'b11111111100111111101111110;
        x_t[55] = 26'b11111111110111011101111101;
        x_t[56] = 26'b11111111111001000101111000;
        x_t[57] = 26'b11111111110000011010001000;
        x_t[58] = 26'b11111111100001011011001111;
        x_t[59] = 26'b11111111011010001101010001;
        x_t[60] = 26'b11111111110101101001001100;
        x_t[61] = 26'b11111111100101110101100100;
        x_t[62] = 26'b11111111010001011111110111;
        x_t[63] = 26'b11111111100010110111001101;
        
        h_t_prev[0] = 26'b00000000000111000010111010;
        h_t_prev[1] = 26'b00000000000110111000111001;
        h_t_prev[2] = 26'b00000000000100101001111011;
        h_t_prev[3] = 26'b00000000000111101100111011;
        h_t_prev[4] = 26'b00000000001010010111000001;
        h_t_prev[5] = 26'b00000000000101101110110010;
        h_t_prev[6] = 26'b00000000000000001100000010;
        h_t_prev[7] = 26'b00000000000000000010001111;
        h_t_prev[8] = 26'b00000000000010010110111100;
        h_t_prev[9] = 26'b00000000000111101000011100;
        h_t_prev[10] = 26'b00000000001101110010111110;
        h_t_prev[11] = 26'b00000000000110010100010001;
        h_t_prev[12] = 26'b00000000000111001001110111;
        h_t_prev[13] = 26'b00000000000110111100010111;
        h_t_prev[14] = 26'b00000000000010000000101010;
        h_t_prev[15] = 26'b00000000000011101010010110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 90 timeout!");
                $fdisplay(fd_cycles, "Test Vector  90: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  90: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 90");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 91
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000100010001010101;
        x_t[1] = 26'b00000000001001000001111100;
        x_t[2] = 26'b00000000001010101110011000;
        x_t[3] = 26'b00000000001110010110010100;
        x_t[4] = 26'b00000000001110011101101110;
        x_t[5] = 26'b00000000001000100000010010;
        x_t[6] = 26'b00000000000101101000100011;
        x_t[7] = 26'b00000000000000000010001111;
        x_t[8] = 26'b00000000000011111110000101;
        x_t[9] = 26'b00000000001100000001000100;
        x_t[10] = 26'b00000000010010111111101010;
        x_t[11] = 26'b00000000000111100101110100;
        x_t[12] = 26'b00000000000110000011101000;
        x_t[13] = 26'b00000000000101001111010110;
        x_t[14] = 26'b11111111111101011001010110;
        x_t[15] = 26'b00000000000011111110101100;
        x_t[16] = 26'b00000000000101111110011011;
        x_t[17] = 26'b00000000000110000110100011;
        x_t[18] = 26'b00000000000010001010000011;
        x_t[19] = 26'b11111111111110010000111111;
        x_t[20] = 26'b11111111111000101011100100;
        x_t[21] = 26'b00000000000011011100011000;
        x_t[22] = 26'b00000000000100001010110010;
        x_t[23] = 26'b00000000000001001101011100;
        x_t[24] = 26'b11111111111101011101000100;
        x_t[25] = 26'b11111111111101010010111110;
        x_t[26] = 26'b00000000000011011001010100;
        x_t[27] = 26'b00000000000011000011000110;
        x_t[28] = 26'b00000000000101001000111111;
        x_t[29] = 26'b11111111111101101101010011;
        x_t[30] = 26'b11111111111111100111101111;
        x_t[31] = 26'b00000000000010101110101101;
        x_t[32] = 26'b00000000001000000111000011;
        x_t[33] = 26'b00000000001000011110011010;
        x_t[34] = 26'b00000000000100111110001101;
        x_t[35] = 26'b00000000000100110100001001;
        x_t[36] = 26'b00000000000010101101010110;
        x_t[37] = 26'b00000000000000100100001001;
        x_t[38] = 26'b11111111111100110011100110;
        x_t[39] = 26'b00000000001100010010101011;
        x_t[40] = 26'b11111111111011000101110100;
        x_t[41] = 26'b11111111111110110100010101;
        x_t[42] = 26'b11111111111011011100111011;
        x_t[43] = 26'b00000000001110110111100100;
        x_t[44] = 26'b11111111111010010011101010;
        x_t[45] = 26'b00000000000001011011000011;
        x_t[46] = 26'b11111111111011010000111010;
        x_t[47] = 26'b11111111111110001111110111;
        x_t[48] = 26'b11111111111100111001100110;
        x_t[49] = 26'b00000000000011011111100000;
        x_t[50] = 26'b00000000000001111110111011;
        x_t[51] = 26'b11111111110111000101110000;
        x_t[52] = 26'b11111111110101010001100111;
        x_t[53] = 26'b11111111110001010010010011;
        x_t[54] = 26'b11111111101101001101100101;
        x_t[55] = 26'b11111111111000110100010001;
        x_t[56] = 26'b11111111111010111110001011;
        x_t[57] = 26'b11111111110111100110100010;
        x_t[58] = 26'b11111111101001100110101010;
        x_t[59] = 26'b11111111100011100101010000;
        x_t[60] = 26'b11111111101110111011110100;
        x_t[61] = 26'b11111111100000001001011001;
        x_t[62] = 26'b11111111001011011111001100;
        x_t[63] = 26'b11111111011111000000110000;
        
        h_t_prev[0] = 26'b00000000000100010001010101;
        h_t_prev[1] = 26'b00000000001001000001111100;
        h_t_prev[2] = 26'b00000000001010101110011000;
        h_t_prev[3] = 26'b00000000001110010110010100;
        h_t_prev[4] = 26'b00000000001110011101101110;
        h_t_prev[5] = 26'b00000000001000100000010010;
        h_t_prev[6] = 26'b00000000000101101000100011;
        h_t_prev[7] = 26'b00000000000000000010001111;
        h_t_prev[8] = 26'b00000000000011111110000101;
        h_t_prev[9] = 26'b00000000001100000001000100;
        h_t_prev[10] = 26'b00000000010010111111101010;
        h_t_prev[11] = 26'b00000000000111100101110100;
        h_t_prev[12] = 26'b00000000000110000011101000;
        h_t_prev[13] = 26'b00000000000101001111010110;
        h_t_prev[14] = 26'b11111111111101011001010110;
        h_t_prev[15] = 26'b00000000000011111110101100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 91 timeout!");
                $fdisplay(fd_cycles, "Test Vector  91: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  91: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 91");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 92
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000111000010111010;
        x_t[1] = 26'b00000000001101010100000001;
        x_t[2] = 26'b00000000001111010001101111;
        x_t[3] = 26'b00000000010010010001101100;
        x_t[4] = 26'b00000000010000101011001011;
        x_t[5] = 26'b00000000001001111001000011;
        x_t[6] = 26'b00000000000101101000100011;
        x_t[7] = 26'b00000000000000101010111101;
        x_t[8] = 26'b00000000001010101111010011;
        x_t[9] = 26'b00000000010010111010000011;
        x_t[10] = 26'b00000000011000110011011111;
        x_t[11] = 26'b00000000001001100000000111;
        x_t[12] = 26'b00000000001000010000000110;
        x_t[13] = 26'b00000000001010110001101100;
        x_t[14] = 26'b00000000000011010101000010;
        x_t[15] = 26'b00000000001010111110001101;
        x_t[16] = 26'b00000000001110010101110000;
        x_t[17] = 26'b00000000001101110100000011;
        x_t[18] = 26'b00000000001000000101100011;
        x_t[19] = 26'b00000000000011011010011111;
        x_t[20] = 26'b11111111111101010111111001;
        x_t[21] = 26'b00000000000101101100000011;
        x_t[22] = 26'b00000000000100010111011110;
        x_t[23] = 26'b11111111111111001101110100;
        x_t[24] = 26'b00000000000010100101111010;
        x_t[25] = 26'b00000000000010001001110001;
        x_t[26] = 26'b00000000000011001000011011;
        x_t[27] = 26'b00000000000001100100110001;
        x_t[28] = 26'b00000000000010110001110110;
        x_t[29] = 26'b00000000001001001001010111;
        x_t[30] = 26'b11111111111110011001101100;
        x_t[31] = 26'b00000000000001111001011110;
        x_t[32] = 26'b00000000001000101011011001;
        x_t[33] = 26'b00000000000111100110111010;
        x_t[34] = 26'b00000000000101010001010000;
        x_t[35] = 26'b00000000000101011011100111;
        x_t[36] = 26'b00000000000000110110000100;
        x_t[37] = 26'b11111111111010011100110001;
        x_t[38] = 26'b00000000000111001101001100;
        x_t[39] = 26'b00000000001100010010101011;
        x_t[40] = 26'b00000000001010011000000100;
        x_t[41] = 26'b11111111111101111100101100;
        x_t[42] = 26'b00000000001000011011000000;
        x_t[43] = 26'b00000000000011111001011001;
        x_t[44] = 26'b00000000000011000010001111;
        x_t[45] = 26'b00000000000001011011000011;
        x_t[46] = 26'b00000000000010011000110011;
        x_t[47] = 26'b00000000000100110001100111;
        x_t[48] = 26'b00000000000010010000101001;
        x_t[49] = 26'b00000000001001110111001111;
        x_t[50] = 26'b00000000001010010011000101;
        x_t[51] = 26'b11111111111111110101111111;
        x_t[52] = 26'b11111111111101100101101001;
        x_t[53] = 26'b11111111110111111001011010;
        x_t[54] = 26'b11111111110001101101001111;
        x_t[55] = 26'b11111111111100100101111101;
        x_t[56] = 26'b00000000000000000100101110;
        x_t[57] = 26'b00000000000000101010010100;
        x_t[58] = 26'b11111111110100100000100011;
        x_t[59] = 26'b11111111101110001100001100;
        x_t[60] = 26'b11111111110000100111001010;
        x_t[61] = 26'b11111111100110010110101011;
        x_t[62] = 26'b11111111010011010110001110;
        x_t[63] = 26'b11111111011111010010010111;
        
        h_t_prev[0] = 26'b00000000000111000010111010;
        h_t_prev[1] = 26'b00000000001101010100000001;
        h_t_prev[2] = 26'b00000000001111010001101111;
        h_t_prev[3] = 26'b00000000010010010001101100;
        h_t_prev[4] = 26'b00000000010000101011001011;
        h_t_prev[5] = 26'b00000000001001111001000011;
        h_t_prev[6] = 26'b00000000000101101000100011;
        h_t_prev[7] = 26'b00000000000000101010111101;
        h_t_prev[8] = 26'b00000000001010101111010011;
        h_t_prev[9] = 26'b00000000010010111010000011;
        h_t_prev[10] = 26'b00000000011000110011011111;
        h_t_prev[11] = 26'b00000000001001100000000111;
        h_t_prev[12] = 26'b00000000001000010000000110;
        h_t_prev[13] = 26'b00000000001010110001101100;
        h_t_prev[14] = 26'b00000000000011010101000010;
        h_t_prev[15] = 26'b00000000001010111110001101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 92 timeout!");
                $fdisplay(fd_cycles, "Test Vector  92: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  92: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 92");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 93
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001101001101100010;
        x_t[1] = 26'b00000000010010110100011010;
        x_t[2] = 26'b00000000010011100001101010;
        x_t[3] = 26'b00000000010101100110011000;
        x_t[4] = 26'b00000000010011100001000011;
        x_t[5] = 26'b00000000001101101101000111;
        x_t[6] = 26'b00000000001001001000100110;
        x_t[7] = 26'b00000000001010110110011011;
        x_t[8] = 26'b00000000010011011100010010;
        x_t[9] = 26'b00000000011010101111001010;
        x_t[10] = 26'b00000000100000110000010011;
        x_t[11] = 26'b00000000010011000011100111;
        x_t[12] = 26'b00000000001110011110000111;
        x_t[13] = 26'b00000000001110001011101111;
        x_t[14] = 26'b00000000001111110110100111;
        x_t[15] = 26'b00000000010110101110110110;
        x_t[16] = 26'b00000000011001011111100010;
        x_t[17] = 26'b00000000011000100110111100;
        x_t[18] = 26'b00000000010011100111011111;
        x_t[19] = 26'b00000000001111000101011000;
        x_t[20] = 26'b00000000000101111110100000;
        x_t[21] = 26'b00000000001001010100000111;
        x_t[22] = 26'b00000000001000001000101000;
        x_t[23] = 26'b00000000000011001101000100;
        x_t[24] = 26'b00000000000110000001001000;
        x_t[25] = 26'b00000000000101101001100010;
        x_t[26] = 26'b00000000000111010110110001;
        x_t[27] = 26'b00000000000111011110000110;
        x_t[28] = 26'b00000000000111100000001000;
        x_t[29] = 26'b00000000001100010001000001;
        x_t[30] = 26'b00000000000010100011000100;
        x_t[31] = 26'b00000000001000100011010011;
        x_t[32] = 26'b00000000001101110010011111;
        x_t[33] = 26'b00000000001101000110011101;
        x_t[34] = 26'b00000000001010010101001001;
        x_t[35] = 26'b00000000001011010010101000;
        x_t[36] = 26'b00000000001000010011001011;
        x_t[37] = 26'b00000000000000100100001001;
        x_t[38] = 26'b00000000001110011101000110;
        x_t[39] = 26'b00000000010000011011001111;
        x_t[40] = 26'b00000000010110111100011001;
        x_t[41] = 26'b00000000000001011011001111;
        x_t[42] = 26'b00000000001000110010101110;
        x_t[43] = 26'b11111111111100010110101001;
        x_t[44] = 26'b00000000001111100110100111;
        x_t[45] = 26'b00000000001100100010111100;
        x_t[46] = 26'b00000000001110000010110100;
        x_t[47] = 26'b00000000010001100001001110;
        x_t[48] = 26'b00000000001110011110000011;
        x_t[49] = 26'b00000000010101001010000010;
        x_t[50] = 26'b00000000010110001011010010;
        x_t[51] = 26'b00000000001111110101110111;
        x_t[52] = 26'b00000000001101100100110001;
        x_t[53] = 26'b00000000000111001101010001;
        x_t[54] = 26'b00000000000001011100000011;
        x_t[55] = 26'b00000000000111000111001111;
        x_t[56] = 26'b00000000001010010001110101;
        x_t[57] = 26'b00000000001100101001101011;
        x_t[58] = 26'b00000000000101001000110110;
        x_t[59] = 26'b11111111111110011110010001;
        x_t[60] = 26'b11111111111011011001001110;
        x_t[61] = 26'b11111111110101010110110011;
        x_t[62] = 26'b11111111100110111111110010;
        x_t[63] = 26'b11111111100111100010011100;
        
        h_t_prev[0] = 26'b00000000001101001101100010;
        h_t_prev[1] = 26'b00000000010010110100011010;
        h_t_prev[2] = 26'b00000000010011100001101010;
        h_t_prev[3] = 26'b00000000010101100110011000;
        h_t_prev[4] = 26'b00000000010011100001000011;
        h_t_prev[5] = 26'b00000000001101101101000111;
        h_t_prev[6] = 26'b00000000001001001000100110;
        h_t_prev[7] = 26'b00000000001010110110011011;
        h_t_prev[8] = 26'b00000000010011011100010010;
        h_t_prev[9] = 26'b00000000011010101111001010;
        h_t_prev[10] = 26'b00000000100000110000010011;
        h_t_prev[11] = 26'b00000000010011000011100111;
        h_t_prev[12] = 26'b00000000001110011110000111;
        h_t_prev[13] = 26'b00000000001110001011101111;
        h_t_prev[14] = 26'b00000000001111110110100111;
        h_t_prev[15] = 26'b00000000010110101110110110;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 93 timeout!");
                $fdisplay(fd_cycles, "Test Vector  93: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  93: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 93");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 94
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000010010001001001110;
        x_t[1] = 26'b00000000010111101101101001;
        x_t[2] = 26'b00000000010111011110001010;
        x_t[3] = 26'b00000000011000010100011010;
        x_t[4] = 26'b00000000010110111111010101;
        x_t[5] = 26'b00000000010000110100110100;
        x_t[6] = 26'b00000000001100001111110000;
        x_t[7] = 26'b00000000010000100100111000;
        x_t[8] = 26'b00000000010111111101000110;
        x_t[9] = 26'b00000000011100010011011000;
        x_t[10] = 26'b00000000100000011100101110;
        x_t[11] = 26'b00000000010110111000001110;
        x_t[12] = 26'b00000000010011111101010011;
        x_t[13] = 26'b00000000010011010010110101;
        x_t[14] = 26'b00000000010011110011101111;
        x_t[15] = 26'b00000000011000101000111001;
        x_t[16] = 26'b00000000011010101110110110;
        x_t[17] = 26'b00000000010111111111011101;
        x_t[18] = 26'b00000000010110010000001010;
        x_t[19] = 26'b00000000010101010000110010;
        x_t[20] = 26'b00000000001101000001000000;
        x_t[21] = 26'b00000000000110011000010000;
        x_t[22] = 26'b00000000000100110000110111;
        x_t[23] = 26'b11111111111110011111011010;
        x_t[24] = 26'b00000000000001000100011110;
        x_t[25] = 26'b00000000000000111111001011;
        x_t[26] = 26'b00000000000011101010001110;
        x_t[27] = 26'b00000000000001110100011111;
        x_t[28] = 26'b11111111111111000010100010;
        x_t[29] = 26'b00000000000110000001101101;
        x_t[30] = 26'b00000000000000000110111101;
        x_t[31] = 26'b00000000000011010010001100;
        x_t[32] = 26'b00000000001001001111101111;
        x_t[33] = 26'b00000000000111100110111010;
        x_t[34] = 26'b00000000000011110010000000;
        x_t[35] = 26'b00000000000100100000011010;
        x_t[36] = 26'b11111111111110101010111010;
        x_t[37] = 26'b11111111111001111100001010;
        x_t[38] = 26'b00000000001001000110001101;
        x_t[39] = 26'b00000000001010011101000101;
        x_t[40] = 26'b00000000001110011100111011;
        x_t[41] = 26'b11111111111011110001100110;
        x_t[42] = 26'b00000000000000101000111101;
        x_t[43] = 26'b11111111101111010100110100;
        x_t[44] = 26'b00000000000111001110010111;
        x_t[45] = 26'b00000000001001001010010010;
        x_t[46] = 26'b00000000001011001000010100;
        x_t[47] = 26'b00000000001101110010100000;
        x_t[48] = 26'b00000000001010000000001011;
        x_t[49] = 26'b00000000010000001110111110;
        x_t[50] = 26'b00000000001111010110001010;
        x_t[51] = 26'b00000000001110111011111010;
        x_t[52] = 26'b00000000001100111011110101;
        x_t[53] = 26'b00000000001000010000000101;
        x_t[54] = 26'b00000000000010001100000000;
        x_t[55] = 26'b00000000000110000010001011;
        x_t[56] = 26'b00000000000111010100110001;
        x_t[57] = 26'b00000000001011110110100001;
        x_t[58] = 26'b00000000001000111101000111;
        x_t[59] = 26'b00000000000100111000110010;
        x_t[60] = 26'b00000000000101001101111100;
        x_t[61] = 26'b00000000000010010010011111;
        x_t[62] = 26'b11111111111001000001110011;
        x_t[63] = 26'b11111111110001011100001001;
        
        h_t_prev[0] = 26'b00000000010010001001001110;
        h_t_prev[1] = 26'b00000000010111101101101001;
        h_t_prev[2] = 26'b00000000010111011110001010;
        h_t_prev[3] = 26'b00000000011000010100011010;
        h_t_prev[4] = 26'b00000000010110111111010101;
        h_t_prev[5] = 26'b00000000010000110100110100;
        h_t_prev[6] = 26'b00000000001100001111110000;
        h_t_prev[7] = 26'b00000000010000100100111000;
        h_t_prev[8] = 26'b00000000010111111101000110;
        h_t_prev[9] = 26'b00000000011100010011011000;
        h_t_prev[10] = 26'b00000000100000011100101110;
        h_t_prev[11] = 26'b00000000010110111000001110;
        h_t_prev[12] = 26'b00000000010011111101010011;
        h_t_prev[13] = 26'b00000000010011010010110101;
        h_t_prev[14] = 26'b00000000010011110011101111;
        h_t_prev[15] = 26'b00000000011000101000111001;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 94 timeout!");
                $fdisplay(fd_cycles, "Test Vector  94: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  94: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 94");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 95
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000001000111001010011;
        x_t[1] = 26'b00000000001101000000011100;
        x_t[2] = 26'b00000000001011000001110011;
        x_t[3] = 26'b00000000001010011010111100;
        x_t[4] = 26'b00000000001000011101110001;
        x_t[5] = 26'b00000000000001100100100001;
        x_t[6] = 26'b11111111111001111101101110;
        x_t[7] = 26'b00000000000111101010110110;
        x_t[8] = 26'b00000000001110100110110110;
        x_t[9] = 26'b00000000001111110001100110;
        x_t[10] = 26'b00000000010011100110110011;
        x_t[11] = 26'b00000000001010110001101001;
        x_t[12] = 26'b00000000001010000101001010;
        x_t[13] = 26'b00000000000110100001000111;
        x_t[14] = 26'b00000000001011111001011111;
        x_t[15] = 26'b00000000010000011000000000;
        x_t[16] = 26'b00000000010001101111110111;
        x_t[17] = 26'b00000000001111000011000000;
        x_t[18] = 26'b00000000001111101010011111;
        x_t[19] = 26'b00000000001111011011010110;
        x_t[20] = 26'b00000000001000010100101011;
        x_t[21] = 26'b11111111111101100100101001;
        x_t[22] = 26'b11111111111100110101001001;
        x_t[23] = 26'b11111111111000101100001010;
        x_t[24] = 26'b11111111111000111000110000;
        x_t[25] = 26'b11111111111001001101111010;
        x_t[26] = 26'b11111111111001000110010110;
        x_t[27] = 26'b11111111111000101110110010;
        x_t[28] = 26'b11111111111110000011100100;
        x_t[29] = 26'b11111111111110001110100100;
        x_t[30] = 26'b11111111111000110010101001;
        x_t[31] = 26'b11111111110111101001000000;
        x_t[32] = 26'b11111111111111010011101110;
        x_t[33] = 26'b11111111111011011101110011;
        x_t[34] = 26'b11111111110111100100110111;
        x_t[35] = 26'b11111111111001101101100101;
        x_t[36] = 26'b11111111110011011111010000;
        x_t[37] = 26'b11111111110100110110000000;
        x_t[38] = 26'b11111111111111111101010010;
        x_t[39] = 26'b11111111111111111000111110;
        x_t[40] = 26'b00000000000011100101010010;
        x_t[41] = 26'b11111111101011101100010101;
        x_t[42] = 26'b00000000000000010001001111;
        x_t[43] = 26'b00000000001010110000001111;
        x_t[44] = 26'b00000000000011101110111011;
        x_t[45] = 26'b00000000001101000001111001;
        x_t[46] = 26'b00000000001101101110000110;
        x_t[47] = 26'b00000000001110000110011001;
        x_t[48] = 26'b00000000001100000101100101;
        x_t[49] = 26'b00000000010010010000101101;
        x_t[50] = 26'b00000000010001101110001101;
        x_t[51] = 26'b00000000010011110001000000;
        x_t[52] = 26'b00000000010010010111101101;
        x_t[53] = 26'b00000000001111111010000000;
        x_t[54] = 26'b00000000001100010011001111;
        x_t[55] = 26'b00000000001100100000100000;
        x_t[56] = 26'b00000000001110010011101000;
        x_t[57] = 26'b00000000010011110110000101;
        x_t[58] = 26'b00000000010011010100000111;
        x_t[59] = 26'b00000000010010101100111110;
        x_t[60] = 26'b00000000001101100110101010;
        x_t[61] = 26'b00000000001111001110001011;
        x_t[62] = 26'b00000000000110101010101101;
        x_t[63] = 26'b11111111111111001100010010;
        
        h_t_prev[0] = 26'b00000000001000111001010011;
        h_t_prev[1] = 26'b00000000001101000000011100;
        h_t_prev[2] = 26'b00000000001011000001110011;
        h_t_prev[3] = 26'b00000000001010011010111100;
        h_t_prev[4] = 26'b00000000001000011101110001;
        h_t_prev[5] = 26'b00000000000001100100100001;
        h_t_prev[6] = 26'b11111111111001111101101110;
        h_t_prev[7] = 26'b00000000000111101010110110;
        h_t_prev[8] = 26'b00000000001110100110110110;
        h_t_prev[9] = 26'b00000000001111110001100110;
        h_t_prev[10] = 26'b00000000010011100110110011;
        h_t_prev[11] = 26'b00000000001010110001101001;
        h_t_prev[12] = 26'b00000000001010000101001010;
        h_t_prev[13] = 26'b00000000000110100001000111;
        h_t_prev[14] = 26'b00000000001011111001011111;
        h_t_prev[15] = 26'b00000000010000011000000000;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 95 timeout!");
                $fdisplay(fd_cycles, "Test Vector  95: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  95: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 95");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 96
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000100010001010101;
        x_t[1] = 26'b00000000000111110011101000;
        x_t[2] = 26'b00000000000101100100001100;
        x_t[3] = 26'b00000000000101010010001110;
        x_t[4] = 26'b00000000000011000110001110;
        x_t[5] = 26'b11111111111100101101111001;
        x_t[6] = 26'b11111111110110110110100101;
        x_t[7] = 26'b00000000000100011111010000;
        x_t[8] = 26'b00000000001001110001011010;
        x_t[9] = 26'b00000000001100111101001101;
        x_t[10] = 26'b00000000010001110001011000;
        x_t[11] = 26'b00000000001001100000000111;
        x_t[12] = 26'b00000000001000111110111011;
        x_t[13] = 26'b00000000000101001111010110;
        x_t[14] = 26'b00000000001010010000000001;
        x_t[15] = 26'b00000000001110110010010011;
        x_t[16] = 26'b00000000001111111000111001;
        x_t[17] = 26'b00000000010000100101101101;
        x_t[18] = 26'b00000000010001010011111001;
        x_t[19] = 26'b00000000010010001011000101;
        x_t[20] = 26'b00000000001011011100111001;
        x_t[21] = 26'b11111111111011101011000101;
        x_t[22] = 26'b11111111111001110110110000;
        x_t[23] = 26'b11111111110110001001101111;
        x_t[24] = 26'b11111111110111100011100000;
        x_t[25] = 26'b11111111110111110110111001;
        x_t[26] = 26'b11111111110101101010101100;
        x_t[27] = 26'b11111111110110000001110110;
        x_t[28] = 26'b11111111111101010001001100;
        x_t[29] = 26'b11111111111110011111001101;
        x_t[30] = 26'b11111111111000100011000010;
        x_t[31] = 26'b11111111110110110011110001;
        x_t[32] = 26'b11111111111100110000001011;
        x_t[33] = 26'b11111111111010000001010010;
        x_t[34] = 26'b11111111110101011111011111;
        x_t[35] = 26'b11111111110110101000001101;
        x_t[36] = 26'b11111111110011001011011000;
        x_t[37] = 26'b11111111110011100100011110;
        x_t[38] = 26'b11111111111111010100111101;
        x_t[39] = 26'b11111111111011010011000000;
        x_t[40] = 26'b00000000000011111011000001;
        x_t[41] = 26'b11111111100111010110001001;
        x_t[42] = 26'b00000000000011111110011010;
        x_t[43] = 26'b00000000001110110111100100;
        x_t[44] = 26'b11111111111110011111110010;
        x_t[45] = 26'b00000000010100010010001011;
        x_t[46] = 26'b00000000001000110111010000;
        x_t[47] = 26'b00000000001100100010111011;
        x_t[48] = 26'b00000000001010111001010110;
        x_t[49] = 26'b00000000010010110101110001;
        x_t[50] = 26'b00000000010011110011001111;
        x_t[51] = 26'b00000000010110011110110111;
        x_t[52] = 26'b00000000010100100110111100;
        x_t[53] = 26'b00000000010011101110111110;
        x_t[54] = 26'b00000000010011000010101110;
        x_t[55] = 26'b00000000001110101010100111;
        x_t[56] = 26'b00000000001111000111001100;
        x_t[57] = 26'b00000000010111110101110111;
        x_t[58] = 26'b00000000010110110110111011;
        x_t[59] = 26'b00000000010111111000100010;
        x_t[60] = 26'b00000000010100010100000010;
        x_t[61] = 26'b00000000011001100100010100;
        x_t[62] = 26'b00000000001111101011101101;
        x_t[63] = 26'b00000000001100101010110100;
        
        h_t_prev[0] = 26'b00000000000100010001010101;
        h_t_prev[1] = 26'b00000000000111110011101000;
        h_t_prev[2] = 26'b00000000000101100100001100;
        h_t_prev[3] = 26'b00000000000101010010001110;
        h_t_prev[4] = 26'b00000000000011000110001110;
        h_t_prev[5] = 26'b11111111111100101101111001;
        h_t_prev[6] = 26'b11111111110110110110100101;
        h_t_prev[7] = 26'b00000000000100011111010000;
        h_t_prev[8] = 26'b00000000001001110001011010;
        h_t_prev[9] = 26'b00000000001100111101001101;
        h_t_prev[10] = 26'b00000000010001110001011000;
        h_t_prev[11] = 26'b00000000001001100000000111;
        h_t_prev[12] = 26'b00000000001000111110111011;
        h_t_prev[13] = 26'b00000000000101001111010110;
        h_t_prev[14] = 26'b00000000001010010000000001;
        h_t_prev[15] = 26'b00000000001110110010010011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 96 timeout!");
                $fdisplay(fd_cycles, "Test Vector  96: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  96: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 96");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 97
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111111100010000010101;
        x_t[1] = 26'b11111111111100011111010001;
        x_t[2] = 26'b11111111110111100110101111;
        x_t[3] = 26'b11111111111010011010001000;
        x_t[4] = 26'b11111111111011110101011100;
        x_t[5] = 26'b11111111111001111100011000;
        x_t[6] = 26'b11111111111100101011111111;
        x_t[7] = 26'b11111111111111101101111000;
        x_t[8] = 26'b11111111111001000000101100;
        x_t[9] = 26'b11111111110101011101110111;
        x_t[10] = 26'b11111111110110110111001111;
        x_t[11] = 26'b11111111110110011001000110;
        x_t[12] = 26'b11111111111011110100000100;
        x_t[13] = 26'b00000000000010101011110011;
        x_t[14] = 26'b11111111111001000111001000;
        x_t[15] = 26'b11111111111001011111011011;
        x_t[16] = 26'b11111111110111000110101101;
        x_t[17] = 26'b11111111110101110000010101;
        x_t[18] = 26'b11111111111010010000000010;
        x_t[19] = 26'b11111111111000011011100011;
        x_t[20] = 26'b00000000000010110110010010;
        x_t[21] = 26'b00000000000110000010001001;
        x_t[22] = 26'b00000000000101111101000001;
        x_t[23] = 26'b00000000000011100100010001;
        x_t[24] = 26'b00000000000011101110111110;
        x_t[25] = 26'b00000000000011010100010111;
        x_t[26] = 26'b00000000000001100011000010;
        x_t[27] = 26'b11111111111101101001001110;
        x_t[28] = 26'b11111111111011101100011011;
        x_t[29] = 26'b00000000000000110100111101;
        x_t[30] = 26'b00000000000100000000101111;
        x_t[31] = 26'b11111111111110010010110101;
        x_t[32] = 26'b00000000000001000000110000;
        x_t[33] = 26'b11111111111101001100110100;
        x_t[34] = 26'b11111111111100111011110011;
        x_t[35] = 26'b11111111111110000001111010;
        x_t[36] = 26'b11111111111100001011111000;
        x_t[37] = 26'b11111111111100101111100010;
        x_t[38] = 26'b11111111111111111101010010;
        x_t[39] = 26'b00000000001001000100111001;
        x_t[40] = 26'b11111111111111001010101011;
        x_t[41] = 26'b00000000011000011101100110;
        x_t[42] = 26'b11111111111100111011110011;
        x_t[43] = 26'b00000000001000000000101101;
        x_t[44] = 26'b11111111111000001101100110;
        x_t[45] = 26'b00000000001010100111001000;
        x_t[46] = 26'b11111111110011110100010011;
        x_t[47] = 26'b11111111111001010001100100;
        x_t[48] = 26'b11111111111001100111111100;
        x_t[49] = 26'b11111111111010100000111101;
        x_t[50] = 26'b11111111111001010111110010;
        x_t[51] = 26'b11111111111011010100001101;
        x_t[52] = 26'b11111111111011101010110111;
        x_t[53] = 26'b11111111111111001101000101;
        x_t[54] = 26'b00000000000010111011111100;
        x_t[55] = 26'b11111111110101000010100101;
        x_t[56] = 26'b11111111111010011011110011;
        x_t[57] = 26'b11111111111100001000011011;
        x_t[58] = 26'b11111111111100111101011011;
        x_t[59] = 26'b11111111111100011111111101;
        x_t[60] = 26'b11111111111100100101111001;
        x_t[61] = 26'b11111111111010000000110001;
        x_t[62] = 26'b11111111111010011010100100;
        x_t[63] = 26'b00000000000000110101111001;
        
        h_t_prev[0] = 26'b11111111111100010000010101;
        h_t_prev[1] = 26'b11111111111100011111010001;
        h_t_prev[2] = 26'b11111111110111100110101111;
        h_t_prev[3] = 26'b11111111111010011010001000;
        h_t_prev[4] = 26'b11111111111011110101011100;
        h_t_prev[5] = 26'b11111111111001111100011000;
        h_t_prev[6] = 26'b11111111111100101011111111;
        h_t_prev[7] = 26'b11111111111111101101111000;
        h_t_prev[8] = 26'b11111111111001000000101100;
        h_t_prev[9] = 26'b11111111110101011101110111;
        h_t_prev[10] = 26'b11111111110110110111001111;
        h_t_prev[11] = 26'b11111111110110011001000110;
        h_t_prev[12] = 26'b11111111111011110100000100;
        h_t_prev[13] = 26'b00000000000010101011110011;
        h_t_prev[14] = 26'b11111111111001000111001000;
        h_t_prev[15] = 26'b11111111111001011111011011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 97 timeout!");
                $fdisplay(fd_cycles, "Test Vector  97: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  97: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 97");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 98
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b00000000000000010000110101;
        x_t[1] = 26'b11111111111111110110100111;
        x_t[2] = 26'b11111111111010101000111101;
        x_t[3] = 26'b11111111111110010101100000;
        x_t[4] = 26'b11111111111110000010111001;
        x_t[5] = 26'b11111111111011101011010101;
        x_t[6] = 26'b11111111111101000100111000;
        x_t[7] = 26'b00000000000001101000000010;
        x_t[8] = 26'b11111111111001111110100101;
        x_t[9] = 26'b11111111110111000010000101;
        x_t[10] = 26'b11111111111001100111010111;
        x_t[11] = 26'b11111111111001100100111100;
        x_t[12] = 26'b11111111111100111010010100;
        x_t[13] = 26'b00000000000101101010100110;
        x_t[14] = 26'b11111111111001011100001110;
        x_t[15] = 26'b11111111111000001110000011;
        x_t[16] = 26'b11111111110110110010111000;
        x_t[17] = 26'b11111111110110111111010010;
        x_t[18] = 26'b11111111111010100101000111;
        x_t[19] = 26'b11111111110111011001101001;
        x_t[20] = 26'b00000000000001010010001011;
        x_t[21] = 26'b00000000000110011000010000;
        x_t[22] = 26'b00000000000101100011101000;
        x_t[23] = 26'b00000000000011001101000100;
        x_t[24] = 26'b00000000000011111011001010;
        x_t[25] = 26'b00000000000011101101001110;
        x_t[26] = 26'b00000000000000110000010110;
        x_t[27] = 26'b11111111111110001000101010;
        x_t[28] = 26'b11111111111010101101011101;
        x_t[29] = 26'b00000000000000110100111101;
        x_t[30] = 26'b00000000000100000000101111;
        x_t[31] = 26'b11111111111111001000000011;
        x_t[32] = 26'b00000000000001000000110000;
        x_t[33] = 26'b11111111111100100111110011;
        x_t[34] = 26'b11111111111100010101101100;
        x_t[35] = 26'b11111111111100011111001110;
        x_t[36] = 26'b11111111111011010000001111;
        x_t[37] = 26'b11111111111010001100011101;
        x_t[38] = 26'b11111111111111010100111101;
        x_t[39] = 26'b00000000000100011110111011;
        x_t[40] = 26'b11111111111011011011100011;
        x_t[41] = 26'b00000000000010101110101100;
        x_t[42] = 26'b11111111111001100110010110;
        x_t[43] = 26'b00000000000100100101010001;
        x_t[44] = 26'b11111111110100000001011110;
        x_t[45] = 26'b00000000000100110011101101;
        x_t[46] = 26'b11111111110000100101000100;
        x_t[47] = 26'b11111111110101001110111101;
        x_t[48] = 26'b11111111110101011101001000;
        x_t[49] = 26'b11111111110111000010100011;
        x_t[50] = 26'b11111111110110101100101110;
        x_t[51] = 26'b11111111110111111111101101;
        x_t[52] = 26'b11111111111000001001110001;
        x_t[53] = 26'b11111111111001111111000010;
        x_t[54] = 26'b11111111111011011100100000;
        x_t[55] = 26'b11111111101111101001010100;
        x_t[56] = 26'b11111111110101000100000100;
        x_t[57] = 26'b11111111110111100110100010;
        x_t[58] = 26'b11111111111001101100000011;
        x_t[59] = 26'b11111111111010000010000100;
        x_t[60] = 26'b11111111111000110000100010;
        x_t[61] = 26'b11111111110111111100010101;
        x_t[62] = 26'b11111111111001111100111110;
        x_t[63] = 26'b11111111111110101001000101;
        
        h_t_prev[0] = 26'b00000000000000010000110101;
        h_t_prev[1] = 26'b11111111111111110110100111;
        h_t_prev[2] = 26'b11111111111010101000111101;
        h_t_prev[3] = 26'b11111111111110010101100000;
        h_t_prev[4] = 26'b11111111111110000010111001;
        h_t_prev[5] = 26'b11111111111011101011010101;
        h_t_prev[6] = 26'b11111111111101000100111000;
        h_t_prev[7] = 26'b00000000000001101000000010;
        h_t_prev[8] = 26'b11111111111001111110100101;
        h_t_prev[9] = 26'b11111111110111000010000101;
        h_t_prev[10] = 26'b11111111111001100111010111;
        h_t_prev[11] = 26'b11111111111001100100111100;
        h_t_prev[12] = 26'b11111111111100111010010100;
        h_t_prev[13] = 26'b00000000000101101010100110;
        h_t_prev[14] = 26'b11111111111001011100001110;
        h_t_prev[15] = 26'b11111111111000001110000011;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 98 timeout!");
                $fdisplay(fd_cycles, "Test Vector  98: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  98: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 98");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 99
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111111011101000110111;
        x_t[1] = 26'b11111111111010010110001110;
        x_t[2] = 26'b11111111110101110010001100;
        x_t[3] = 26'b11111111111001110011011101;
        x_t[4] = 26'b11111111111001010011110010;
        x_t[5] = 26'b11111111110110110100101100;
        x_t[6] = 26'b11111111110110110110100101;
        x_t[7] = 26'b11111111111010101000001001;
        x_t[8] = 26'b11111111110010100100000111;
        x_t[9] = 26'b11111111110000001001000111;
        x_t[10] = 26'b11111111110010111000110101;
        x_t[11] = 26'b11111111110001111011101111;
        x_t[12] = 26'b11111111110011110000111111;
        x_t[13] = 26'b11111111111000111000111000;
        x_t[14] = 26'b11111111110010110110010110;
        x_t[15] = 26'b11111111101111101000110101;
        x_t[16] = 26'b11111111101110000111101101;
        x_t[17] = 26'b11111111101111100101100010;
        x_t[18] = 26'b11111111110001101011110110;
        x_t[19] = 26'b11111111101100110000101010;
        x_t[20] = 26'b11111111110010110100001001;
        x_t[21] = 26'b00000000000100101001101111;
        x_t[22] = 26'b00000000000011011000000000;
        x_t[23] = 26'b00000000000001011001000010;
        x_t[24] = 26'b00000000000000101100000111;
        x_t[25] = 26'b00000000000000011001111000;
        x_t[26] = 26'b11111111111100110010111001;
        x_t[27] = 26'b11111111111010101100100100;
        x_t[28] = 26'b11111111110111110000100001;
        x_t[29] = 26'b11111111111101101101010011;
        x_t[30] = 26'b00000000000000010110100101;
        x_t[31] = 26'b11111111111010101100001011;
        x_t[32] = 26'b11111111111011010101010100;
        x_t[33] = 26'b11111111110111011010110000;
        x_t[34] = 26'b11111111111000001010111101;
        x_t[35] = 26'b11111111111000011110101000;
        x_t[36] = 26'b11111111110101111110010011;
        x_t[37] = 26'b11111111110101110111001111;
        x_t[38] = 26'b11111111111100001011010000;
        x_t[39] = 26'b11111111111001000000000001;
        x_t[40] = 26'b11111111111000010111111010;
        x_t[41] = 26'b11111111110001010101111110;
        x_t[42] = 26'b11111111110111000000010101;
        x_t[43] = 26'b11111111111010111110111000;
        x_t[44] = 26'b11111111110000111000011001;
        x_t[45] = 26'b11111111110000011111101110;
        x_t[46] = 26'b11111111101100101100011010;
        x_t[47] = 26'b11111111101110000101011011;
        x_t[48] = 26'b11111111101100110100011011;
        x_t[49] = 26'b11111111101100100111010110;
        x_t[50] = 26'b11111111101100010011100011;
        x_t[51] = 26'b11111111101100001110010010;
        x_t[52] = 26'b11111111101010101110010110;
        x_t[53] = 26'b11111111101001101000010111;
        x_t[54] = 26'b11111111100110110110000100;
        x_t[55] = 26'b11111111101001011100010001;
        x_t[56] = 26'b11111111101101000000011110;
        x_t[57] = 26'b11111111101110000000101010;
        x_t[58] = 26'b11111111101101111101110100;
        x_t[59] = 26'b11111111101100101101011101;
        x_t[60] = 26'b11111111110011101110100001;
        x_t[61] = 26'b11111111110001101111000011;
        x_t[62] = 26'b11111111110100011001111001;
        x_t[63] = 26'b11111111111000000010100111;
        
        h_t_prev[0] = 26'b11111111111011101000110111;
        h_t_prev[1] = 26'b11111111111010010110001110;
        h_t_prev[2] = 26'b11111111110101110010001100;
        h_t_prev[3] = 26'b11111111111001110011011101;
        h_t_prev[4] = 26'b11111111111001010011110010;
        h_t_prev[5] = 26'b11111111110110110100101100;
        h_t_prev[6] = 26'b11111111110110110110100101;
        h_t_prev[7] = 26'b11111111111010101000001001;
        h_t_prev[8] = 26'b11111111110010100100000111;
        h_t_prev[9] = 26'b11111111110000001001000111;
        h_t_prev[10] = 26'b11111111110010111000110101;
        h_t_prev[11] = 26'b11111111110001111011101111;
        h_t_prev[12] = 26'b11111111110011110000111111;
        h_t_prev[13] = 26'b11111111111000111000111000;
        h_t_prev[14] = 26'b11111111110010110110010110;
        h_t_prev[15] = 26'b11111111101111101000110101;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 99 timeout!");
                $fdisplay(fd_cycles, "Test Vector  99: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector  99: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 99");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Test Vector 100
    if (!test_timeout) begin
        test_start_cycle = cycle_count;
        
        // Load input data
        x_t[0] = 26'b11111111111011101000110111;
        x_t[1] = 26'b11111111111001000111111010;
        x_t[2] = 26'b11111111110010101111111101;
        x_t[3] = 26'b11111111110111011000110001;
        x_t[4] = 26'b11111111110111011010100010;
        x_t[5] = 26'b11111111110100101111100100;
        x_t[6] = 26'b11111111110110000100110010;
        x_t[7] = 26'b11111111111100100010010010;
        x_t[8] = 26'b11111111101111010101110100;
        x_t[9] = 26'b11111111101100000100100010;
        x_t[10] = 26'b11111111101101011000100101;
        x_t[11] = 26'b11111111101100001100110101;
        x_t[12] = 26'b11111111101100011100101111;
        x_t[13] = 26'b11111111110001001110010000;
        x_t[14] = 26'b11111111110011100000100010;
        x_t[15] = 26'b11111111101101011010011100;
        x_t[16] = 26'b11111111101001001010011110;
        x_t[17] = 26'b11111111101001011010101111;
        x_t[18] = 26'b11111111101011110000010110;
        x_t[19] = 26'b11111111100100100001011101;
        x_t[20] = 26'b11111111101001000010011101;
        x_t[21] = 26'b00000000001000100111111010;
        x_t[22] = 26'b00000000001001001000000110;
        x_t[23] = 26'b00000000000110010010010010;
        x_t[24] = 26'b00000000000101101000110001;
        x_t[25] = 26'b00000000000100110111110100;
        x_t[26] = 26'b00000000000011001000011011;
        x_t[27] = 26'b00000000000000100101111000;
        x_t[28] = 26'b11111111111100101011011001;
        x_t[29] = 26'b00000000000100101110100001;
        x_t[30] = 26'b00000000000100010000010110;
        x_t[31] = 26'b11111111111110110110010100;
        x_t[32] = 26'b11111111111111000001100011;
        x_t[33] = 26'b11111111111101011111010100;
        x_t[34] = 26'b11111111111110101110000111;
        x_t[35] = 26'b11111111111110101001011001;
        x_t[36] = 26'b11111111111101101111010010;
        x_t[37] = 26'b11111111111100111111110110;
        x_t[38] = 26'b00000000000010110010110100;
        x_t[39] = 26'b11111111111110100000110001;
        x_t[40] = 26'b00000000000001100010110110;
        x_t[41] = 26'b11111111111100001101011011;
        x_t[42] = 26'b00000000000001110000000111;
        x_t[43] = 26'b11111111101101010001001010;
        x_t[44] = 26'b11111111110100101110001010;
        x_t[45] = 26'b11111111100001111111001010;
        x_t[46] = 26'b11111111101110101000101111;
        x_t[47] = 26'b11111111101101110001100010;
        x_t[48] = 26'b11111111101011010101001000;
        x_t[49] = 26'b11111111101001001000111100;
        x_t[50] = 26'b11111111101000001001011110;
        x_t[51] = 26'b11111111100111011001001100;
        x_t[52] = 26'b11111111100111001101010000;
        x_t[53] = 26'b11111111100100000100000011;
        x_t[54] = 26'b11111111100001001110011111;
        x_t[55] = 26'b11111111100111100011011011;
        x_t[56] = 26'b11111111101000111110101011;
        x_t[57] = 26'b11111111101010000000110111;
        x_t[58] = 26'b11111111101001010101001101;
        x_t[59] = 26'b11111111100111110001101011;
        x_t[60] = 26'b11111111101110111011110100;
        x_t[61] = 26'b11111111101100000010110111;
        x_t[62] = 26'b11111111101110110110110100;
        x_t[63] = 26'b11111111110101010010100101;
        
        h_t_prev[0] = 26'b11111111111011101000110111;
        h_t_prev[1] = 26'b11111111111001000111111010;
        h_t_prev[2] = 26'b11111111110010101111111101;
        h_t_prev[3] = 26'b11111111110111011000110001;
        h_t_prev[4] = 26'b11111111110111011010100010;
        h_t_prev[5] = 26'b11111111110100101111100100;
        h_t_prev[6] = 26'b11111111110110000100110010;
        h_t_prev[7] = 26'b11111111111100100010010010;
        h_t_prev[8] = 26'b11111111101111010101110100;
        h_t_prev[9] = 26'b11111111101100000100100010;
        h_t_prev[10] = 26'b11111111101101011000100101;
        h_t_prev[11] = 26'b11111111101100001100110101;
        h_t_prev[12] = 26'b11111111101100011100101111;
        h_t_prev[13] = 26'b11111111110001001110010000;
        h_t_prev[14] = 26'b11111111110011100000100010;
        h_t_prev[15] = 26'b11111111101101011010011100;
        
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;
        
        // Wait for completion with timeout
        fork
            begin
                wait(done);
                test_cycles = cycle_count - test_start_cycle;
            end
            begin
                repeat(200000) @(posedge clk);
                $display("ERROR: Test 100 timeout!");
                $fdisplay(fd_cycles, "Test Vector 100: TIMEOUT");
                test_cycles = -1;
                test_timeout = 1;
            end
        join_any
        disable fork;
        
        if (test_cycles > 0) begin
            repeat(5) @(posedge clk); // Extra cycles for stability
            total_cycles = total_cycles + test_cycles;
            $fdisplay(fd_cycles, "Test Vector 100: %0d cycles (%.2f us @ 100MHz)", test_cycles, test_cycles * 0.01);
            
            // Write outputs
            $fdisplay(fd_output, "%026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b %026b", h_t[0], h_t[1], h_t[2], h_t[3], h_t[4], h_t[5], h_t[6], h_t[7], h_t[8], h_t[9], h_t[10], h_t[11], h_t[12], h_t[13], h_t[14], h_t[15]);
        end else begin
            $display("Stopping simulation due to timeout on test 100");
        end
        
        repeat(5) @(posedge clk); // Wait between tests
    end

    // Write summary to cycles file
    $fdisplay(fd_cycles, "");
    $fdisplay(fd_cycles, "==========================================================");
    $fdisplay(fd_cycles, "SUMMARY");
    $fdisplay(fd_cycles, "==========================================================");
    $fdisplay(fd_cycles, "Total Test Vectors: %0d", 100);
    $fdisplay(fd_cycles, "Total Cycles:       %0d", total_cycles);
    $fdisplay(fd_cycles, "Average Cycles:     %.2f", real'(total_cycles) / 100);
    $fdisplay(fd_cycles, "Total Time:         %.2f us @ 100MHz", total_cycles * 0.01);
    $fdisplay(fd_cycles, "Average Time:       %.2f us @ 100MHz", (total_cycles * 0.01) / 100);
    $fdisplay(fd_cycles, "Throughput:         %.2f computations/ms @ 100MHz", 100000.0 / (real'(total_cycles) / 100));
    $fdisplay(fd_cycles, "==========================================================");
    
    $fclose(fd_output);
    $fclose(fd_cycles);
    
    $display("");
    $display("==========================================================");
    $display("Simulation Complete");
    $display("==========================================================");
    $display("Test Vectors:   %0d", 100);
    $display("Total Cycles:   %0d", total_cycles);
    $display("Average Cycles: %.2f", real'(total_cycles) / 100);
    $display("==========================================================");
    $display("Output file:    output_d64_h16_dw26_fb16_np16.txt");
    $display("Cycles file:    cycles_d64_h16_dw26_fb16_np16.txt");
    $display("==========================================================");
    
    $finish;
end

endmodule