`timescale 1ns / 1ps

module gru_tb;

// Parameters
parameter int INT_WIDTH  = 4;
parameter int FRAC_WIDTH = 5;
parameter int WIDTH      = INT_WIDTH + FRAC_WIDTH;
parameter real CLK_PERIOD = 10.0;

// Clock and reset
logic clk;
logic reset;

// Inputs
logic signed [WIDTH-1:0] x_0 = 0;
logic signed [WIDTH-1:0] x_1 = 0;
logic signed [WIDTH-1:0] x_2 = 0;
logic signed [WIDTH-1:0] x_3 = 0;
logic signed [WIDTH-1:0] x_4 = 0;
logic signed [WIDTH-1:0] x_5 = 0;
logic signed [WIDTH-1:0] x_6 = 0;
logic signed [WIDTH-1:0] x_7 = 0;
logic signed [WIDTH-1:0] x_8 = 0;
logic signed [WIDTH-1:0] x_9 = 0;
logic signed [WIDTH-1:0] x_10 = 0;
logic signed [WIDTH-1:0] x_11 = 0;
logic signed [WIDTH-1:0] x_12 = 0;
logic signed [WIDTH-1:0] x_13 = 0;
logic signed [WIDTH-1:0] x_14 = 0;
logic signed [WIDTH-1:0] x_15 = 0;
logic signed [WIDTH-1:0] x_16 = 0;
logic signed [WIDTH-1:0] x_17 = 0;
logic signed [WIDTH-1:0] x_18 = 0;
logic signed [WIDTH-1:0] x_19 = 0;
logic signed [WIDTH-1:0] x_20 = 0;
logic signed [WIDTH-1:0] x_21 = 0;
logic signed [WIDTH-1:0] x_22 = 0;
logic signed [WIDTH-1:0] x_23 = 0;
logic signed [WIDTH-1:0] x_24 = 0;
logic signed [WIDTH-1:0] x_25 = 0;
logic signed [WIDTH-1:0] x_26 = 0;
logic signed [WIDTH-1:0] x_27 = 0;
logic signed [WIDTH-1:0] x_28 = 0;
logic signed [WIDTH-1:0] x_29 = 0;
logic signed [WIDTH-1:0] x_30 = 0;
logic signed [WIDTH-1:0] x_31 = 0;
logic signed [WIDTH-1:0] x_32 = 0;
logic signed [WIDTH-1:0] x_33 = 0;
logic signed [WIDTH-1:0] x_34 = 0;
logic signed [WIDTH-1:0] x_35 = 0;
logic signed [WIDTH-1:0] x_36 = 0;
logic signed [WIDTH-1:0] x_37 = 0;
logic signed [WIDTH-1:0] x_38 = 0;
logic signed [WIDTH-1:0] x_39 = 0;
logic signed [WIDTH-1:0] x_40 = 0;
logic signed [WIDTH-1:0] x_41 = 0;
logic signed [WIDTH-1:0] x_42 = 0;
logic signed [WIDTH-1:0] x_43 = 0;
logic signed [WIDTH-1:0] x_44 = 0;
logic signed [WIDTH-1:0] x_45 = 0;
logic signed [WIDTH-1:0] x_46 = 0;
logic signed [WIDTH-1:0] x_47 = 0;
logic signed [WIDTH-1:0] x_48 = 0;
logic signed [WIDTH-1:0] x_49 = 0;
logic signed [WIDTH-1:0] x_50 = 0;
logic signed [WIDTH-1:0] x_51 = 0;
logic signed [WIDTH-1:0] x_52 = 0;
logic signed [WIDTH-1:0] x_53 = 0;
logic signed [WIDTH-1:0] x_54 = 0;
logic signed [WIDTH-1:0] x_55 = 0;
logic signed [WIDTH-1:0] x_56 = 0;
logic signed [WIDTH-1:0] x_57 = 0;
logic signed [WIDTH-1:0] x_58 = 0;
logic signed [WIDTH-1:0] x_59 = 0;
logic signed [WIDTH-1:0] x_60 = 0;
logic signed [WIDTH-1:0] x_61 = 0;
logic signed [WIDTH-1:0] x_62 = 0;
logic signed [WIDTH-1:0] x_63 = 0;

logic signed [WIDTH-1:0] h_0 = 0;
logic signed [WIDTH-1:0] h_1 = 0;
logic signed [WIDTH-1:0] h_2 = 0;
logic signed [WIDTH-1:0] h_3 = 0;

// Input weights (h×d for each gate)
logic signed [WIDTH-1:0] w_ir_0_0 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_1 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_0_2 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_3 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_4 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_5 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_0_6 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_7 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_8 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_0_9 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_10 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_0_11 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_12 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_0_13 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_14 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_15 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_0_16 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_17 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_0_18 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_19 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_0_20 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_21 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_22 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_23 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_24 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_0_25 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_26 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_27 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_28 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_0_29 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_0_30 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_31 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_32 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_33 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_34 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_35 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_0_36 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_0_37 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_38 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_39 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_40 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_0_41 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_0_42 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_43 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_44 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_45 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_0_46 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_0_47 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_0_48 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_0_49 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_50 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_0_51 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_0_52 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_0_53 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_54 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_0_55 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_56 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_0_57 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_58 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_0_59 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_60 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_0_61 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_0_62 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_0_63 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_1_0 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_1 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_2 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_1_3 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_1_4 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_5 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_6 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_7 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_8 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_9 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_10 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_11 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_12 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_13 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_1_14 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_1_15 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_16 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_17 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_18 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_19 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_20 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_21 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_22 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_23 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_24 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_25 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_1_26 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_1_27 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_1_28 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_1_29 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_30 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_31 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_32 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_33 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_34 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_35 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_36 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_37 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_38 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_39 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_1_40 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_41 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_42 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_43 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_44 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_1_45 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_46 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_1_47 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_48 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_49 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_1_50 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_1_51 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_1_52 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_53 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_54 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_55 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_1_56 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_57 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_1_58 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_1_59 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_1_60 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_1_61 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_62 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_1_63 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_2_0 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_2_1 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_2 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_2_3 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_2_4 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_5 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_6 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_7 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_2_8 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_9 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_10 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_11 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_2_12 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_13 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_14 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_15 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_2_16 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_2_17 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_2_18 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_19 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_20 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_21 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_22 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_23 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_2_24 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_2_25 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_26 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_27 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_2_28 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_29 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_2_30 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_2_31 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_2_32 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_33 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_2_34 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_2_35 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_36 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_37 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_38 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_39 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_40 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_41 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_2_42 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_2_43 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_44 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_45 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_46 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_47 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_48 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_49 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_50 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_2_51 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_2_52 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_2_53 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_54 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_2_55 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_56 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_57 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_2_58 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_2_59 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_2_60 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_2_61 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_2_62 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_2_63 = 'b000001001;
logic signed [WIDTH-1:0] w_ir_3_0 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_1 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_3_2 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_3 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_3_4 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_3_5 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_6 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_7 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_8 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_9 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_3_10 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_11 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_12 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_13 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_14 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_15 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_16 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_17 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_18 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_19 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_20 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_21 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_22 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_3_23 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_24 = 'b000000111;
logic signed [WIDTH-1:0] w_ir_3_25 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_26 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_27 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_28 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_29 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_30 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_31 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_3_32 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_33 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_3_34 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_3_35 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_36 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_37 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_3_38 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_3_39 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_40 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_3_41 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_3_42 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_3_43 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_3_44 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_45 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_46 = 'b000000110;
logic signed [WIDTH-1:0] w_ir_3_47 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_48 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_49 = 'b111111111;
logic signed [WIDTH-1:0] w_ir_3_50 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_51 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_52 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_53 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_54 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_3_55 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_3_56 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_57 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_3_58 = 'b111111100;
logic signed [WIDTH-1:0] w_ir_3_59 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_60 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_61 = 'b111111101;
logic signed [WIDTH-1:0] w_ir_3_62 = 'b111111010;
logic signed [WIDTH-1:0] w_ir_3_63 = 'b111111110;

logic signed [WIDTH-1:0] w_iz_0_0 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_1 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_2 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_3 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_4 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_5 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_0_6 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_0_7 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_0_8 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_0_9 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_10 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_0_11 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_12 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_13 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_0_14 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_0_15 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_16 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_0_17 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_18 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_0_19 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_0_20 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_21 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_0_22 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_0_23 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_0_24 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_0_25 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_0_26 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_27 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_0_28 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_0_29 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_30 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_0_31 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_0_32 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_0_33 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_0_34 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_0_35 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_0_36 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_0_37 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_0_38 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_39 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_0_40 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_0_41 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_0_42 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_43 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_44 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_0_45 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_46 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_47 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_48 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_0_49 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_0_50 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_0_51 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_0_52 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_0_53 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_54 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_0_55 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_0_56 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_0_57 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_0_58 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_0_59 = 'b000001110;
logic signed [WIDTH-1:0] w_iz_0_60 = 'b000001010;
logic signed [WIDTH-1:0] w_iz_0_61 = 'b000001011;
logic signed [WIDTH-1:0] w_iz_0_62 = 'b000001101;
logic signed [WIDTH-1:0] w_iz_0_63 = 'b000001100;
logic signed [WIDTH-1:0] w_iz_1_0 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_1 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_2 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_3 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_4 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_5 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_1_6 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_1_7 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_1_8 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_1_9 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_10 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_11 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_12 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_13 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_14 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_15 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_16 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_1_17 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_1_18 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_19 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_1_20 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_21 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_22 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_1_23 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_24 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_25 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_26 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_27 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_1_28 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_29 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_30 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_31 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_1_32 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_33 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_1_34 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_35 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_36 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_37 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_1_38 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_1_39 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_1_40 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_41 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_42 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_43 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_44 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_45 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_46 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_47 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_48 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_49 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_50 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_51 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_52 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_53 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_1_54 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_1_55 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_1_56 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_1_57 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_1_58 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_1_59 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_60 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_1_61 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_1_62 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_1_63 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_2_0 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_2_1 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_2 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_2_3 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_4 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_2_5 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_2_6 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_2_7 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_2_8 = 'b000001011;
logic signed [WIDTH-1:0] w_iz_2_9 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_2_10 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_2_11 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_12 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_13 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_2_14 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_15 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_2_16 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_17 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_2_18 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_19 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_20 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_21 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_22 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_2_23 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_24 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_25 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_2_26 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_2_27 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_28 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_2_29 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_2_30 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_31 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_2_32 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_2_33 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_2_34 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_2_35 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_2_36 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_37 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_2_38 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_2_39 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_40 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_2_41 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_2_42 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_2_43 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_2_44 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_2_45 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_46 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_2_47 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_2_48 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_2_49 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_2_50 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_2_51 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_2_52 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_2_53 = 'b111110010;
logic signed [WIDTH-1:0] w_iz_2_54 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_55 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_2_56 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_57 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_58 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_59 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_2_60 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_2_61 = 'b111110100;
logic signed [WIDTH-1:0] w_iz_2_62 = 'b111110001;
logic signed [WIDTH-1:0] w_iz_2_63 = 'b111110000;
logic signed [WIDTH-1:0] w_iz_3_0 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_3_1 = 'b111110101;
logic signed [WIDTH-1:0] w_iz_3_2 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_3_3 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_4 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_3_5 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_3_6 = 'b111111001;
logic signed [WIDTH-1:0] w_iz_3_7 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_3_8 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_3_9 = 'b111110100;
logic signed [WIDTH-1:0] w_iz_3_10 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_3_11 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_3_12 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_3_13 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_3_14 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_3_15 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_3_16 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_3_17 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_3_18 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_3_19 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_3_20 = 'b111111100;
logic signed [WIDTH-1:0] w_iz_3_21 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_3_22 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_3_23 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_3_24 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_3_25 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_3_26 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_3_27 = 'b111111110;
logic signed [WIDTH-1:0] w_iz_3_28 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_3_29 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_3_30 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_3_31 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_3_32 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_3_33 = 'b111111101;
logic signed [WIDTH-1:0] w_iz_3_34 = 'b111110100;
logic signed [WIDTH-1:0] w_iz_3_35 = 'b111111010;
logic signed [WIDTH-1:0] w_iz_3_36 = 'b000001000;
logic signed [WIDTH-1:0] w_iz_3_37 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_3_38 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_3_39 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_3_40 = 'b000000000;
logic signed [WIDTH-1:0] w_iz_3_41 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_3_42 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_3_43 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_3_44 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_3_45 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_3_46 = 'b000010010;
logic signed [WIDTH-1:0] w_iz_3_47 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_3_48 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_3_49 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_3_50 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_3_51 = 'b000001100;
logic signed [WIDTH-1:0] w_iz_3_52 = 'b111110111;
logic signed [WIDTH-1:0] w_iz_3_53 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_3_54 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_3_55 = 'b000000001;
logic signed [WIDTH-1:0] w_iz_3_56 = 'b000010010;
logic signed [WIDTH-1:0] w_iz_3_57 = 'b000000010;
logic signed [WIDTH-1:0] w_iz_3_58 = 'b000010011;
logic signed [WIDTH-1:0] w_iz_3_59 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_3_60 = 'b111111000;
logic signed [WIDTH-1:0] w_iz_3_61 = 'b000001001;
logic signed [WIDTH-1:0] w_iz_3_62 = 'b000001100;
logic signed [WIDTH-1:0] w_iz_3_63 = 'b111111000;

logic signed [WIDTH-1:0] w_in_0_0 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_1 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_2 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_3 = 'b000000100;
logic signed [WIDTH-1:0] w_in_0_4 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_5 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_6 = 'b111111001;
logic signed [WIDTH-1:0] w_in_0_7 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_8 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_9 = 'b000000101;
logic signed [WIDTH-1:0] w_in_0_10 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_11 = 'b000000111;
logic signed [WIDTH-1:0] w_in_0_12 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_13 = 'b000000100;
logic signed [WIDTH-1:0] w_in_0_14 = 'b000000100;
logic signed [WIDTH-1:0] w_in_0_15 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_16 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_17 = 'b000000101;
logic signed [WIDTH-1:0] w_in_0_18 = 'b000001000;
logic signed [WIDTH-1:0] w_in_0_19 = 'b000000100;
logic signed [WIDTH-1:0] w_in_0_20 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_21 = 'b000000001;
logic signed [WIDTH-1:0] w_in_0_22 = 'b000000110;
logic signed [WIDTH-1:0] w_in_0_23 = 'b000000001;
logic signed [WIDTH-1:0] w_in_0_24 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_25 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_26 = 'b111111001;
logic signed [WIDTH-1:0] w_in_0_27 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_28 = 'b000000100;
logic signed [WIDTH-1:0] w_in_0_29 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_30 = 'b000000101;
logic signed [WIDTH-1:0] w_in_0_31 = 'b000000100;
logic signed [WIDTH-1:0] w_in_0_32 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_33 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_34 = 'b111111010;
logic signed [WIDTH-1:0] w_in_0_35 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_36 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_37 = 'b111110110;
logic signed [WIDTH-1:0] w_in_0_38 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_39 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_40 = 'b111111111;
logic signed [WIDTH-1:0] w_in_0_41 = 'b000000111;
logic signed [WIDTH-1:0] w_in_0_42 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_43 = 'b000000100;
logic signed [WIDTH-1:0] w_in_0_44 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_45 = 'b111111100;
logic signed [WIDTH-1:0] w_in_0_46 = 'b111111011;
logic signed [WIDTH-1:0] w_in_0_47 = 'b000000101;
logic signed [WIDTH-1:0] w_in_0_48 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_49 = 'b000001001;
logic signed [WIDTH-1:0] w_in_0_50 = 'b000000000;
logic signed [WIDTH-1:0] w_in_0_51 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_52 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_53 = 'b111111010;
logic signed [WIDTH-1:0] w_in_0_54 = 'b111111001;
logic signed [WIDTH-1:0] w_in_0_55 = 'b111111101;
logic signed [WIDTH-1:0] w_in_0_56 = 'b000000111;
logic signed [WIDTH-1:0] w_in_0_57 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_58 = 'b000001000;
logic signed [WIDTH-1:0] w_in_0_59 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_60 = 'b111110111;
logic signed [WIDTH-1:0] w_in_0_61 = 'b111110010;
logic signed [WIDTH-1:0] w_in_0_62 = 'b111110000;
logic signed [WIDTH-1:0] w_in_0_63 = 'b000000011;
logic signed [WIDTH-1:0] w_in_1_0 = 'b000000110;
logic signed [WIDTH-1:0] w_in_1_1 = 'b000000010;
logic signed [WIDTH-1:0] w_in_1_2 = 'b000000001;
logic signed [WIDTH-1:0] w_in_1_3 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_4 = 'b000000001;
logic signed [WIDTH-1:0] w_in_1_5 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_6 = 'b111111010;
logic signed [WIDTH-1:0] w_in_1_7 = 'b111111011;
logic signed [WIDTH-1:0] w_in_1_8 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_9 = 'b000001000;
logic signed [WIDTH-1:0] w_in_1_10 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_11 = 'b111111000;
logic signed [WIDTH-1:0] w_in_1_12 = 'b111111011;
logic signed [WIDTH-1:0] w_in_1_13 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_14 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_15 = 'b000000110;
logic signed [WIDTH-1:0] w_in_1_16 = 'b111111000;
logic signed [WIDTH-1:0] w_in_1_17 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_18 = 'b000001001;
logic signed [WIDTH-1:0] w_in_1_19 = 'b111111011;
logic signed [WIDTH-1:0] w_in_1_20 = 'b111111011;
logic signed [WIDTH-1:0] w_in_1_21 = 'b111111001;
logic signed [WIDTH-1:0] w_in_1_22 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_23 = 'b000001010;
logic signed [WIDTH-1:0] w_in_1_24 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_25 = 'b111111100;
logic signed [WIDTH-1:0] w_in_1_26 = 'b111111101;
logic signed [WIDTH-1:0] w_in_1_27 = 'b111111100;
logic signed [WIDTH-1:0] w_in_1_28 = 'b111111101;
logic signed [WIDTH-1:0] w_in_1_29 = 'b111111010;
logic signed [WIDTH-1:0] w_in_1_30 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_31 = 'b111111010;
logic signed [WIDTH-1:0] w_in_1_32 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_33 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_34 = 'b111111100;
logic signed [WIDTH-1:0] w_in_1_35 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_36 = 'b111110111;
logic signed [WIDTH-1:0] w_in_1_37 = 'b000000001;
logic signed [WIDTH-1:0] w_in_1_38 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_39 = 'b111111100;
logic signed [WIDTH-1:0] w_in_1_40 = 'b000000110;
logic signed [WIDTH-1:0] w_in_1_41 = 'b000000011;
logic signed [WIDTH-1:0] w_in_1_42 = 'b000000111;
logic signed [WIDTH-1:0] w_in_1_43 = 'b000000110;
logic signed [WIDTH-1:0] w_in_1_44 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_45 = 'b000000111;
logic signed [WIDTH-1:0] w_in_1_46 = 'b000000010;
logic signed [WIDTH-1:0] w_in_1_47 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_48 = 'b111111010;
logic signed [WIDTH-1:0] w_in_1_49 = 'b111111111;
logic signed [WIDTH-1:0] w_in_1_50 = 'b111111101;
logic signed [WIDTH-1:0] w_in_1_51 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_52 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_53 = 'b000000011;
logic signed [WIDTH-1:0] w_in_1_54 = 'b111111000;
logic signed [WIDTH-1:0] w_in_1_55 = 'b000001010;
logic signed [WIDTH-1:0] w_in_1_56 = 'b000000101;
logic signed [WIDTH-1:0] w_in_1_57 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_58 = 'b111111111;
logic signed [WIDTH-1:0] w_in_1_59 = 'b000000111;
logic signed [WIDTH-1:0] w_in_1_60 = 'b111110111;
logic signed [WIDTH-1:0] w_in_1_61 = 'b000000000;
logic signed [WIDTH-1:0] w_in_1_62 = 'b111111101;
logic signed [WIDTH-1:0] w_in_1_63 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_0 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_1 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_2 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_3 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_4 = 'b000000110;
logic signed [WIDTH-1:0] w_in_2_5 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_6 = 'b111110111;
logic signed [WIDTH-1:0] w_in_2_7 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_8 = 'b111110100;
logic signed [WIDTH-1:0] w_in_2_9 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_10 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_11 = 'b111111100;
logic signed [WIDTH-1:0] w_in_2_12 = 'b111111001;
logic signed [WIDTH-1:0] w_in_2_13 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_14 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_15 = 'b111110101;
logic signed [WIDTH-1:0] w_in_2_16 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_17 = 'b000000101;
logic signed [WIDTH-1:0] w_in_2_18 = 'b111110100;
logic signed [WIDTH-1:0] w_in_2_19 = 'b111111000;
logic signed [WIDTH-1:0] w_in_2_20 = 'b000000111;
logic signed [WIDTH-1:0] w_in_2_21 = 'b111111010;
logic signed [WIDTH-1:0] w_in_2_22 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_23 = 'b111111010;
logic signed [WIDTH-1:0] w_in_2_24 = 'b000000011;
logic signed [WIDTH-1:0] w_in_2_25 = 'b111111011;
logic signed [WIDTH-1:0] w_in_2_26 = 'b000001001;
logic signed [WIDTH-1:0] w_in_2_27 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_28 = 'b000000110;
logic signed [WIDTH-1:0] w_in_2_29 = 'b000001001;
logic signed [WIDTH-1:0] w_in_2_30 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_31 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_32 = 'b000001011;
logic signed [WIDTH-1:0] w_in_2_33 = 'b111111000;
logic signed [WIDTH-1:0] w_in_2_34 = 'b111111000;
logic signed [WIDTH-1:0] w_in_2_35 = 'b111111100;
logic signed [WIDTH-1:0] w_in_2_36 = 'b000001010;
logic signed [WIDTH-1:0] w_in_2_37 = 'b000001000;
logic signed [WIDTH-1:0] w_in_2_38 = 'b111111011;
logic signed [WIDTH-1:0] w_in_2_39 = 'b111110101;
logic signed [WIDTH-1:0] w_in_2_40 = 'b000000100;
logic signed [WIDTH-1:0] w_in_2_41 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_42 = 'b111111000;
logic signed [WIDTH-1:0] w_in_2_43 = 'b000000001;
logic signed [WIDTH-1:0] w_in_2_44 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_45 = 'b000000101;
logic signed [WIDTH-1:0] w_in_2_46 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_47 = 'b111111110;
logic signed [WIDTH-1:0] w_in_2_48 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_49 = 'b000000000;
logic signed [WIDTH-1:0] w_in_2_50 = 'b111111000;
logic signed [WIDTH-1:0] w_in_2_51 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_52 = 'b111111000;
logic signed [WIDTH-1:0] w_in_2_53 = 'b000000111;
logic signed [WIDTH-1:0] w_in_2_54 = 'b111111111;
logic signed [WIDTH-1:0] w_in_2_55 = 'b111111100;
logic signed [WIDTH-1:0] w_in_2_56 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_57 = 'b000000111;
logic signed [WIDTH-1:0] w_in_2_58 = 'b000001000;
logic signed [WIDTH-1:0] w_in_2_59 = 'b000001010;
logic signed [WIDTH-1:0] w_in_2_60 = 'b000001111;
logic signed [WIDTH-1:0] w_in_2_61 = 'b000001010;
logic signed [WIDTH-1:0] w_in_2_62 = 'b000010001;
logic signed [WIDTH-1:0] w_in_2_63 = 'b000001101;
logic signed [WIDTH-1:0] w_in_3_0 = 'b111110101;
logic signed [WIDTH-1:0] w_in_3_1 = 'b000001000;
logic signed [WIDTH-1:0] w_in_3_2 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_3 = 'b000001001;
logic signed [WIDTH-1:0] w_in_3_4 = 'b111110110;
logic signed [WIDTH-1:0] w_in_3_5 = 'b000000010;
logic signed [WIDTH-1:0] w_in_3_6 = 'b111110111;
logic signed [WIDTH-1:0] w_in_3_7 = 'b000000101;
logic signed [WIDTH-1:0] w_in_3_8 = 'b111110010;
logic signed [WIDTH-1:0] w_in_3_9 = 'b111110101;
logic signed [WIDTH-1:0] w_in_3_10 = 'b000001001;
logic signed [WIDTH-1:0] w_in_3_11 = 'b111110101;
logic signed [WIDTH-1:0] w_in_3_12 = 'b111110101;
logic signed [WIDTH-1:0] w_in_3_13 = 'b000000101;
logic signed [WIDTH-1:0] w_in_3_14 = 'b000000100;
logic signed [WIDTH-1:0] w_in_3_15 = 'b000000100;
logic signed [WIDTH-1:0] w_in_3_16 = 'b000001011;
logic signed [WIDTH-1:0] w_in_3_17 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_18 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_19 = 'b000001101;
logic signed [WIDTH-1:0] w_in_3_20 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_21 = 'b111111000;
logic signed [WIDTH-1:0] w_in_3_22 = 'b111111101;
logic signed [WIDTH-1:0] w_in_3_23 = 'b111111100;
logic signed [WIDTH-1:0] w_in_3_24 = 'b111110110;
logic signed [WIDTH-1:0] w_in_3_25 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_26 = 'b111111000;
logic signed [WIDTH-1:0] w_in_3_27 = 'b111110110;
logic signed [WIDTH-1:0] w_in_3_28 = 'b000001101;
logic signed [WIDTH-1:0] w_in_3_29 = 'b000000100;
logic signed [WIDTH-1:0] w_in_3_30 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_31 = 'b000000111;
logic signed [WIDTH-1:0] w_in_3_32 = 'b000000100;
logic signed [WIDTH-1:0] w_in_3_33 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_34 = 'b000000111;
logic signed [WIDTH-1:0] w_in_3_35 = 'b000000100;
logic signed [WIDTH-1:0] w_in_3_36 = 'b111110111;
logic signed [WIDTH-1:0] w_in_3_37 = 'b111110110;
logic signed [WIDTH-1:0] w_in_3_38 = 'b000000100;
logic signed [WIDTH-1:0] w_in_3_39 = 'b000000000;
logic signed [WIDTH-1:0] w_in_3_40 = 'b111110100;
logic signed [WIDTH-1:0] w_in_3_41 = 'b111110110;
logic signed [WIDTH-1:0] w_in_3_42 = 'b000001000;
logic signed [WIDTH-1:0] w_in_3_43 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_44 = 'b000000011;
logic signed [WIDTH-1:0] w_in_3_45 = 'b000001100;
logic signed [WIDTH-1:0] w_in_3_46 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_47 = 'b000001010;
logic signed [WIDTH-1:0] w_in_3_48 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_49 = 'b111111111;
logic signed [WIDTH-1:0] w_in_3_50 = 'b111111011;
logic signed [WIDTH-1:0] w_in_3_51 = 'b000000110;
logic signed [WIDTH-1:0] w_in_3_52 = 'b111111110;
logic signed [WIDTH-1:0] w_in_3_53 = 'b111110110;
logic signed [WIDTH-1:0] w_in_3_54 = 'b000001100;
logic signed [WIDTH-1:0] w_in_3_55 = 'b000000010;
logic signed [WIDTH-1:0] w_in_3_56 = 'b111111010;
logic signed [WIDTH-1:0] w_in_3_57 = 'b000000110;
logic signed [WIDTH-1:0] w_in_3_58 = 'b111111011;
logic signed [WIDTH-1:0] w_in_3_59 = 'b000001011;
logic signed [WIDTH-1:0] w_in_3_60 = 'b000001011;
logic signed [WIDTH-1:0] w_in_3_61 = 'b000000011;
logic signed [WIDTH-1:0] w_in_3_62 = 'b000000001;
logic signed [WIDTH-1:0] w_in_3_63 = 'b000001001;

// Recurrent weights (h×h for each gate)
logic signed [WIDTH-1:0] w_hr_0_0 = 'b000000000;
logic signed [WIDTH-1:0] w_hr_0_1 = 'b000000001;
logic signed [WIDTH-1:0] w_hr_0_2 = 'b000000010;
logic signed [WIDTH-1:0] w_hr_0_3 = 'b111111011;
logic signed [WIDTH-1:0] w_hr_1_0 = 'b000001001;
logic signed [WIDTH-1:0] w_hr_1_1 = 'b000001001;
logic signed [WIDTH-1:0] w_hr_1_2 = 'b000001001;
logic signed [WIDTH-1:0] w_hr_1_3 = 'b111110111;
logic signed [WIDTH-1:0] w_hr_2_0 = 'b000001000;
logic signed [WIDTH-1:0] w_hr_2_1 = 'b000001001;
logic signed [WIDTH-1:0] w_hr_2_2 = 'b111111100;
logic signed [WIDTH-1:0] w_hr_2_3 = 'b111111011;
logic signed [WIDTH-1:0] w_hr_3_0 = 'b000000100;
logic signed [WIDTH-1:0] w_hr_3_1 = 'b000000101;
logic signed [WIDTH-1:0] w_hr_3_2 = 'b000001011;
logic signed [WIDTH-1:0] w_hr_3_3 = 'b111111000;

logic signed [WIDTH-1:0] w_hz_0_0 = 'b000000111;
logic signed [WIDTH-1:0] w_hz_0_1 = 'b000000100;
logic signed [WIDTH-1:0] w_hz_0_2 = 'b111111101;
logic signed [WIDTH-1:0] w_hz_0_3 = 'b000000100;
logic signed [WIDTH-1:0] w_hz_1_0 = 'b000001101;
logic signed [WIDTH-1:0] w_hz_1_1 = 'b111110100;
logic signed [WIDTH-1:0] w_hz_1_2 = 'b000000000;
logic signed [WIDTH-1:0] w_hz_1_3 = 'b000001001;
logic signed [WIDTH-1:0] w_hz_2_0 = 'b000000111;
logic signed [WIDTH-1:0] w_hz_2_1 = 'b000000000;
logic signed [WIDTH-1:0] w_hz_2_2 = 'b111110000;
logic signed [WIDTH-1:0] w_hz_2_3 = 'b000001110;
logic signed [WIDTH-1:0] w_hz_3_0 = 'b000001100;
logic signed [WIDTH-1:0] w_hz_3_1 = 'b000000100;
logic signed [WIDTH-1:0] w_hz_3_2 = 'b111110111;
logic signed [WIDTH-1:0] w_hz_3_3 = 'b000010101;

logic signed [WIDTH-1:0] w_hn_0_0 = 'b111111111;
logic signed [WIDTH-1:0] w_hn_0_1 = 'b111111110;
logic signed [WIDTH-1:0] w_hn_0_2 = 'b000000101;
logic signed [WIDTH-1:0] w_hn_0_3 = 'b111111010;
logic signed [WIDTH-1:0] w_hn_1_0 = 'b111111010;
logic signed [WIDTH-1:0] w_hn_1_1 = 'b111111111;
logic signed [WIDTH-1:0] w_hn_1_2 = 'b000010111;
logic signed [WIDTH-1:0] w_hn_1_3 = 'b111110100;
logic signed [WIDTH-1:0] w_hn_2_0 = 'b111111111;
logic signed [WIDTH-1:0] w_hn_2_1 = 'b000001110;
logic signed [WIDTH-1:0] w_hn_2_2 = 'b000010100;
logic signed [WIDTH-1:0] w_hn_2_3 = 'b111110010;
logic signed [WIDTH-1:0] w_hn_3_0 = 'b111111011;
logic signed [WIDTH-1:0] w_hn_3_1 = 'b111110110;
logic signed [WIDTH-1:0] w_hn_3_2 = 'b111111001;
logic signed [WIDTH-1:0] w_hn_3_3 = 'b000001010;

// Biases (h for each gate type)
logic signed [WIDTH-1:0] b_ir_0 = 'b000000001;
logic signed [WIDTH-1:0] b_ir_1 = 'b000001000;
logic signed [WIDTH-1:0] b_ir_2 = 'b000001111;
logic signed [WIDTH-1:0] b_ir_3 = 'b000000101;

logic signed [WIDTH-1:0] b_iz_0 = 'b000000110;
logic signed [WIDTH-1:0] b_iz_1 = 'b000000100;
logic signed [WIDTH-1:0] b_iz_2 = 'b000010000;
logic signed [WIDTH-1:0] b_iz_3 = 'b000000000;

logic signed [WIDTH-1:0] b_in_0 = 'b000001011;
logic signed [WIDTH-1:0] b_in_1 = 'b000000010;
logic signed [WIDTH-1:0] b_in_2 = 'b000001110;
logic signed [WIDTH-1:0] b_in_3 = 'b000000010;

logic signed [WIDTH-1:0] b_hr_0 = 'b000000010;
logic signed [WIDTH-1:0] b_hr_1 = 'b000001010;
logic signed [WIDTH-1:0] b_hr_2 = 'b000000111;
logic signed [WIDTH-1:0] b_hr_3 = 'b000001101;

logic signed [WIDTH-1:0] b_hz_0 = 'b000000111;
logic signed [WIDTH-1:0] b_hz_1 = 'b000001001;
logic signed [WIDTH-1:0] b_hz_2 = 'b000000101;
logic signed [WIDTH-1:0] b_hz_3 = 'b000011010;

logic signed [WIDTH-1:0] b_hn_0 = 'b000000011;
logic signed [WIDTH-1:0] b_hn_1 = 'b000010011;
logic signed [WIDTH-1:0] b_hn_2 = 'b000000111;
logic signed [WIDTH-1:0] b_hn_3 = 'b111110001;

// Outputs (h=4)
logic signed [WIDTH-1:0]  y_0 = 0;
logic signed [WIDTH-1:0]  y_1 = 0;
logic signed [WIDTH-1:0]  y_2 = 0;
logic signed [WIDTH-1:0]  y_3 = 0;

gru #(
        .INT_WIDTH(INT_WIDTH),
        .FRAC_WIDTH(FRAC_WIDTH)
    ) gru_inst (
        .clk(clk),
        .reset(reset),
        // Input features (d=64)
        	
.x_0(x_0), .x_1(x_1), .x_2(x_2), .x_3(x_3), .x_4(x_4), .x_5(x_5), .x_6(x_6), .x_7(x_7), .x_8(x_8), .x_9(x_9), .x_10(x_10), .x_11(x_11), .x_12(x_12), .x_13(x_13), .x_14(x_14), .x_15(x_15), .x_16(x_16), .x_17(x_17), .x_18(x_18), .x_19(x_19), .x_20(x_20), .x_21(x_21), .x_22(x_22), .x_23(x_23), .x_24(x_24), .x_25(x_25), .x_26(x_26), .x_27(x_27), .x_28(x_28), .x_29(x_29), .x_30(x_30), .x_31(x_31), .x_32(x_32), .x_33(x_33), .x_34(x_34), .x_35(x_35), .x_36(x_36), .x_37(x_37), .x_38(x_38), .x_39(x_39), .x_40(x_40), .x_41(x_41), .x_42(x_42), .x_43(x_43), .x_44(x_44), .x_45(x_45), .x_46(x_46), .x_47(x_47), .x_48(x_48), .x_49(x_49), .x_50(x_50), .x_51(x_51), .x_52(x_52), .x_53(x_53), .x_54(x_54), .x_55(x_55), .x_56(x_56), .x_57(x_57), .x_58(x_58), .x_59(x_59), .x_60(x_60), .x_61(x_61), .x_62(x_62), .x_63(x_63), 	
.h_0(h_0), .h_1(h_1), .h_2(h_2), .h_3(h_3), 	
.w_ir_0_0(w_ir_0_0), .w_ir_0_1(w_ir_0_1), .w_ir_0_2(w_ir_0_2), .w_ir_0_3(w_ir_0_3), .w_ir_0_4(w_ir_0_4), .w_ir_0_5(w_ir_0_5), .w_ir_0_6(w_ir_0_6), .w_ir_0_7(w_ir_0_7), .w_ir_0_8(w_ir_0_8), .w_ir_0_9(w_ir_0_9), .w_ir_0_10(w_ir_0_10), .w_ir_0_11(w_ir_0_11), .w_ir_0_12(w_ir_0_12), .w_ir_0_13(w_ir_0_13), .w_ir_0_14(w_ir_0_14), .w_ir_0_15(w_ir_0_15), .w_ir_0_16(w_ir_0_16), .w_ir_0_17(w_ir_0_17), .w_ir_0_18(w_ir_0_18), .w_ir_0_19(w_ir_0_19), .w_ir_0_20(w_ir_0_20), .w_ir_0_21(w_ir_0_21), .w_ir_0_22(w_ir_0_22), .w_ir_0_23(w_ir_0_23), .w_ir_0_24(w_ir_0_24), .w_ir_0_25(w_ir_0_25), .w_ir_0_26(w_ir_0_26), .w_ir_0_27(w_ir_0_27), .w_ir_0_28(w_ir_0_28), .w_ir_0_29(w_ir_0_29), .w_ir_0_30(w_ir_0_30), .w_ir_0_31(w_ir_0_31), .w_ir_0_32(w_ir_0_32), .w_ir_0_33(w_ir_0_33), .w_ir_0_34(w_ir_0_34), .w_ir_0_35(w_ir_0_35), .w_ir_0_36(w_ir_0_36), .w_ir_0_37(w_ir_0_37), .w_ir_0_38(w_ir_0_38), .w_ir_0_39(w_ir_0_39), .w_ir_0_40(w_ir_0_40), .w_ir_0_41(w_ir_0_41), .w_ir_0_42(w_ir_0_42), .w_ir_0_43(w_ir_0_43), .w_ir_0_44(w_ir_0_44), .w_ir_0_45(w_ir_0_45), .w_ir_0_46(w_ir_0_46), .w_ir_0_47(w_ir_0_47), .w_ir_0_48(w_ir_0_48), .w_ir_0_49(w_ir_0_49), .w_ir_0_50(w_ir_0_50), .w_ir_0_51(w_ir_0_51), .w_ir_0_52(w_ir_0_52), .w_ir_0_53(w_ir_0_53), .w_ir_0_54(w_ir_0_54), .w_ir_0_55(w_ir_0_55), .w_ir_0_56(w_ir_0_56), .w_ir_0_57(w_ir_0_57), .w_ir_0_58(w_ir_0_58), .w_ir_0_59(w_ir_0_59), .w_ir_0_60(w_ir_0_60), .w_ir_0_61(w_ir_0_61), .w_ir_0_62(w_ir_0_62), .w_ir_0_63(w_ir_0_63), .w_ir_1_0(w_ir_1_0), .w_ir_1_1(w_ir_1_1), .w_ir_1_2(w_ir_1_2), .w_ir_1_3(w_ir_1_3), .w_ir_1_4(w_ir_1_4), .w_ir_1_5(w_ir_1_5), .w_ir_1_6(w_ir_1_6), .w_ir_1_7(w_ir_1_7), .w_ir_1_8(w_ir_1_8), .w_ir_1_9(w_ir_1_9), .w_ir_1_10(w_ir_1_10), .w_ir_1_11(w_ir_1_11), .w_ir_1_12(w_ir_1_12), .w_ir_1_13(w_ir_1_13), .w_ir_1_14(w_ir_1_14), .w_ir_1_15(w_ir_1_15), .w_ir_1_16(w_ir_1_16), .w_ir_1_17(w_ir_1_17), .w_ir_1_18(w_ir_1_18), .w_ir_1_19(w_ir_1_19), .w_ir_1_20(w_ir_1_20), .w_ir_1_21(w_ir_1_21), .w_ir_1_22(w_ir_1_22), .w_ir_1_23(w_ir_1_23), .w_ir_1_24(w_ir_1_24), .w_ir_1_25(w_ir_1_25), .w_ir_1_26(w_ir_1_26), .w_ir_1_27(w_ir_1_27), .w_ir_1_28(w_ir_1_28), .w_ir_1_29(w_ir_1_29), .w_ir_1_30(w_ir_1_30), .w_ir_1_31(w_ir_1_31), .w_ir_1_32(w_ir_1_32), .w_ir_1_33(w_ir_1_33), .w_ir_1_34(w_ir_1_34), .w_ir_1_35(w_ir_1_35), .w_ir_1_36(w_ir_1_36), .w_ir_1_37(w_ir_1_37), .w_ir_1_38(w_ir_1_38), .w_ir_1_39(w_ir_1_39), .w_ir_1_40(w_ir_1_40), .w_ir_1_41(w_ir_1_41), .w_ir_1_42(w_ir_1_42), .w_ir_1_43(w_ir_1_43), .w_ir_1_44(w_ir_1_44), .w_ir_1_45(w_ir_1_45), .w_ir_1_46(w_ir_1_46), .w_ir_1_47(w_ir_1_47), .w_ir_1_48(w_ir_1_48), .w_ir_1_49(w_ir_1_49), .w_ir_1_50(w_ir_1_50), .w_ir_1_51(w_ir_1_51), .w_ir_1_52(w_ir_1_52), .w_ir_1_53(w_ir_1_53), .w_ir_1_54(w_ir_1_54), .w_ir_1_55(w_ir_1_55), .w_ir_1_56(w_ir_1_56), .w_ir_1_57(w_ir_1_57), .w_ir_1_58(w_ir_1_58), .w_ir_1_59(w_ir_1_59), .w_ir_1_60(w_ir_1_60), .w_ir_1_61(w_ir_1_61), .w_ir_1_62(w_ir_1_62), .w_ir_1_63(w_ir_1_63), .w_ir_2_0(w_ir_2_0), .w_ir_2_1(w_ir_2_1), .w_ir_2_2(w_ir_2_2), .w_ir_2_3(w_ir_2_3), .w_ir_2_4(w_ir_2_4), .w_ir_2_5(w_ir_2_5), .w_ir_2_6(w_ir_2_6), .w_ir_2_7(w_ir_2_7), .w_ir_2_8(w_ir_2_8), .w_ir_2_9(w_ir_2_9), .w_ir_2_10(w_ir_2_10), .w_ir_2_11(w_ir_2_11), .w_ir_2_12(w_ir_2_12), .w_ir_2_13(w_ir_2_13), .w_ir_2_14(w_ir_2_14), .w_ir_2_15(w_ir_2_15), .w_ir_2_16(w_ir_2_16), .w_ir_2_17(w_ir_2_17), .w_ir_2_18(w_ir_2_18), .w_ir_2_19(w_ir_2_19), .w_ir_2_20(w_ir_2_20), .w_ir_2_21(w_ir_2_21), .w_ir_2_22(w_ir_2_22), .w_ir_2_23(w_ir_2_23), .w_ir_2_24(w_ir_2_24), .w_ir_2_25(w_ir_2_25), .w_ir_2_26(w_ir_2_26), .w_ir_2_27(w_ir_2_27), .w_ir_2_28(w_ir_2_28), .w_ir_2_29(w_ir_2_29), .w_ir_2_30(w_ir_2_30), .w_ir_2_31(w_ir_2_31), .w_ir_2_32(w_ir_2_32), .w_ir_2_33(w_ir_2_33), .w_ir_2_34(w_ir_2_34), .w_ir_2_35(w_ir_2_35), .w_ir_2_36(w_ir_2_36), .w_ir_2_37(w_ir_2_37), .w_ir_2_38(w_ir_2_38), .w_ir_2_39(w_ir_2_39), .w_ir_2_40(w_ir_2_40), .w_ir_2_41(w_ir_2_41), .w_ir_2_42(w_ir_2_42), .w_ir_2_43(w_ir_2_43), .w_ir_2_44(w_ir_2_44), .w_ir_2_45(w_ir_2_45), .w_ir_2_46(w_ir_2_46), .w_ir_2_47(w_ir_2_47), .w_ir_2_48(w_ir_2_48), .w_ir_2_49(w_ir_2_49), .w_ir_2_50(w_ir_2_50), .w_ir_2_51(w_ir_2_51), .w_ir_2_52(w_ir_2_52), .w_ir_2_53(w_ir_2_53), .w_ir_2_54(w_ir_2_54), .w_ir_2_55(w_ir_2_55), .w_ir_2_56(w_ir_2_56), .w_ir_2_57(w_ir_2_57), .w_ir_2_58(w_ir_2_58), .w_ir_2_59(w_ir_2_59), .w_ir_2_60(w_ir_2_60), .w_ir_2_61(w_ir_2_61), .w_ir_2_62(w_ir_2_62), .w_ir_2_63(w_ir_2_63), .w_ir_3_0(w_ir_3_0), .w_ir_3_1(w_ir_3_1), .w_ir_3_2(w_ir_3_2), .w_ir_3_3(w_ir_3_3), .w_ir_3_4(w_ir_3_4), .w_ir_3_5(w_ir_3_5), .w_ir_3_6(w_ir_3_6), .w_ir_3_7(w_ir_3_7), .w_ir_3_8(w_ir_3_8), .w_ir_3_9(w_ir_3_9), .w_ir_3_10(w_ir_3_10), .w_ir_3_11(w_ir_3_11), .w_ir_3_12(w_ir_3_12), .w_ir_3_13(w_ir_3_13), .w_ir_3_14(w_ir_3_14), .w_ir_3_15(w_ir_3_15), .w_ir_3_16(w_ir_3_16), .w_ir_3_17(w_ir_3_17), .w_ir_3_18(w_ir_3_18), .w_ir_3_19(w_ir_3_19), .w_ir_3_20(w_ir_3_20), .w_ir_3_21(w_ir_3_21), .w_ir_3_22(w_ir_3_22), .w_ir_3_23(w_ir_3_23), .w_ir_3_24(w_ir_3_24), .w_ir_3_25(w_ir_3_25), .w_ir_3_26(w_ir_3_26), .w_ir_3_27(w_ir_3_27), .w_ir_3_28(w_ir_3_28), .w_ir_3_29(w_ir_3_29), .w_ir_3_30(w_ir_3_30), .w_ir_3_31(w_ir_3_31), .w_ir_3_32(w_ir_3_32), .w_ir_3_33(w_ir_3_33), .w_ir_3_34(w_ir_3_34), .w_ir_3_35(w_ir_3_35), .w_ir_3_36(w_ir_3_36), .w_ir_3_37(w_ir_3_37), .w_ir_3_38(w_ir_3_38), .w_ir_3_39(w_ir_3_39), .w_ir_3_40(w_ir_3_40), .w_ir_3_41(w_ir_3_41), .w_ir_3_42(w_ir_3_42), .w_ir_3_43(w_ir_3_43), .w_ir_3_44(w_ir_3_44), .w_ir_3_45(w_ir_3_45), .w_ir_3_46(w_ir_3_46), .w_ir_3_47(w_ir_3_47), .w_ir_3_48(w_ir_3_48), .w_ir_3_49(w_ir_3_49), .w_ir_3_50(w_ir_3_50), .w_ir_3_51(w_ir_3_51), .w_ir_3_52(w_ir_3_52), .w_ir_3_53(w_ir_3_53), .w_ir_3_54(w_ir_3_54), .w_ir_3_55(w_ir_3_55), .w_ir_3_56(w_ir_3_56), .w_ir_3_57(w_ir_3_57), .w_ir_3_58(w_ir_3_58), .w_ir_3_59(w_ir_3_59), .w_ir_3_60(w_ir_3_60), .w_ir_3_61(w_ir_3_61), .w_ir_3_62(w_ir_3_62), .w_ir_3_63(w_ir_3_63), 	
.w_iz_0_0(w_iz_0_0), .w_iz_0_1(w_iz_0_1), .w_iz_0_2(w_iz_0_2), .w_iz_0_3(w_iz_0_3), .w_iz_0_4(w_iz_0_4), .w_iz_0_5(w_iz_0_5), .w_iz_0_6(w_iz_0_6), .w_iz_0_7(w_iz_0_7), .w_iz_0_8(w_iz_0_8), .w_iz_0_9(w_iz_0_9), .w_iz_0_10(w_iz_0_10), .w_iz_0_11(w_iz_0_11), .w_iz_0_12(w_iz_0_12), .w_iz_0_13(w_iz_0_13), .w_iz_0_14(w_iz_0_14), .w_iz_0_15(w_iz_0_15), .w_iz_0_16(w_iz_0_16), .w_iz_0_17(w_iz_0_17), .w_iz_0_18(w_iz_0_18), .w_iz_0_19(w_iz_0_19), .w_iz_0_20(w_iz_0_20), .w_iz_0_21(w_iz_0_21), .w_iz_0_22(w_iz_0_22), .w_iz_0_23(w_iz_0_23), .w_iz_0_24(w_iz_0_24), .w_iz_0_25(w_iz_0_25), .w_iz_0_26(w_iz_0_26), .w_iz_0_27(w_iz_0_27), .w_iz_0_28(w_iz_0_28), .w_iz_0_29(w_iz_0_29), .w_iz_0_30(w_iz_0_30), .w_iz_0_31(w_iz_0_31), .w_iz_0_32(w_iz_0_32), .w_iz_0_33(w_iz_0_33), .w_iz_0_34(w_iz_0_34), .w_iz_0_35(w_iz_0_35), .w_iz_0_36(w_iz_0_36), .w_iz_0_37(w_iz_0_37), .w_iz_0_38(w_iz_0_38), .w_iz_0_39(w_iz_0_39), .w_iz_0_40(w_iz_0_40), .w_iz_0_41(w_iz_0_41), .w_iz_0_42(w_iz_0_42), .w_iz_0_43(w_iz_0_43), .w_iz_0_44(w_iz_0_44), .w_iz_0_45(w_iz_0_45), .w_iz_0_46(w_iz_0_46), .w_iz_0_47(w_iz_0_47), .w_iz_0_48(w_iz_0_48), .w_iz_0_49(w_iz_0_49), .w_iz_0_50(w_iz_0_50), .w_iz_0_51(w_iz_0_51), .w_iz_0_52(w_iz_0_52), .w_iz_0_53(w_iz_0_53), .w_iz_0_54(w_iz_0_54), .w_iz_0_55(w_iz_0_55), .w_iz_0_56(w_iz_0_56), .w_iz_0_57(w_iz_0_57), .w_iz_0_58(w_iz_0_58), .w_iz_0_59(w_iz_0_59), .w_iz_0_60(w_iz_0_60), .w_iz_0_61(w_iz_0_61), .w_iz_0_62(w_iz_0_62), .w_iz_0_63(w_iz_0_63), .w_iz_1_0(w_iz_1_0), .w_iz_1_1(w_iz_1_1), .w_iz_1_2(w_iz_1_2), .w_iz_1_3(w_iz_1_3), .w_iz_1_4(w_iz_1_4), .w_iz_1_5(w_iz_1_5), .w_iz_1_6(w_iz_1_6), .w_iz_1_7(w_iz_1_7), .w_iz_1_8(w_iz_1_8), .w_iz_1_9(w_iz_1_9), .w_iz_1_10(w_iz_1_10), .w_iz_1_11(w_iz_1_11), .w_iz_1_12(w_iz_1_12), .w_iz_1_13(w_iz_1_13), .w_iz_1_14(w_iz_1_14), .w_iz_1_15(w_iz_1_15), .w_iz_1_16(w_iz_1_16), .w_iz_1_17(w_iz_1_17), .w_iz_1_18(w_iz_1_18), .w_iz_1_19(w_iz_1_19), .w_iz_1_20(w_iz_1_20), .w_iz_1_21(w_iz_1_21), .w_iz_1_22(w_iz_1_22), .w_iz_1_23(w_iz_1_23), .w_iz_1_24(w_iz_1_24), .w_iz_1_25(w_iz_1_25), .w_iz_1_26(w_iz_1_26), .w_iz_1_27(w_iz_1_27), .w_iz_1_28(w_iz_1_28), .w_iz_1_29(w_iz_1_29), .w_iz_1_30(w_iz_1_30), .w_iz_1_31(w_iz_1_31), .w_iz_1_32(w_iz_1_32), .w_iz_1_33(w_iz_1_33), .w_iz_1_34(w_iz_1_34), .w_iz_1_35(w_iz_1_35), .w_iz_1_36(w_iz_1_36), .w_iz_1_37(w_iz_1_37), .w_iz_1_38(w_iz_1_38), .w_iz_1_39(w_iz_1_39), .w_iz_1_40(w_iz_1_40), .w_iz_1_41(w_iz_1_41), .w_iz_1_42(w_iz_1_42), .w_iz_1_43(w_iz_1_43), .w_iz_1_44(w_iz_1_44), .w_iz_1_45(w_iz_1_45), .w_iz_1_46(w_iz_1_46), .w_iz_1_47(w_iz_1_47), .w_iz_1_48(w_iz_1_48), .w_iz_1_49(w_iz_1_49), .w_iz_1_50(w_iz_1_50), .w_iz_1_51(w_iz_1_51), .w_iz_1_52(w_iz_1_52), .w_iz_1_53(w_iz_1_53), .w_iz_1_54(w_iz_1_54), .w_iz_1_55(w_iz_1_55), .w_iz_1_56(w_iz_1_56), .w_iz_1_57(w_iz_1_57), .w_iz_1_58(w_iz_1_58), .w_iz_1_59(w_iz_1_59), .w_iz_1_60(w_iz_1_60), .w_iz_1_61(w_iz_1_61), .w_iz_1_62(w_iz_1_62), .w_iz_1_63(w_iz_1_63), .w_iz_2_0(w_iz_2_0), .w_iz_2_1(w_iz_2_1), .w_iz_2_2(w_iz_2_2), .w_iz_2_3(w_iz_2_3), .w_iz_2_4(w_iz_2_4), .w_iz_2_5(w_iz_2_5), .w_iz_2_6(w_iz_2_6), .w_iz_2_7(w_iz_2_7), .w_iz_2_8(w_iz_2_8), .w_iz_2_9(w_iz_2_9), .w_iz_2_10(w_iz_2_10), .w_iz_2_11(w_iz_2_11), .w_iz_2_12(w_iz_2_12), .w_iz_2_13(w_iz_2_13), .w_iz_2_14(w_iz_2_14), .w_iz_2_15(w_iz_2_15), .w_iz_2_16(w_iz_2_16), .w_iz_2_17(w_iz_2_17), .w_iz_2_18(w_iz_2_18), .w_iz_2_19(w_iz_2_19), .w_iz_2_20(w_iz_2_20), .w_iz_2_21(w_iz_2_21), .w_iz_2_22(w_iz_2_22), .w_iz_2_23(w_iz_2_23), .w_iz_2_24(w_iz_2_24), .w_iz_2_25(w_iz_2_25), .w_iz_2_26(w_iz_2_26), .w_iz_2_27(w_iz_2_27), .w_iz_2_28(w_iz_2_28), .w_iz_2_29(w_iz_2_29), .w_iz_2_30(w_iz_2_30), .w_iz_2_31(w_iz_2_31), .w_iz_2_32(w_iz_2_32), .w_iz_2_33(w_iz_2_33), .w_iz_2_34(w_iz_2_34), .w_iz_2_35(w_iz_2_35), .w_iz_2_36(w_iz_2_36), .w_iz_2_37(w_iz_2_37), .w_iz_2_38(w_iz_2_38), .w_iz_2_39(w_iz_2_39), .w_iz_2_40(w_iz_2_40), .w_iz_2_41(w_iz_2_41), .w_iz_2_42(w_iz_2_42), .w_iz_2_43(w_iz_2_43), .w_iz_2_44(w_iz_2_44), .w_iz_2_45(w_iz_2_45), .w_iz_2_46(w_iz_2_46), .w_iz_2_47(w_iz_2_47), .w_iz_2_48(w_iz_2_48), .w_iz_2_49(w_iz_2_49), .w_iz_2_50(w_iz_2_50), .w_iz_2_51(w_iz_2_51), .w_iz_2_52(w_iz_2_52), .w_iz_2_53(w_iz_2_53), .w_iz_2_54(w_iz_2_54), .w_iz_2_55(w_iz_2_55), .w_iz_2_56(w_iz_2_56), .w_iz_2_57(w_iz_2_57), .w_iz_2_58(w_iz_2_58), .w_iz_2_59(w_iz_2_59), .w_iz_2_60(w_iz_2_60), .w_iz_2_61(w_iz_2_61), .w_iz_2_62(w_iz_2_62), .w_iz_2_63(w_iz_2_63), .w_iz_3_0(w_iz_3_0), .w_iz_3_1(w_iz_3_1), .w_iz_3_2(w_iz_3_2), .w_iz_3_3(w_iz_3_3), .w_iz_3_4(w_iz_3_4), .w_iz_3_5(w_iz_3_5), .w_iz_3_6(w_iz_3_6), .w_iz_3_7(w_iz_3_7), .w_iz_3_8(w_iz_3_8), .w_iz_3_9(w_iz_3_9), .w_iz_3_10(w_iz_3_10), .w_iz_3_11(w_iz_3_11), .w_iz_3_12(w_iz_3_12), .w_iz_3_13(w_iz_3_13), .w_iz_3_14(w_iz_3_14), .w_iz_3_15(w_iz_3_15), .w_iz_3_16(w_iz_3_16), .w_iz_3_17(w_iz_3_17), .w_iz_3_18(w_iz_3_18), .w_iz_3_19(w_iz_3_19), .w_iz_3_20(w_iz_3_20), .w_iz_3_21(w_iz_3_21), .w_iz_3_22(w_iz_3_22), .w_iz_3_23(w_iz_3_23), .w_iz_3_24(w_iz_3_24), .w_iz_3_25(w_iz_3_25), .w_iz_3_26(w_iz_3_26), .w_iz_3_27(w_iz_3_27), .w_iz_3_28(w_iz_3_28), .w_iz_3_29(w_iz_3_29), .w_iz_3_30(w_iz_3_30), .w_iz_3_31(w_iz_3_31), .w_iz_3_32(w_iz_3_32), .w_iz_3_33(w_iz_3_33), .w_iz_3_34(w_iz_3_34), .w_iz_3_35(w_iz_3_35), .w_iz_3_36(w_iz_3_36), .w_iz_3_37(w_iz_3_37), .w_iz_3_38(w_iz_3_38), .w_iz_3_39(w_iz_3_39), .w_iz_3_40(w_iz_3_40), .w_iz_3_41(w_iz_3_41), .w_iz_3_42(w_iz_3_42), .w_iz_3_43(w_iz_3_43), .w_iz_3_44(w_iz_3_44), .w_iz_3_45(w_iz_3_45), .w_iz_3_46(w_iz_3_46), .w_iz_3_47(w_iz_3_47), .w_iz_3_48(w_iz_3_48), .w_iz_3_49(w_iz_3_49), .w_iz_3_50(w_iz_3_50), .w_iz_3_51(w_iz_3_51), .w_iz_3_52(w_iz_3_52), .w_iz_3_53(w_iz_3_53), .w_iz_3_54(w_iz_3_54), .w_iz_3_55(w_iz_3_55), .w_iz_3_56(w_iz_3_56), .w_iz_3_57(w_iz_3_57), .w_iz_3_58(w_iz_3_58), .w_iz_3_59(w_iz_3_59), .w_iz_3_60(w_iz_3_60), .w_iz_3_61(w_iz_3_61), .w_iz_3_62(w_iz_3_62), .w_iz_3_63(w_iz_3_63), 
.w_in_0_0(w_in_0_0), .w_in_0_1(w_in_0_1), .w_in_0_2(w_in_0_2), .w_in_0_3(w_in_0_3), .w_in_0_4(w_in_0_4), .w_in_0_5(w_in_0_5), .w_in_0_6(w_in_0_6), .w_in_0_7(w_in_0_7), .w_in_0_8(w_in_0_8), .w_in_0_9(w_in_0_9), .w_in_0_10(w_in_0_10), .w_in_0_11(w_in_0_11), .w_in_0_12(w_in_0_12), .w_in_0_13(w_in_0_13), .w_in_0_14(w_in_0_14), .w_in_0_15(w_in_0_15), .w_in_0_16(w_in_0_16), .w_in_0_17(w_in_0_17), .w_in_0_18(w_in_0_18), .w_in_0_19(w_in_0_19), .w_in_0_20(w_in_0_20), .w_in_0_21(w_in_0_21), .w_in_0_22(w_in_0_22), .w_in_0_23(w_in_0_23), .w_in_0_24(w_in_0_24), .w_in_0_25(w_in_0_25), .w_in_0_26(w_in_0_26), .w_in_0_27(w_in_0_27), .w_in_0_28(w_in_0_28), .w_in_0_29(w_in_0_29), .w_in_0_30(w_in_0_30), .w_in_0_31(w_in_0_31), .w_in_0_32(w_in_0_32), .w_in_0_33(w_in_0_33), .w_in_0_34(w_in_0_34), .w_in_0_35(w_in_0_35), .w_in_0_36(w_in_0_36), .w_in_0_37(w_in_0_37), .w_in_0_38(w_in_0_38), .w_in_0_39(w_in_0_39), .w_in_0_40(w_in_0_40), .w_in_0_41(w_in_0_41), .w_in_0_42(w_in_0_42), .w_in_0_43(w_in_0_43), .w_in_0_44(w_in_0_44), .w_in_0_45(w_in_0_45), .w_in_0_46(w_in_0_46), .w_in_0_47(w_in_0_47), .w_in_0_48(w_in_0_48), .w_in_0_49(w_in_0_49), .w_in_0_50(w_in_0_50), .w_in_0_51(w_in_0_51), .w_in_0_52(w_in_0_52), .w_in_0_53(w_in_0_53), .w_in_0_54(w_in_0_54), .w_in_0_55(w_in_0_55), .w_in_0_56(w_in_0_56), .w_in_0_57(w_in_0_57), .w_in_0_58(w_in_0_58), .w_in_0_59(w_in_0_59), .w_in_0_60(w_in_0_60), .w_in_0_61(w_in_0_61), .w_in_0_62(w_in_0_62), .w_in_0_63(w_in_0_63), .w_in_1_0(w_in_1_0), .w_in_1_1(w_in_1_1), .w_in_1_2(w_in_1_2), .w_in_1_3(w_in_1_3), .w_in_1_4(w_in_1_4), .w_in_1_5(w_in_1_5), .w_in_1_6(w_in_1_6), .w_in_1_7(w_in_1_7), .w_in_1_8(w_in_1_8), .w_in_1_9(w_in_1_9), .w_in_1_10(w_in_1_10), .w_in_1_11(w_in_1_11), .w_in_1_12(w_in_1_12), .w_in_1_13(w_in_1_13), .w_in_1_14(w_in_1_14), .w_in_1_15(w_in_1_15), .w_in_1_16(w_in_1_16), .w_in_1_17(w_in_1_17), .w_in_1_18(w_in_1_18), .w_in_1_19(w_in_1_19), .w_in_1_20(w_in_1_20), .w_in_1_21(w_in_1_21), .w_in_1_22(w_in_1_22), .w_in_1_23(w_in_1_23), .w_in_1_24(w_in_1_24), .w_in_1_25(w_in_1_25), .w_in_1_26(w_in_1_26), .w_in_1_27(w_in_1_27), .w_in_1_28(w_in_1_28), .w_in_1_29(w_in_1_29), .w_in_1_30(w_in_1_30), .w_in_1_31(w_in_1_31), .w_in_1_32(w_in_1_32), .w_in_1_33(w_in_1_33), .w_in_1_34(w_in_1_34), .w_in_1_35(w_in_1_35), .w_in_1_36(w_in_1_36), .w_in_1_37(w_in_1_37), .w_in_1_38(w_in_1_38), .w_in_1_39(w_in_1_39), .w_in_1_40(w_in_1_40), .w_in_1_41(w_in_1_41), .w_in_1_42(w_in_1_42), .w_in_1_43(w_in_1_43), .w_in_1_44(w_in_1_44), .w_in_1_45(w_in_1_45), .w_in_1_46(w_in_1_46), .w_in_1_47(w_in_1_47), .w_in_1_48(w_in_1_48), .w_in_1_49(w_in_1_49), .w_in_1_50(w_in_1_50), .w_in_1_51(w_in_1_51), .w_in_1_52(w_in_1_52), .w_in_1_53(w_in_1_53), .w_in_1_54(w_in_1_54), .w_in_1_55(w_in_1_55), .w_in_1_56(w_in_1_56), .w_in_1_57(w_in_1_57), .w_in_1_58(w_in_1_58), .w_in_1_59(w_in_1_59), .w_in_1_60(w_in_1_60), .w_in_1_61(w_in_1_61), .w_in_1_62(w_in_1_62), .w_in_1_63(w_in_1_63), .w_in_2_0(w_in_2_0), .w_in_2_1(w_in_2_1), .w_in_2_2(w_in_2_2), .w_in_2_3(w_in_2_3), .w_in_2_4(w_in_2_4), .w_in_2_5(w_in_2_5), .w_in_2_6(w_in_2_6), .w_in_2_7(w_in_2_7), .w_in_2_8(w_in_2_8), .w_in_2_9(w_in_2_9), .w_in_2_10(w_in_2_10), .w_in_2_11(w_in_2_11), .w_in_2_12(w_in_2_12), .w_in_2_13(w_in_2_13), .w_in_2_14(w_in_2_14), .w_in_2_15(w_in_2_15), .w_in_2_16(w_in_2_16), .w_in_2_17(w_in_2_17), .w_in_2_18(w_in_2_18), .w_in_2_19(w_in_2_19), .w_in_2_20(w_in_2_20), .w_in_2_21(w_in_2_21), .w_in_2_22(w_in_2_22), .w_in_2_23(w_in_2_23), .w_in_2_24(w_in_2_24), .w_in_2_25(w_in_2_25), .w_in_2_26(w_in_2_26), .w_in_2_27(w_in_2_27), .w_in_2_28(w_in_2_28), .w_in_2_29(w_in_2_29), .w_in_2_30(w_in_2_30), .w_in_2_31(w_in_2_31), .w_in_2_32(w_in_2_32), .w_in_2_33(w_in_2_33), .w_in_2_34(w_in_2_34), .w_in_2_35(w_in_2_35), .w_in_2_36(w_in_2_36), .w_in_2_37(w_in_2_37), .w_in_2_38(w_in_2_38), .w_in_2_39(w_in_2_39), .w_in_2_40(w_in_2_40), .w_in_2_41(w_in_2_41), .w_in_2_42(w_in_2_42), .w_in_2_43(w_in_2_43), .w_in_2_44(w_in_2_44), .w_in_2_45(w_in_2_45), .w_in_2_46(w_in_2_46), .w_in_2_47(w_in_2_47), .w_in_2_48(w_in_2_48), .w_in_2_49(w_in_2_49), .w_in_2_50(w_in_2_50), .w_in_2_51(w_in_2_51), .w_in_2_52(w_in_2_52), .w_in_2_53(w_in_2_53), .w_in_2_54(w_in_2_54), .w_in_2_55(w_in_2_55), .w_in_2_56(w_in_2_56), .w_in_2_57(w_in_2_57), .w_in_2_58(w_in_2_58), .w_in_2_59(w_in_2_59), .w_in_2_60(w_in_2_60), .w_in_2_61(w_in_2_61), .w_in_2_62(w_in_2_62), .w_in_2_63(w_in_2_63), .w_in_3_0(w_in_3_0), .w_in_3_1(w_in_3_1), .w_in_3_2(w_in_3_2), .w_in_3_3(w_in_3_3), .w_in_3_4(w_in_3_4), .w_in_3_5(w_in_3_5), .w_in_3_6(w_in_3_6), .w_in_3_7(w_in_3_7), .w_in_3_8(w_in_3_8), .w_in_3_9(w_in_3_9), .w_in_3_10(w_in_3_10), .w_in_3_11(w_in_3_11), .w_in_3_12(w_in_3_12), .w_in_3_13(w_in_3_13), .w_in_3_14(w_in_3_14), .w_in_3_15(w_in_3_15), .w_in_3_16(w_in_3_16), .w_in_3_17(w_in_3_17), .w_in_3_18(w_in_3_18), .w_in_3_19(w_in_3_19), .w_in_3_20(w_in_3_20), .w_in_3_21(w_in_3_21), .w_in_3_22(w_in_3_22), .w_in_3_23(w_in_3_23), .w_in_3_24(w_in_3_24), .w_in_3_25(w_in_3_25), .w_in_3_26(w_in_3_26), .w_in_3_27(w_in_3_27), .w_in_3_28(w_in_3_28), .w_in_3_29(w_in_3_29), .w_in_3_30(w_in_3_30), .w_in_3_31(w_in_3_31), .w_in_3_32(w_in_3_32), .w_in_3_33(w_in_3_33), .w_in_3_34(w_in_3_34), .w_in_3_35(w_in_3_35), .w_in_3_36(w_in_3_36), .w_in_3_37(w_in_3_37), .w_in_3_38(w_in_3_38), .w_in_3_39(w_in_3_39), .w_in_3_40(w_in_3_40), .w_in_3_41(w_in_3_41), .w_in_3_42(w_in_3_42), .w_in_3_43(w_in_3_43), .w_in_3_44(w_in_3_44), .w_in_3_45(w_in_3_45), .w_in_3_46(w_in_3_46), .w_in_3_47(w_in_3_47), .w_in_3_48(w_in_3_48), .w_in_3_49(w_in_3_49), .w_in_3_50(w_in_3_50), .w_in_3_51(w_in_3_51), .w_in_3_52(w_in_3_52), .w_in_3_53(w_in_3_53), .w_in_3_54(w_in_3_54), .w_in_3_55(w_in_3_55), .w_in_3_56(w_in_3_56), .w_in_3_57(w_in_3_57), .w_in_3_58(w_in_3_58), .w_in_3_59(w_in_3_59), .w_in_3_60(w_in_3_60), .w_in_3_61(w_in_3_61), .w_in_3_62(w_in_3_62), .w_in_3_63(w_in_3_63), 
.w_hr_0_0(w_hr_0_0), .w_hr_0_1(w_hr_0_1), .w_hr_0_2(w_hr_0_2), .w_hr_0_3(w_hr_0_3), .w_hr_1_0(w_hr_1_0), .w_hr_1_1(w_hr_1_1), .w_hr_1_2(w_hr_1_2), .w_hr_1_3(w_hr_1_3), .w_hr_2_0(w_hr_2_0), .w_hr_2_1(w_hr_2_1), .w_hr_2_2(w_hr_2_2), .w_hr_2_3(w_hr_2_3), .w_hr_3_0(w_hr_3_0), .w_hr_3_1(w_hr_3_1), .w_hr_3_2(w_hr_3_2), .w_hr_3_3(w_hr_3_3), 
.w_hz_0_0(w_hz_0_0), .w_hz_0_1(w_hz_0_1), .w_hz_0_2(w_hz_0_2), .w_hz_0_3(w_hz_0_3), .w_hz_1_0(w_hz_1_0), .w_hz_1_1(w_hz_1_1), .w_hz_1_2(w_hz_1_2), .w_hz_1_3(w_hz_1_3), .w_hz_2_0(w_hz_2_0), .w_hz_2_1(w_hz_2_1), .w_hz_2_2(w_hz_2_2), .w_hz_2_3(w_hz_2_3), .w_hz_3_0(w_hz_3_0), .w_hz_3_1(w_hz_3_1), .w_hz_3_2(w_hz_3_2), .w_hz_3_3(w_hz_3_3), 
.w_hn_0_0(w_hn_0_0), .w_hn_0_1(w_hn_0_1), .w_hn_0_2(w_hn_0_2), .w_hn_0_3(w_hn_0_3), .w_hn_1_0(w_hn_1_0), .w_hn_1_1(w_hn_1_1), .w_hn_1_2(w_hn_1_2), .w_hn_1_3(w_hn_1_3), .w_hn_2_0(w_hn_2_0), .w_hn_2_1(w_hn_2_1), .w_hn_2_2(w_hn_2_2), .w_hn_2_3(w_hn_2_3), .w_hn_3_0(w_hn_3_0), .w_hn_3_1(w_hn_3_1), .w_hn_3_2(w_hn_3_2), .w_hn_3_3(w_hn_3_3), 
.b_ir_0(b_ir_0), .b_ir_1(b_ir_1), .b_ir_2(b_ir_2), .b_ir_3(b_ir_3), 
.b_iz_0(b_iz_0), .b_iz_1(b_iz_1), .b_iz_2(b_iz_2), .b_iz_3(b_iz_3), 
.b_in_0(b_in_0), .b_in_1(b_in_1), .b_in_2(b_in_2), .b_in_3(b_in_3), 
.b_hr_0(b_hr_0), .b_hr_1(b_hr_1), .b_hr_2(b_hr_2), .b_hr_3(b_hr_3), 
.b_hz_0(b_hz_0), .b_hz_1(b_hz_1), .b_hz_2(b_hz_2), .b_hz_3(b_hz_3), 
.b_hn_0(b_hn_0), .b_hn_1(b_hn_1), .b_hn_2(b_hn_2), .b_hn_3(b_hn_3), 
.y_0(y_0), .y_1(y_1), .y_2(y_2), .y_3(y_3)
);

    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end
    
    initial begin
        // Open file for writing (overwrite existing)
        integer fd;
        fd = $fopen("../../../../../output_d64_h4_int4_frac5.txt", "w+");
        if (fd == 0) begin
            $display("ERROR: Failed to open file!");
            $finish;
        end
        x_0 = 'b000100100;
    x_1 = 'b000110111;
    x_2 = 'b001000001;
    x_3 = 'b001001001;
    x_4 = 'b000111011;
    x_5 = 'b000110110;
    x_6 = 'b000100111;
    x_7 = 'b000100101;
    x_8 = 'b000111100;
    x_9 = 'b001001000;
    x_10 = 'b001001011;
    x_11 = 'b001001001;
    x_12 = 'b001000111;
    x_13 = 'b000101101;
    x_14 = 'b000111011;
    x_15 = 'b001000110;
    x_16 = 'b001001010;
    x_17 = 'b001001101;
    x_18 = 'b001001111;
    x_19 = 'b001001110;
    x_20 = 'b000110111;
    x_21 = 'b000010001;
    x_22 = 'b000010100;
    x_23 = 'b000010111;
    x_24 = 'b000001100;
    x_25 = 'b000001110;
    x_26 = 'b000101001;
    x_27 = 'b000011100;
    x_28 = 'b000011110;
    x_29 = 'b000001100;
    x_30 = 'b000011000;
    x_31 = 'b000110010;
    x_32 = 'b000111110;
    x_33 = 'b000111110;
    x_34 = 'b000111000;
    x_35 = 'b000101111;
    x_36 = 'b000101000;
    x_37 = 'b000010100;
    x_38 = 'b000010111;
    x_39 = 'b000100100;
    x_40 = 'b000101010;
    x_41 = 'b000110100;
    x_42 = 'b000100000;
    x_43 = 'b000011011;
    x_44 = 'b000110001;
    x_45 = 'b000010111;
    x_46 = 'b000111011;
    x_47 = 'b001000011;
    x_48 = 'b000111111;
    x_49 = 'b001000110;
    x_50 = 'b001010001;
    x_51 = 'b001010101;
    x_52 = 'b001010001;
    x_53 = 'b001000110;
    x_54 = 'b000110111;
    x_55 = 'b000110111;
    x_56 = 'b001000011;
    x_57 = 'b001000110;
    x_58 = 'b001001001;
    x_59 = 'b000101111;
    x_60 = 'b000110000;
    x_61 = 'b000110011;
    x_62 = 'b000100101;
    x_63 = 'b000110000;

    h_0 = 'b000100100;
    h_1 = 'b000110111;
    h_2 = 'b001000001;
    h_3 = 'b001001001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000101110;
    x_1 = 'b001001001;
    x_2 = 'b001010010;
    x_3 = 'b001010101;
    x_4 = 'b001001111;
    x_5 = 'b001001100;
    x_6 = 'b000111111;
    x_7 = 'b000110111;
    x_8 = 'b001010001;
    x_9 = 'b001011010;
    x_10 = 'b001011011;
    x_11 = 'b001011111;
    x_12 = 'b001011010;
    x_13 = 'b001000000;
    x_14 = 'b001001101;
    x_15 = 'b001010111;
    x_16 = 'b001011000;
    x_17 = 'b001011101;
    x_18 = 'b001011110;
    x_19 = 'b001011101;
    x_20 = 'b001000011;
    x_21 = 'b000010011;
    x_22 = 'b000010100;
    x_23 = 'b000010110;
    x_24 = 'b000011000;
    x_25 = 'b000011010;
    x_26 = 'b000101101;
    x_27 = 'b000100001;
    x_28 = 'b000011010;
    x_29 = 'b000100011;
    x_30 = 'b000101010;
    x_31 = 'b000111000;
    x_32 = 'b001000010;
    x_33 = 'b001000000;
    x_34 = 'b000111010;
    x_35 = 'b000110101;
    x_36 = 'b000101001;
    x_37 = 'b000011001;
    x_38 = 'b000110101;
    x_39 = 'b000010110;
    x_40 = 'b001000010;
    x_41 = 'b111111101;
    x_42 = 'b000111010;
    x_43 = 'b000100101;
    x_44 = 'b001001000;
    x_45 = 'b000000101;
    x_46 = 'b001001001;
    x_47 = 'b001001001;
    x_48 = 'b001000000;
    x_49 = 'b001000001;
    x_50 = 'b001001110;
    x_51 = 'b001010010;
    x_52 = 'b001001001;
    x_53 = 'b000111100;
    x_54 = 'b000101010;
    x_55 = 'b000110101;
    x_56 = 'b000111110;
    x_57 = 'b000111110;
    x_58 = 'b001000010;
    x_59 = 'b000101001;
    x_60 = 'b000101110;
    x_61 = 'b000110100;
    x_62 = 'b000100110;
    x_63 = 'b000101101;

    h_0 = 'b000101110;
    h_1 = 'b001001001;
    h_2 = 'b001010010;
    h_3 = 'b001010101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000111111;
    x_1 = 'b001000011;
    x_2 = 'b001000001;
    x_3 = 'b001000000;
    x_4 = 'b000110111;
    x_5 = 'b000101101;
    x_6 = 'b000011110;
    x_7 = 'b000110010;
    x_8 = 'b001000010;
    x_9 = 'b001000001;
    x_10 = 'b001000000;
    x_11 = 'b001000011;
    x_12 = 'b000110100;
    x_13 = 'b000001110;
    x_14 = 'b001000001;
    x_15 = 'b001000010;
    x_16 = 'b001000001;
    x_17 = 'b001000011;
    x_18 = 'b001000001;
    x_19 = 'b000111100;
    x_20 = 'b000011101;
    x_21 = 'b000100001;
    x_22 = 'b000011010;
    x_23 = 'b000010111;
    x_24 = 'b000101100;
    x_25 = 'b000101101;
    x_26 = 'b000100100;
    x_27 = 'b000011100;
    x_28 = 'b000011000;
    x_29 = 'b000111011;
    x_30 = 'b000101011;
    x_31 = 'b000101001;
    x_32 = 'b000110011;
    x_33 = 'b000101110;
    x_34 = 'b000100111;
    x_35 = 'b000100010;
    x_36 = 'b000011001;
    x_37 = 'b000010010;
    x_38 = 'b000110100;
    x_39 = 'b000000010;
    x_40 = 'b000111000;
    x_41 = 'b000000001;
    x_42 = 'b000110110;
    x_43 = 'b000100010;
    x_44 = 'b000111100;
    x_45 = 'b000000100;
    x_46 = 'b000111010;
    x_47 = 'b000110111;
    x_48 = 'b000101011;
    x_49 = 'b000101100;
    x_50 = 'b000111000;
    x_51 = 'b000111011;
    x_52 = 'b000110011;
    x_53 = 'b000101011;
    x_54 = 'b000100010;
    x_55 = 'b000100101;
    x_56 = 'b000110000;
    x_57 = 'b000101110;
    x_58 = 'b000110101;
    x_59 = 'b000100101;
    x_60 = 'b000100110;
    x_61 = 'b000101110;
    x_62 = 'b000100010;
    x_63 = 'b000101110;

    h_0 = 'b000111111;
    h_1 = 'b001000011;
    h_2 = 'b001000001;
    h_3 = 'b001000000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000101101;
    x_1 = 'b000101111;
    x_2 = 'b000110100;
    x_3 = 'b000111010;
    x_4 = 'b000110001;
    x_5 = 'b000100100;
    x_6 = 'b000011100;
    x_7 = 'b000011111;
    x_8 = 'b000110001;
    x_9 = 'b000110101;
    x_10 = 'b000111000;
    x_11 = 'b000111100;
    x_12 = 'b000101011;
    x_13 = 'b000010001;
    x_14 = 'b000101110;
    x_15 = 'b000110110;
    x_16 = 'b000110101;
    x_17 = 'b000110110;
    x_18 = 'b000110111;
    x_19 = 'b000110010;
    x_20 = 'b000011100;
    x_21 = 'b000011011;
    x_22 = 'b000011001;
    x_23 = 'b000011111;
    x_24 = 'b000100000;
    x_25 = 'b000100010;
    x_26 = 'b000100110;
    x_27 = 'b000100010;
    x_28 = 'b000100100;
    x_29 = 'b000100001;
    x_30 = 'b000011111;
    x_31 = 'b000101000;
    x_32 = 'b000110001;
    x_33 = 'b000110000;
    x_34 = 'b000101100;
    x_35 = 'b000100101;
    x_36 = 'b000100011;
    x_37 = 'b000011011;
    x_38 = 'b000011100;
    x_39 = 'b000011100;
    x_40 = 'b000110001;
    x_41 = 'b000101101;
    x_42 = 'b000100001;
    x_43 = 'b000001101;
    x_44 = 'b000100010;
    x_45 = 'b000001111;
    x_46 = 'b000100011;
    x_47 = 'b000101001;
    x_48 = 'b000100011;
    x_49 = 'b000100100;
    x_50 = 'b000101100;
    x_51 = 'b000101110;
    x_52 = 'b000100111;
    x_53 = 'b000100100;
    x_54 = 'b000011111;
    x_55 = 'b000011101;
    x_56 = 'b000100111;
    x_57 = 'b000100111;
    x_58 = 'b000101100;
    x_59 = 'b000100001;
    x_60 = 'b000011101;
    x_61 = 'b000100111;
    x_62 = 'b000011010;
    x_63 = 'b000101110;

    h_0 = 'b000101101;
    h_1 = 'b000101111;
    h_2 = 'b000110100;
    h_3 = 'b000111010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000011100;
    x_1 = 'b000100110;
    x_2 = 'b000101001;
    x_3 = 'b000110001;
    x_4 = 'b000101100;
    x_5 = 'b000100000;
    x_6 = 'b000011101;
    x_7 = 'b000010100;
    x_8 = 'b000100001;
    x_9 = 'b000100111;
    x_10 = 'b000101010;
    x_11 = 'b000110000;
    x_12 = 'b000100001;
    x_13 = 'b000010000;
    x_14 = 'b000100010;
    x_15 = 'b000101000;
    x_16 = 'b000101000;
    x_17 = 'b000101000;
    x_18 = 'b000100111;
    x_19 = 'b000100010;
    x_20 = 'b000010010;
    x_21 = 'b000011111;
    x_22 = 'b000010101;
    x_23 = 'b000011011;
    x_24 = 'b000010110;
    x_25 = 'b000010111;
    x_26 = 'b000100000;
    x_27 = 'b000011101;
    x_28 = 'b000011111;
    x_29 = 'b000001110;
    x_30 = 'b000011001;
    x_31 = 'b000100001;
    x_32 = 'b000101000;
    x_33 = 'b000100110;
    x_34 = 'b000100101;
    x_35 = 'b000011011;
    x_36 = 'b000011010;
    x_37 = 'b000010100;
    x_38 = 'b000001100;
    x_39 = 'b000001110;
    x_40 = 'b000000110;
    x_41 = 'b000001100;
    x_42 = 'b000000100;
    x_43 = 'b111111011;
    x_44 = 'b000010001;
    x_45 = 'b000000100;
    x_46 = 'b000011101;
    x_47 = 'b000100100;
    x_48 = 'b000011101;
    x_49 = 'b000011111;
    x_50 = 'b000100101;
    x_51 = 'b000100101;
    x_52 = 'b000011101;
    x_53 = 'b000011010;
    x_54 = 'b000010011;
    x_55 = 'b000011010;
    x_56 = 'b000100100;
    x_57 = 'b000100011;
    x_58 = 'b000100101;
    x_59 = 'b000011010;
    x_60 = 'b000011000;
    x_61 = 'b000100001;
    x_62 = 'b000010010;
    x_63 = 'b000101010;

    h_0 = 'b000011100;
    h_1 = 'b000100110;
    h_2 = 'b000101001;
    h_3 = 'b000110001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000010011;
    x_1 = 'b000011111;
    x_2 = 'b000100100;
    x_3 = 'b000101100;
    x_4 = 'b000100101;
    x_5 = 'b000010111;
    x_6 = 'b000010101;
    x_7 = 'b000001011;
    x_8 = 'b000011101;
    x_9 = 'b000100101;
    x_10 = 'b000101000;
    x_11 = 'b000101111;
    x_12 = 'b000011110;
    x_13 = 'b000001101;
    x_14 = 'b000100000;
    x_15 = 'b000100111;
    x_16 = 'b000100111;
    x_17 = 'b000101001;
    x_18 = 'b000100111;
    x_19 = 'b000100100;
    x_20 = 'b000010101;
    x_21 = 'b000010011;
    x_22 = 'b000010000;
    x_23 = 'b000010010;
    x_24 = 'b000010010;
    x_25 = 'b000010011;
    x_26 = 'b000011010;
    x_27 = 'b000010011;
    x_28 = 'b000010011;
    x_29 = 'b000001100;
    x_30 = 'b000011101;
    x_31 = 'b000011110;
    x_32 = 'b000101000;
    x_33 = 'b000100101;
    x_34 = 'b000100001;
    x_35 = 'b000011010;
    x_36 = 'b000010100;
    x_37 = 'b000001101;
    x_38 = 'b000001011;
    x_39 = 'b000001001;
    x_40 = 'b000010001;
    x_41 = 'b000000101;
    x_42 = 'b000010101;
    x_43 = 'b000011011;
    x_44 = 'b000011010;
    x_45 = 'b000001010;
    x_46 = 'b000011001;
    x_47 = 'b000011101;
    x_48 = 'b000010101;
    x_49 = 'b000011100;
    x_50 = 'b000100101;
    x_51 = 'b000101001;
    x_52 = 'b000100100;
    x_53 = 'b000100101;
    x_54 = 'b000011011;
    x_55 = 'b000010001;
    x_56 = 'b000011100;
    x_57 = 'b000011111;
    x_58 = 'b000100111;
    x_59 = 'b000011001;
    x_60 = 'b000010100;
    x_61 = 'b000011011;
    x_62 = 'b000001011;
    x_63 = 'b000100011;

    h_0 = 'b000010011;
    h_1 = 'b000011111;
    h_2 = 'b000100100;
    h_3 = 'b000101100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000011001;
    x_1 = 'b000100101;
    x_2 = 'b000101100;
    x_3 = 'b000110101;
    x_4 = 'b000101111;
    x_5 = 'b000100010;
    x_6 = 'b000011100;
    x_7 = 'b000000110;
    x_8 = 'b000100000;
    x_9 = 'b000101011;
    x_10 = 'b000110001;
    x_11 = 'b000111010;
    x_12 = 'b000101111;
    x_13 = 'b000011100;
    x_14 = 'b000010011;
    x_15 = 'b000100101;
    x_16 = 'b000101000;
    x_17 = 'b000101010;
    x_18 = 'b000101110;
    x_19 = 'b000110010;
    x_20 = 'b000101001;
    x_21 = 'b000010001;
    x_22 = 'b000001111;
    x_23 = 'b000001111;
    x_24 = 'b000010110;
    x_25 = 'b000010111;
    x_26 = 'b000011101;
    x_27 = 'b000010110;
    x_28 = 'b000010010;
    x_29 = 'b000010001;
    x_30 = 'b000100100;
    x_31 = 'b000100011;
    x_32 = 'b000101010;
    x_33 = 'b000101010;
    x_34 = 'b000100110;
    x_35 = 'b000100000;
    x_36 = 'b000011101;
    x_37 = 'b000010100;
    x_38 = 'b000010011;
    x_39 = 'b000010011;
    x_40 = 'b000100000;
    x_41 = 'b000010011;
    x_42 = 'b000010101;
    x_43 = 'b001001010;
    x_44 = 'b000011001;
    x_45 = 'b000100001;
    x_46 = 'b000010011;
    x_47 = 'b000010101;
    x_48 = 'b000001101;
    x_49 = 'b000010100;
    x_50 = 'b000100011;
    x_51 = 'b000101101;
    x_52 = 'b000101111;
    x_53 = 'b000110011;
    x_54 = 'b000101111;
    x_55 = 'b000001001;
    x_56 = 'b000010101;
    x_57 = 'b000011011;
    x_58 = 'b000101101;
    x_59 = 'b000100000;
    x_60 = 'b000001110;
    x_61 = 'b000010100;
    x_62 = 'b000000111;
    x_63 = 'b000011000;

    h_0 = 'b000011001;
    h_1 = 'b000100101;
    h_2 = 'b000101100;
    h_3 = 'b000110101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000011001;
    x_1 = 'b000100011;
    x_2 = 'b000101001;
    x_3 = 'b000110101;
    x_4 = 'b000110001;
    x_5 = 'b000100111;
    x_6 = 'b000100110;
    x_7 = 'b000001001;
    x_8 = 'b000011100;
    x_9 = 'b000100101;
    x_10 = 'b000101110;
    x_11 = 'b000111010;
    x_12 = 'b000110011;
    x_13 = 'b000100111;
    x_14 = 'b000010011;
    x_15 = 'b000100000;
    x_16 = 'b000100010;
    x_17 = 'b000100110;
    x_18 = 'b000101110;
    x_19 = 'b000110100;
    x_20 = 'b000110000;
    x_21 = 'b000010110;
    x_22 = 'b000010010;
    x_23 = 'b000010101;
    x_24 = 'b000010110;
    x_25 = 'b000011000;
    x_26 = 'b000100001;
    x_27 = 'b000011011;
    x_28 = 'b000011000;
    x_29 = 'b000010001;
    x_30 = 'b000100001;
    x_31 = 'b000100110;
    x_32 = 'b000101011;
    x_33 = 'b000101001;
    x_34 = 'b000100111;
    x_35 = 'b000100001;
    x_36 = 'b000100011;
    x_37 = 'b000011100;
    x_38 = 'b000001101;
    x_39 = 'b000011000;
    x_40 = 'b000011000;
    x_41 = 'b000011001;
    x_42 = 'b000001110;
    x_43 = 'b000101010;
    x_44 = 'b000001110;
    x_45 = 'b000100100;
    x_46 = 'b000001101;
    x_47 = 'b000010010;
    x_48 = 'b000001011;
    x_49 = 'b000010011;
    x_50 = 'b000100001;
    x_51 = 'b000101100;
    x_52 = 'b000101011;
    x_53 = 'b000110001;
    x_54 = 'b000101010;
    x_55 = 'b000001001;
    x_56 = 'b000010100;
    x_57 = 'b000011010;
    x_58 = 'b000101000;
    x_59 = 'b000010111;
    x_60 = 'b000001001;
    x_61 = 'b000001110;
    x_62 = 'b000000011;
    x_63 = 'b000001100;

    h_0 = 'b000011001;
    h_1 = 'b000100011;
    h_2 = 'b000101001;
    h_3 = 'b000110101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000010111;
    x_1 = 'b000011110;
    x_2 = 'b000100110;
    x_3 = 'b000101111;
    x_4 = 'b000101011;
    x_5 = 'b000100100;
    x_6 = 'b000100110;
    x_7 = 'b000000110;
    x_8 = 'b000010101;
    x_9 = 'b000011101;
    x_10 = 'b000100101;
    x_11 = 'b000110100;
    x_12 = 'b000101100;
    x_13 = 'b000101001;
    x_14 = 'b000001110;
    x_15 = 'b000011000;
    x_16 = 'b000011011;
    x_17 = 'b000100001;
    x_18 = 'b000100111;
    x_19 = 'b000101100;
    x_20 = 'b000101000;
    x_21 = 'b000011011;
    x_22 = 'b000010011;
    x_23 = 'b000010110;
    x_24 = 'b000011001;
    x_25 = 'b000011011;
    x_26 = 'b000100001;
    x_27 = 'b000011010;
    x_28 = 'b000010010;
    x_29 = 'b000010011;
    x_30 = 'b000100001;
    x_31 = 'b000100010;
    x_32 = 'b000101001;
    x_33 = 'b000100110;
    x_34 = 'b000100011;
    x_35 = 'b000011111;
    x_36 = 'b000011001;
    x_37 = 'b000010111;
    x_38 = 'b000010000;
    x_39 = 'b000001110;
    x_40 = 'b000010111;
    x_41 = 'b000001101;
    x_42 = 'b000001110;
    x_43 = 'b000100101;
    x_44 = 'b000000011;
    x_45 = 'b000010000;
    x_46 = 'b000010010;
    x_47 = 'b000010110;
    x_48 = 'b000001100;
    x_49 = 'b000010101;
    x_50 = 'b000011110;
    x_51 = 'b000100110;
    x_52 = 'b000100010;
    x_53 = 'b000100011;
    x_54 = 'b000011111;
    x_55 = 'b000010101;
    x_56 = 'b000011101;
    x_57 = 'b000011110;
    x_58 = 'b000100011;
    x_59 = 'b000010010;
    x_60 = 'b000001101;
    x_61 = 'b000001110;
    x_62 = 'b000000001;
    x_63 = 'b000001011;

    h_0 = 'b000010111;
    h_1 = 'b000011110;
    h_2 = 'b000100110;
    h_3 = 'b000101111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000010001;
    x_1 = 'b000010011;
    x_2 = 'b000011010;
    x_3 = 'b000100010;
    x_4 = 'b000011111;
    x_5 = 'b000010011;
    x_6 = 'b000001110;
    x_7 = 'b000001000;
    x_8 = 'b000010000;
    x_9 = 'b000010100;
    x_10 = 'b000011010;
    x_11 = 'b000100101;
    x_12 = 'b000011010;
    x_13 = 'b000001001;
    x_14 = 'b000010011;
    x_15 = 'b000011010;
    x_16 = 'b000011001;
    x_17 = 'b000011010;
    x_18 = 'b000011011;
    x_19 = 'b000011100;
    x_20 = 'b000010011;
    x_21 = 'b000010100;
    x_22 = 'b000001100;
    x_23 = 'b000001111;
    x_24 = 'b000001101;
    x_25 = 'b000001111;
    x_26 = 'b000010011;
    x_27 = 'b000001101;
    x_28 = 'b000010001;
    x_29 = 'b000000111;
    x_30 = 'b000010011;
    x_31 = 'b000001111;
    x_32 = 'b000010110;
    x_33 = 'b000010011;
    x_34 = 'b000010000;
    x_35 = 'b000001001;
    x_36 = 'b000000010;
    x_37 = 'b000001001;
    x_38 = 'b000000111;
    x_39 = 'b111111010;
    x_40 = 'b000001001;
    x_41 = 'b111111101;
    x_42 = 'b000001100;
    x_43 = 'b000100011;
    x_44 = 'b000011000;
    x_45 = 'b000010011;
    x_46 = 'b000101010;
    x_47 = 'b000100010;
    x_48 = 'b000010011;
    x_49 = 'b000011011;
    x_50 = 'b000011101;
    x_51 = 'b000011111;
    x_52 = 'b000011001;
    x_53 = 'b000011100;
    x_54 = 'b000011100;
    x_55 = 'b000100011;
    x_56 = 'b000101010;
    x_57 = 'b000100010;
    x_58 = 'b000100001;
    x_59 = 'b000010101;
    x_60 = 'b000011000;
    x_61 = 'b000011001;
    x_62 = 'b000000110;
    x_63 = 'b000011001;

    h_0 = 'b000010001;
    h_1 = 'b000010011;
    h_2 = 'b000011010;
    h_3 = 'b000100010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000000110;
    x_1 = 'b000000111;
    x_2 = 'b000001011;
    x_3 = 'b000010001;
    x_4 = 'b000001101;
    x_5 = 'b000000000;
    x_6 = 'b111111100;
    x_7 = 'b111111111;
    x_8 = 'b000001100;
    x_9 = 'b000001111;
    x_10 = 'b000010001;
    x_11 = 'b000010010;
    x_12 = 'b000001011;
    x_13 = 'b111111100;
    x_14 = 'b000011000;
    x_15 = 'b000011100;
    x_16 = 'b000011000;
    x_17 = 'b000010111;
    x_18 = 'b000010001;
    x_19 = 'b000010001;
    x_20 = 'b000001011;
    x_21 = 'b000000111;
    x_22 = 'b000000010;
    x_23 = 'b000000110;
    x_24 = 'b000000111;
    x_25 = 'b000001000;
    x_26 = 'b000000100;
    x_27 = 'b111111110;
    x_28 = 'b000000111;
    x_29 = 'b000000011;
    x_30 = 'b000001111;
    x_31 = 'b000000110;
    x_32 = 'b000001101;
    x_33 = 'b000001000;
    x_34 = 'b000000011;
    x_35 = 'b111111110;
    x_36 = 'b111110110;
    x_37 = 'b000000000;
    x_38 = 'b000001110;
    x_39 = 'b111110011;
    x_40 = 'b000011110;
    x_41 = 'b000010010;
    x_42 = 'b000100001;
    x_43 = 'b000000110;
    x_44 = 'b000100111;
    x_45 = 'b000001111;
    x_46 = 'b000101101;
    x_47 = 'b000101001;
    x_48 = 'b000010111;
    x_49 = 'b000011111;
    x_50 = 'b000011100;
    x_51 = 'b000011011;
    x_52 = 'b000010100;
    x_53 = 'b000011000;
    x_54 = 'b000011010;
    x_55 = 'b000101011;
    x_56 = 'b000110000;
    x_57 = 'b000100110;
    x_58 = 'b000011110;
    x_59 = 'b000010110;
    x_60 = 'b000100110;
    x_61 = 'b000100101;
    x_62 = 'b000001100;
    x_63 = 'b000101010;

    h_0 = 'b000000110;
    h_1 = 'b000000111;
    h_2 = 'b000001011;
    h_3 = 'b000010001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000010101;
    x_1 = 'b000010000;
    x_2 = 'b000010000;
    x_3 = 'b000010001;
    x_4 = 'b000001101;
    x_5 = 'b111111101;
    x_6 = 'b111111011;
    x_7 = 'b000001101;
    x_8 = 'b000010100;
    x_9 = 'b000010001;
    x_10 = 'b000001110;
    x_11 = 'b000001111;
    x_12 = 'b000000110;
    x_13 = 'b111111011;
    x_14 = 'b000100000;
    x_15 = 'b000011111;
    x_16 = 'b000011000;
    x_17 = 'b000010001;
    x_18 = 'b000001011;
    x_19 = 'b000001100;
    x_20 = 'b000000110;
    x_21 = 'b000001011;
    x_22 = 'b000000100;
    x_23 = 'b000000100;
    x_24 = 'b000001100;
    x_25 = 'b000001101;
    x_26 = 'b000000110;
    x_27 = 'b111111111;
    x_28 = 'b000000100;
    x_29 = 'b000010000;
    x_30 = 'b000010001;
    x_31 = 'b000000111;
    x_32 = 'b000010010;
    x_33 = 'b000001110;
    x_34 = 'b000001000;
    x_35 = 'b000000011;
    x_36 = 'b111111000;
    x_37 = 'b000000010;
    x_38 = 'b000010011;
    x_39 = 'b111101110;
    x_40 = 'b000100110;
    x_41 = 'b111111000;
    x_42 = 'b000101101;
    x_43 = 'b111101010;
    x_44 = 'b000101000;
    x_45 = 'b000000000;
    x_46 = 'b000101010;
    x_47 = 'b000101001;
    x_48 = 'b000010111;
    x_49 = 'b000011011;
    x_50 = 'b000010110;
    x_51 = 'b000010100;
    x_52 = 'b000001011;
    x_53 = 'b000001110;
    x_54 = 'b000001100;
    x_55 = 'b000101010;
    x_56 = 'b000101110;
    x_57 = 'b000100011;
    x_58 = 'b000010110;
    x_59 = 'b000001010;
    x_60 = 'b000101011;
    x_61 = 'b000101000;
    x_62 = 'b000001100;
    x_63 = 'b000101111;

    h_0 = 'b000010101;
    h_1 = 'b000010000;
    h_2 = 'b000010000;
    h_3 = 'b000010001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000010101;
    x_1 = 'b000010010;
    x_2 = 'b000010001;
    x_3 = 'b000010010;
    x_4 = 'b000001010;
    x_5 = 'b111111001;
    x_6 = 'b111111000;
    x_7 = 'b000010000;
    x_8 = 'b000010010;
    x_9 = 'b000001110;
    x_10 = 'b000001101;
    x_11 = 'b000001101;
    x_12 = 'b000000000;
    x_13 = 'b111110010;
    x_14 = 'b000100000;
    x_15 = 'b000011100;
    x_16 = 'b000010100;
    x_17 = 'b000001100;
    x_18 = 'b000001001;
    x_19 = 'b000001001;
    x_20 = 'b000000000;
    x_21 = 'b000001100;
    x_22 = 'b000000001;
    x_23 = 'b000000010;
    x_24 = 'b000001111;
    x_25 = 'b000010000;
    x_26 = 'b000000100;
    x_27 = 'b111111110;
    x_28 = 'b000000100;
    x_29 = 'b000010110;
    x_30 = 'b000001011;
    x_31 = 'b000000110;
    x_32 = 'b000001111;
    x_33 = 'b000001001;
    x_34 = 'b000000011;
    x_35 = 'b111111100;
    x_36 = 'b111110111;
    x_37 = 'b000000010;
    x_38 = 'b000011000;
    x_39 = 'b111100111;
    x_40 = 'b000101011;
    x_41 = 'b111100010;
    x_42 = 'b000100110;
    x_43 = 'b000110000;
    x_44 = 'b000100111;
    x_45 = 'b111111101;
    x_46 = 'b000100101;
    x_47 = 'b000100010;
    x_48 = 'b000010010;
    x_49 = 'b000011000;
    x_50 = 'b000010101;
    x_51 = 'b000010011;
    x_52 = 'b000001010;
    x_53 = 'b000001011;
    x_54 = 'b000000100;
    x_55 = 'b000011101;
    x_56 = 'b000100100;
    x_57 = 'b000011100;
    x_58 = 'b000010000;
    x_59 = 'b000000010;
    x_60 = 'b000100100;
    x_61 = 'b000100001;
    x_62 = 'b000000100;
    x_63 = 'b000100000;

    h_0 = 'b000010101;
    h_1 = 'b000010010;
    h_2 = 'b000010001;
    h_3 = 'b000010010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000001111;
    x_1 = 'b000000110;
    x_2 = 'b000001000;
    x_3 = 'b000001101;
    x_4 = 'b111111110;
    x_5 = 'b111101101;
    x_6 = 'b111101110;
    x_7 = 'b000000001;
    x_8 = 'b000000111;
    x_9 = 'b000000110;
    x_10 = 'b000001000;
    x_11 = 'b000000100;
    x_12 = 'b111110101;
    x_13 = 'b111101100;
    x_14 = 'b000001111;
    x_15 = 'b000001111;
    x_16 = 'b000001001;
    x_17 = 'b000000101;
    x_18 = 'b000000010;
    x_19 = 'b000000001;
    x_20 = 'b111110111;
    x_21 = 'b000000111;
    x_22 = 'b111110101;
    x_23 = 'b111110111;
    x_24 = 'b000001011;
    x_25 = 'b000001100;
    x_26 = 'b111110100;
    x_27 = 'b111101110;
    x_28 = 'b111110111;
    x_29 = 'b000001110;
    x_30 = 'b000000101;
    x_31 = 'b111111001;
    x_32 = 'b000000100;
    x_33 = 'b111111001;
    x_34 = 'b111110010;
    x_35 = 'b111101111;
    x_36 = 'b111100101;
    x_37 = 'b111110101;
    x_38 = 'b000010110;
    x_39 = 'b111011010;
    x_40 = 'b000100100;
    x_41 = 'b111101001;
    x_42 = 'b000001100;
    x_43 = 'b000101011;
    x_44 = 'b000010000;
    x_45 = 'b111011001;
    x_46 = 'b000001110;
    x_47 = 'b000001111;
    x_48 = 'b000000010;
    x_49 = 'b000001001;
    x_50 = 'b000000111;
    x_51 = 'b000000101;
    x_52 = 'b111111011;
    x_53 = 'b111111000;
    x_54 = 'b111101011;
    x_55 = 'b000001100;
    x_56 = 'b000010011;
    x_57 = 'b000001111;
    x_58 = 'b000000010;
    x_59 = 'b111110110;
    x_60 = 'b000010101;
    x_61 = 'b000010000;
    x_62 = 'b111110100;
    x_63 = 'b000001000;

    h_0 = 'b000001111;
    h_1 = 'b000000110;
    h_2 = 'b000001000;
    h_3 = 'b000001101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000010100;
    x_1 = 'b000001011;
    x_2 = 'b000001011;
    x_3 = 'b000001110;
    x_4 = 'b000000001;
    x_5 = 'b111101110;
    x_6 = 'b111100111;
    x_7 = 'b000001101;
    x_8 = 'b000010000;
    x_9 = 'b000010001;
    x_10 = 'b000010011;
    x_11 = 'b000010001;
    x_12 = 'b111111101;
    x_13 = 'b111110000;
    x_14 = 'b000010101;
    x_15 = 'b000011001;
    x_16 = 'b000010011;
    x_17 = 'b000010001;
    x_18 = 'b000010000;
    x_19 = 'b000001110;
    x_20 = 'b111111111;
    x_21 = 'b000000011;
    x_22 = 'b111110111;
    x_23 = 'b111111011;
    x_24 = 'b000001001;
    x_25 = 'b000001011;
    x_26 = 'b111111101;
    x_27 = 'b111110011;
    x_28 = 'b111111011;
    x_29 = 'b000001111;
    x_30 = 'b000000111;
    x_31 = 'b000000100;
    x_32 = 'b000010010;
    x_33 = 'b000001011;
    x_34 = 'b000000010;
    x_35 = 'b111111110;
    x_36 = 'b111110010;
    x_37 = 'b000000110;
    x_38 = 'b000011100;
    x_39 = 'b111110000;
    x_40 = 'b000100000;
    x_41 = 'b000001100;
    x_42 = 'b000011001;
    x_43 = 'b000011011;
    x_44 = 'b000010111;
    x_45 = 'b000001100;
    x_46 = 'b000011001;
    x_47 = 'b000011101;
    x_48 = 'b000010001;
    x_49 = 'b000011010;
    x_50 = 'b000011011;
    x_51 = 'b000011001;
    x_52 = 'b000010001;
    x_53 = 'b000010000;
    x_54 = 'b000001101;
    x_55 = 'b000011000;
    x_56 = 'b000100001;
    x_57 = 'b000011101;
    x_58 = 'b000010010;
    x_59 = 'b000000101;
    x_60 = 'b000010001;
    x_61 = 'b000001111;
    x_62 = 'b111110011;
    x_63 = 'b000001000;

    h_0 = 'b000010100;
    h_1 = 'b000001011;
    h_2 = 'b000001011;
    h_3 = 'b000001110;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000011010;
    x_1 = 'b000011001;
    x_2 = 'b000011100;
    x_3 = 'b000100000;
    x_4 = 'b000011001;
    x_5 = 'b000000101;
    x_6 = 'b111111101;
    x_7 = 'b000010111;
    x_8 = 'b000011101;
    x_9 = 'b000011110;
    x_10 = 'b000100011;
    x_11 = 'b000100100;
    x_12 = 'b000010111;
    x_13 = 'b000001001;
    x_14 = 'b000100101;
    x_15 = 'b000100100;
    x_16 = 'b000100011;
    x_17 = 'b000100001;
    x_18 = 'b000100001;
    x_19 = 'b000100000;
    x_20 = 'b000010011;
    x_21 = 'b000001000;
    x_22 = 'b000000001;
    x_23 = 'b000000010;
    x_24 = 'b000001001;
    x_25 = 'b000001100;
    x_26 = 'b000001000;
    x_27 = 'b111111100;
    x_28 = 'b000000000;
    x_29 = 'b000001110;
    x_30 = 'b000000111;
    x_31 = 'b000001011;
    x_32 = 'b000010110;
    x_33 = 'b000010000;
    x_34 = 'b000001010;
    x_35 = 'b000000010;
    x_36 = 'b111111000;
    x_37 = 'b000001011;
    x_38 = 'b000001101;
    x_39 = 'b111111000;
    x_40 = 'b000001111;
    x_41 = 'b000001100;
    x_42 = 'b000011001;
    x_43 = 'b000011110;
    x_44 = 'b000010101;
    x_45 = 'b000010101;
    x_46 = 'b000011111;
    x_47 = 'b000100010;
    x_48 = 'b000010010;
    x_49 = 'b000011110;
    x_50 = 'b000011110;
    x_51 = 'b000011101;
    x_52 = 'b000010111;
    x_53 = 'b000010011;
    x_54 = 'b000001010;
    x_55 = 'b000011101;
    x_56 = 'b000100101;
    x_57 = 'b000100000;
    x_58 = 'b000010110;
    x_59 = 'b000000110;
    x_60 = 'b000011001;
    x_61 = 'b000011001;
    x_62 = 'b111111111;
    x_63 = 'b000010101;

    h_0 = 'b000011010;
    h_1 = 'b000011001;
    h_2 = 'b000011100;
    h_3 = 'b000100000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000000101;
    x_1 = 'b000000111;
    x_2 = 'b111101000;
    x_3 = 'b111110000;
    x_4 = 'b111101101;
    x_5 = 'b111101001;
    x_6 = 'b111110100;
    x_7 = 'b000010001;
    x_8 = 'b000000001;
    x_9 = 'b111110100;
    x_10 = 'b111101100;
    x_11 = 'b111011111;
    x_12 = 'b111100010;
    x_13 = 'b111100110;
    x_14 = 'b000011000;
    x_15 = 'b000001001;
    x_16 = 'b111111000;
    x_17 = 'b111110000;
    x_18 = 'b111011111;
    x_19 = 'b111100000;
    x_20 = 'b111101010;
    x_21 = 'b111111111;
    x_22 = 'b000001000;
    x_23 = 'b000001010;
    x_24 = 'b000000110;
    x_25 = 'b000000101;
    x_26 = 'b111110001;
    x_27 = 'b111111000;
    x_28 = 'b000001111;
    x_29 = 'b000000011;
    x_30 = 'b000010010;
    x_31 = 'b111111110;
    x_32 = 'b111111001;
    x_33 = 'b111110101;
    x_34 = 'b111110011;
    x_35 = 'b111101110;
    x_36 = 'b111111110;
    x_37 = 'b111011001;
    x_38 = 'b000001001;
    x_39 = 'b000000100;
    x_40 = 'b000010001;
    x_41 = 'b000000111;
    x_42 = 'b000011000;
    x_43 = 'b111111110;
    x_44 = 'b000011100;
    x_45 = 'b000000000;
    x_46 = 'b000011011;
    x_47 = 'b000010110;
    x_48 = 'b000001110;
    x_49 = 'b000000101;
    x_50 = 'b111110101;
    x_51 = 'b111101111;
    x_52 = 'b111110001;
    x_53 = 'b111110111;
    x_54 = 'b000001010;
    x_55 = 'b000001110;
    x_56 = 'b000010101;
    x_57 = 'b111111010;
    x_58 = 'b111111001;
    x_59 = 'b000010101;
    x_60 = 'b000000011;
    x_61 = 'b111111010;
    x_62 = 'b111111101;
    x_63 = 'b000001000;

    h_0 = 'b000000101;
    h_1 = 'b000000111;
    h_2 = 'b111101000;
    h_3 = 'b111110000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000010101;
    x_1 = 'b000011000;
    x_2 = 'b000000000;
    x_3 = 'b000000101;
    x_4 = 'b111111101;
    x_5 = 'b111111001;
    x_6 = 'b111111110;
    x_7 = 'b000100110;
    x_8 = 'b000010010;
    x_9 = 'b000000111;
    x_10 = 'b000000000;
    x_11 = 'b111110110;
    x_12 = 'b111111000;
    x_13 = 'b111111011;
    x_14 = 'b000011000;
    x_15 = 'b000010100;
    x_16 = 'b000001000;
    x_17 = 'b000000110;
    x_18 = 'b111110110;
    x_19 = 'b111111010;
    x_20 = 'b000000000;
    x_21 = 'b000000001;
    x_22 = 'b000001010;
    x_23 = 'b000001101;
    x_24 = 'b000001011;
    x_25 = 'b000001011;
    x_26 = 'b111111100;
    x_27 = 'b111111111;
    x_28 = 'b000010000;
    x_29 = 'b000001111;
    x_30 = 'b000011110;
    x_31 = 'b000001000;
    x_32 = 'b000001001;
    x_33 = 'b000000010;
    x_34 = 'b111111101;
    x_35 = 'b111111011;
    x_36 = 'b000000010;
    x_37 = 'b111010101;
    x_38 = 'b000011101;
    x_39 = 'b000000110;
    x_40 = 'b000100111;
    x_41 = 'b111110011;
    x_42 = 'b000011001;
    x_43 = 'b000010100;
    x_44 = 'b000011100;
    x_45 = 'b000001010;
    x_46 = 'b000010000;
    x_47 = 'b000010011;
    x_48 = 'b000001110;
    x_49 = 'b000001001;
    x_50 = 'b000000010;
    x_51 = 'b000000001;
    x_52 = 'b000000010;
    x_53 = 'b000000100;
    x_54 = 'b000010010;
    x_55 = 'b000001001;
    x_56 = 'b000001111;
    x_57 = 'b000000000;
    x_58 = 'b000001010;
    x_59 = 'b000010110;
    x_60 = 'b111111100;
    x_61 = 'b111111101;
    x_62 = 'b000001001;
    x_63 = 'b111110111;

    h_0 = 'b000010101;
    h_1 = 'b000011000;
    h_2 = 'b000000000;
    h_3 = 'b000000101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000100101;
    x_1 = 'b000100001;
    x_2 = 'b000001010;
    x_3 = 'b000001011;
    x_4 = 'b000000001;
    x_5 = 'b111111101;
    x_6 = 'b111111101;
    x_7 = 'b000101010;
    x_8 = 'b000010100;
    x_9 = 'b000001100;
    x_10 = 'b000000100;
    x_11 = 'b000000001;
    x_12 = 'b000000010;
    x_13 = 'b111111011;
    x_14 = 'b000011100;
    x_15 = 'b000010110;
    x_16 = 'b000001011;
    x_17 = 'b000001101;
    x_18 = 'b000000101;
    x_19 = 'b000001011;
    x_20 = 'b000001110;
    x_21 = 'b000010100;
    x_22 = 'b000011001;
    x_23 = 'b000010110;
    x_24 = 'b000100100;
    x_25 = 'b000100010;
    x_26 = 'b000001000;
    x_27 = 'b000000110;
    x_28 = 'b000010011;
    x_29 = 'b000101000;
    x_30 = 'b000110111;
    x_31 = 'b000010101;
    x_32 = 'b000011000;
    x_33 = 'b000001111;
    x_34 = 'b000001001;
    x_35 = 'b000000110;
    x_36 = 'b000000011;
    x_37 = 'b111001110;
    x_38 = 'b000111001;
    x_39 = 'b111111110;
    x_40 = 'b000110111;
    x_41 = 'b111100001;
    x_42 = 'b000101110;
    x_43 = 'b000000001;
    x_44 = 'b000101001;
    x_45 = 'b000101010;
    x_46 = 'b000011110;
    x_47 = 'b000100000;
    x_48 = 'b000100000;
    x_49 = 'b000011011;
    x_50 = 'b000011100;
    x_51 = 'b000100011;
    x_52 = 'b000101000;
    x_53 = 'b000101001;
    x_54 = 'b000110000;
    x_55 = 'b000010111;
    x_56 = 'b000011101;
    x_57 = 'b000011100;
    x_58 = 'b000110000;
    x_59 = 'b000101110;
    x_60 = 'b111111100;
    x_61 = 'b000000100;
    x_62 = 'b000010000;
    x_63 = 'b111101000;

    h_0 = 'b000100101;
    h_1 = 'b000100001;
    h_2 = 'b000001010;
    h_3 = 'b000001011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000111001;
    x_1 = 'b000110110;
    x_2 = 'b000011111;
    x_3 = 'b000011100;
    x_4 = 'b000010111;
    x_5 = 'b000010110;
    x_6 = 'b000010000;
    x_7 = 'b000111011;
    x_8 = 'b000101010;
    x_9 = 'b000100101;
    x_10 = 'b000100001;
    x_11 = 'b000011101;
    x_12 = 'b000100110;
    x_13 = 'b000100000;
    x_14 = 'b000110001;
    x_15 = 'b000101111;
    x_16 = 'b000100101;
    x_17 = 'b000100111;
    x_18 = 'b000101010;
    x_19 = 'b000110011;
    x_20 = 'b000111001;
    x_21 = 'b000011000;
    x_22 = 'b000011001;
    x_23 = 'b000010110;
    x_24 = 'b000100011;
    x_25 = 'b000100011;
    x_26 = 'b000010000;
    x_27 = 'b000001011;
    x_28 = 'b000010100;
    x_29 = 'b000011111;
    x_30 = 'b000111000;
    x_31 = 'b000011001;
    x_32 = 'b000011010;
    x_33 = 'b000010100;
    x_34 = 'b000001111;
    x_35 = 'b000001011;
    x_36 = 'b000001011;
    x_37 = 'b111010110;
    x_38 = 'b000101101;
    x_39 = 'b000010011;
    x_40 = 'b000101101;
    x_41 = 'b000001110;
    x_42 = 'b000101001;
    x_43 = 'b111111110;
    x_44 = 'b000101100;
    x_45 = 'b001000011;
    x_46 = 'b000100110;
    x_47 = 'b000100100;
    x_48 = 'b000100011;
    x_49 = 'b000100011;
    x_50 = 'b000100110;
    x_51 = 'b000111000;
    x_52 = 'b000111101;
    x_53 = 'b000111110;
    x_54 = 'b001000000;
    x_55 = 'b000011001;
    x_56 = 'b000011100;
    x_57 = 'b000100111;
    x_58 = 'b001000100;
    x_59 = 'b000111010;
    x_60 = 'b000000100;
    x_61 = 'b000010101;
    x_62 = 'b000100001;
    x_63 = 'b111110100;

    h_0 = 'b000111001;
    h_1 = 'b000110110;
    h_2 = 'b000011111;
    h_3 = 'b000011100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000010111;
    x_1 = 'b000011001;
    x_2 = 'b000001000;
    x_3 = 'b000001001;
    x_4 = 'b000001101;
    x_5 = 'b000010000;
    x_6 = 'b000010101;
    x_7 = 'b000011010;
    x_8 = 'b000010000;
    x_9 = 'b000001110;
    x_10 = 'b000001110;
    x_11 = 'b000010000;
    x_12 = 'b000100100;
    x_13 = 'b000100110;
    x_14 = 'b000011000;
    x_15 = 'b000010111;
    x_16 = 'b000010010;
    x_17 = 'b000010111;
    x_18 = 'b000011101;
    x_19 = 'b000101011;
    x_20 = 'b000110110;
    x_21 = 'b111110111;
    x_22 = 'b000000001;
    x_23 = 'b000001011;
    x_24 = 'b111111010;
    x_25 = 'b111111010;
    x_26 = 'b111111001;
    x_27 = 'b000000001;
    x_28 = 'b000001101;
    x_29 = 'b111110110;
    x_30 = 'b000001001;
    x_31 = 'b000000111;
    x_32 = 'b111111011;
    x_33 = 'b111111011;
    x_34 = 'b111111110;
    x_35 = 'b111110111;
    x_36 = 'b000001011;
    x_37 = 'b111011100;
    x_38 = 'b111111101;
    x_39 = 'b000011000;
    x_40 = 'b000010011;
    x_41 = 'b000010111;
    x_42 = 'b000000100;
    x_43 = 'b000100111;
    x_44 = 'b000010001;
    x_45 = 'b000110001;
    x_46 = 'b000010010;
    x_47 = 'b000010010;
    x_48 = 'b000010001;
    x_49 = 'b000010011;
    x_50 = 'b000011011;
    x_51 = 'b000101101;
    x_52 = 'b000110000;
    x_53 = 'b000110001;
    x_54 = 'b000101010;
    x_55 = 'b000001111;
    x_56 = 'b000010011;
    x_57 = 'b000100001;
    x_58 = 'b000111001;
    x_59 = 'b000101110;
    x_60 = 'b000000111;
    x_61 = 'b000100010;
    x_62 = 'b000101101;
    x_63 = 'b000000011;

    h_0 = 'b000010111;
    h_1 = 'b000011001;
    h_2 = 'b000001000;
    h_3 = 'b000001001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000000110;
    x_1 = 'b000001011;
    x_2 = 'b111111101;
    x_3 = 'b000000010;
    x_4 = 'b000001001;
    x_5 = 'b000001110;
    x_6 = 'b000010101;
    x_7 = 'b000010110;
    x_8 = 'b000000111;
    x_9 = 'b000001000;
    x_10 = 'b000001011;
    x_11 = 'b000010000;
    x_12 = 'b000011111;
    x_13 = 'b000100111;
    x_14 = 'b000010110;
    x_15 = 'b000010011;
    x_16 = 'b000001110;
    x_17 = 'b000010101;
    x_18 = 'b000011001;
    x_19 = 'b000100100;
    x_20 = 'b000110001;
    x_21 = 'b000000011;
    x_22 = 'b000001010;
    x_23 = 'b000001110;
    x_24 = 'b000001101;
    x_25 = 'b000001011;
    x_26 = 'b111111110;
    x_27 = 'b000000100;
    x_28 = 'b000010001;
    x_29 = 'b000010000;
    x_30 = 'b000011111;
    x_31 = 'b000001110;
    x_32 = 'b000000101;
    x_33 = 'b000000100;
    x_34 = 'b000000011;
    x_35 = 'b000000000;
    x_36 = 'b000001101;
    x_37 = 'b111010100;
    x_38 = 'b000100001;
    x_39 = 'b000010000;
    x_40 = 'b000011100;
    x_41 = 'b000010000;
    x_42 = 'b000101111;
    x_43 = 'b111111110;
    x_44 = 'b000011110;
    x_45 = 'b000100011;
    x_46 = 'b000100100;
    x_47 = 'b000100100;
    x_48 = 'b000011111;
    x_49 = 'b000011111;
    x_50 = 'b000100010;
    x_51 = 'b000101111;
    x_52 = 'b000110000;
    x_53 = 'b000101101;
    x_54 = 'b000100111;
    x_55 = 'b000100101;
    x_56 = 'b000100111;
    x_57 = 'b000101011;
    x_58 = 'b000111010;
    x_59 = 'b000101110;
    x_60 = 'b000010001;
    x_61 = 'b000101100;
    x_62 = 'b000110010;
    x_63 = 'b000011010;

    h_0 = 'b000000110;
    h_1 = 'b000001011;
    h_2 = 'b111111101;
    h_3 = 'b000000010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000100110;
    x_1 = 'b000100001;
    x_2 = 'b000001011;
    x_3 = 'b000010001;
    x_4 = 'b000001101;
    x_5 = 'b000001110;
    x_6 = 'b000010100;
    x_7 = 'b000110110;
    x_8 = 'b000011101;
    x_9 = 'b000010110;
    x_10 = 'b000010101;
    x_11 = 'b000010011;
    x_12 = 'b000011001;
    x_13 = 'b000011100;
    x_14 = 'b000110001;
    x_15 = 'b000100100;
    x_16 = 'b000011100;
    x_17 = 'b000011101;
    x_18 = 'b000011011;
    x_19 = 'b000100010;
    x_20 = 'b000101001;
    x_21 = 'b000001110;
    x_22 = 'b000010101;
    x_23 = 'b000010111;
    x_24 = 'b000010111;
    x_25 = 'b000010111;
    x_26 = 'b000000011;
    x_27 = 'b000001010;
    x_28 = 'b000011110;
    x_29 = 'b000011010;
    x_30 = 'b000100111;
    x_31 = 'b000001100;
    x_32 = 'b000001001;
    x_33 = 'b000000110;
    x_34 = 'b000000011;
    x_35 = 'b111111111;
    x_36 = 'b000001100;
    x_37 = 'b111011111;
    x_38 = 'b000100001;
    x_39 = 'b000010010;
    x_40 = 'b000100111;
    x_41 = 'b000000110;
    x_42 = 'b000101110;
    x_43 = 'b000001100;
    x_44 = 'b000110110;
    x_45 = 'b000011010;
    x_46 = 'b000110100;
    x_47 = 'b000101011;
    x_48 = 'b000100010;
    x_49 = 'b000011111;
    x_50 = 'b000011111;
    x_51 = 'b000101001;
    x_52 = 'b000100111;
    x_53 = 'b000100101;
    x_54 = 'b000100101;
    x_55 = 'b000100111;
    x_56 = 'b000100101;
    x_57 = 'b000100101;
    x_58 = 'b000110100;
    x_59 = 'b000101100;
    x_60 = 'b000011011;
    x_61 = 'b000110011;
    x_62 = 'b000110010;
    x_63 = 'b000101010;

    h_0 = 'b000100110;
    h_1 = 'b000100001;
    h_2 = 'b000001011;
    h_3 = 'b000010001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000001001;
    x_1 = 'b000001110;
    x_2 = 'b111111111;
    x_3 = 'b000000111;
    x_4 = 'b111111111;
    x_5 = 'b111111100;
    x_6 = 'b000000011;
    x_7 = 'b000011010;
    x_8 = 'b000001011;
    x_9 = 'b000001100;
    x_10 = 'b000001100;
    x_11 = 'b000000001;
    x_12 = 'b000001000;
    x_13 = 'b000000011;
    x_14 = 'b000100100;
    x_15 = 'b000011000;
    x_16 = 'b000010010;
    x_17 = 'b000010101;
    x_18 = 'b000001111;
    x_19 = 'b000010101;
    x_20 = 'b000011000;
    x_21 = 'b111110101;
    x_22 = 'b111111110;
    x_23 = 'b000000101;
    x_24 = 'b111111010;
    x_25 = 'b111111010;
    x_26 = 'b111101111;
    x_27 = 'b111110101;
    x_28 = 'b000001010;
    x_29 = 'b111111000;
    x_30 = 'b000001101;
    x_31 = 'b111111100;
    x_32 = 'b111111010;
    x_33 = 'b111110110;
    x_34 = 'b111110010;
    x_35 = 'b111101011;
    x_36 = 'b111110100;
    x_37 = 'b111010101;
    x_38 = 'b111111111;
    x_39 = 'b111111011;
    x_40 = 'b000101010;
    x_41 = 'b111011101;
    x_42 = 'b000101001;
    x_43 = 'b000010001;
    x_44 = 'b000110110;
    x_45 = 'b000100100;
    x_46 = 'b000110001;
    x_47 = 'b000100111;
    x_48 = 'b000100001;
    x_49 = 'b000011110;
    x_50 = 'b000011100;
    x_51 = 'b000101000;
    x_52 = 'b000100111;
    x_53 = 'b000100110;
    x_54 = 'b000101101;
    x_55 = 'b000011111;
    x_56 = 'b000100001;
    x_57 = 'b000100011;
    x_58 = 'b000110110;
    x_59 = 'b000110011;
    x_60 = 'b000011011;
    x_61 = 'b000110011;
    x_62 = 'b000110000;
    x_63 = 'b000101001;

    h_0 = 'b000001001;
    h_1 = 'b000001110;
    h_2 = 'b111111111;
    h_3 = 'b000000111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000001001;
    x_1 = 'b000010010;
    x_2 = 'b000000100;
    x_3 = 'b000001010;
    x_4 = 'b000000000;
    x_5 = 'b111111001;
    x_6 = 'b111110101;
    x_7 = 'b000101010;
    x_8 = 'b000010110;
    x_9 = 'b000010110;
    x_10 = 'b000010100;
    x_11 = 'b000001010;
    x_12 = 'b000001011;
    x_13 = 'b111111111;
    x_14 = 'b000110001;
    x_15 = 'b000100111;
    x_16 = 'b000011100;
    x_17 = 'b000011111;
    x_18 = 'b000010110;
    x_19 = 'b000011001;
    x_20 = 'b000011101;
    x_21 = 'b111111110;
    x_22 = 'b000000001;
    x_23 = 'b000000101;
    x_24 = 'b000000111;
    x_25 = 'b000000101;
    x_26 = 'b111110111;
    x_27 = 'b111110110;
    x_28 = 'b000000100;
    x_29 = 'b000000000;
    x_30 = 'b000011000;
    x_31 = 'b000000100;
    x_32 = 'b000001000;
    x_33 = 'b000000100;
    x_34 = 'b111111011;
    x_35 = 'b111110111;
    x_36 = 'b111110111;
    x_37 = 'b111010100;
    x_38 = 'b000001011;
    x_39 = 'b111110111;
    x_40 = 'b000010011;
    x_41 = 'b111100100;
    x_42 = 'b000011110;
    x_43 = 'b000010100;
    x_44 = 'b000100011;
    x_45 = 'b000101001;
    x_46 = 'b000101011;
    x_47 = 'b000101011;
    x_48 = 'b000100111;
    x_49 = 'b000100101;
    x_50 = 'b000100100;
    x_51 = 'b000101010;
    x_52 = 'b000101001;
    x_53 = 'b000100111;
    x_54 = 'b000101010;
    x_55 = 'b000100011;
    x_56 = 'b000100011;
    x_57 = 'b000100011;
    x_58 = 'b000110100;
    x_59 = 'b000101110;
    x_60 = 'b000011001;
    x_61 = 'b000110000;
    x_62 = 'b000101100;
    x_63 = 'b000100011;

    h_0 = 'b000001001;
    h_1 = 'b000010010;
    h_2 = 'b000000100;
    h_3 = 'b000001010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000001010;
    x_1 = 'b000011001;
    x_2 = 'b000001110;
    x_3 = 'b000010110;
    x_4 = 'b000001010;
    x_5 = 'b000000110;
    x_6 = 'b000000011;
    x_7 = 'b000100001;
    x_8 = 'b000010111;
    x_9 = 'b000010111;
    x_10 = 'b000010101;
    x_11 = 'b000001111;
    x_12 = 'b000010001;
    x_13 = 'b000000110;
    x_14 = 'b000100000;
    x_15 = 'b000011011;
    x_16 = 'b000010110;
    x_17 = 'b000011100;
    x_18 = 'b000010100;
    x_19 = 'b000010110;
    x_20 = 'b000011010;
    x_21 = 'b111111000;
    x_22 = 'b111111111;
    x_23 = 'b000000100;
    x_24 = 'b111111100;
    x_25 = 'b111111101;
    x_26 = 'b111111100;
    x_27 = 'b111111010;
    x_28 = 'b000000110;
    x_29 = 'b111101011;
    x_30 = 'b000001100;
    x_31 = 'b000000011;
    x_32 = 'b000000110;
    x_33 = 'b000000100;
    x_34 = 'b111111101;
    x_35 = 'b111110101;
    x_36 = 'b111111011;
    x_37 = 'b111010111;
    x_38 = 'b111110101;
    x_39 = 'b000000001;
    x_40 = 'b000000001;
    x_41 = 'b111110110;
    x_42 = 'b000001100;
    x_43 = 'b111101111;
    x_44 = 'b000010010;
    x_45 = 'b000010101;
    x_46 = 'b000010010;
    x_47 = 'b000010010;
    x_48 = 'b000010101;
    x_49 = 'b000010001;
    x_50 = 'b000010101;
    x_51 = 'b000011010;
    x_52 = 'b000011001;
    x_53 = 'b000010111;
    x_54 = 'b000011001;
    x_55 = 'b000010000;
    x_56 = 'b000010010;
    x_57 = 'b000010010;
    x_58 = 'b000100100;
    x_59 = 'b000011111;
    x_60 = 'b000001111;
    x_61 = 'b000100011;
    x_62 = 'b000011101;
    x_63 = 'b000010000;

    h_0 = 'b000001010;
    h_1 = 'b000011001;
    h_2 = 'b000001110;
    h_3 = 'b000010110;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111111010;
    x_1 = 'b000000110;
    x_2 = 'b000000001;
    x_3 = 'b000001001;
    x_4 = 'b000000000;
    x_5 = 'b111111110;
    x_6 = 'b000000001;
    x_7 = 'b000000101;
    x_8 = 'b111111111;
    x_9 = 'b000001000;
    x_10 = 'b000001001;
    x_11 = 'b000000001;
    x_12 = 'b000000110;
    x_13 = 'b000000011;
    x_14 = 'b000000101;
    x_15 = 'b000001001;
    x_16 = 'b000001000;
    x_17 = 'b000001111;
    x_18 = 'b000000110;
    x_19 = 'b000001001;
    x_20 = 'b000010011;
    x_21 = 'b111111110;
    x_22 = 'b000000100;
    x_23 = 'b000001010;
    x_24 = 'b000000001;
    x_25 = 'b000000001;
    x_26 = 'b111111011;
    x_27 = 'b111111101;
    x_28 = 'b000001100;
    x_29 = 'b111111011;
    x_30 = 'b000001100;
    x_31 = 'b000000010;
    x_32 = 'b000000000;
    x_33 = 'b000000000;
    x_34 = 'b111111001;
    x_35 = 'b111110010;
    x_36 = 'b111111111;
    x_37 = 'b111011111;
    x_38 = 'b000000100;
    x_39 = 'b000000111;
    x_40 = 'b000010101;
    x_41 = 'b111101111;
    x_42 = 'b000010010;
    x_43 = 'b111110101;
    x_44 = 'b000010001;
    x_45 = 'b000100100;
    x_46 = 'b000010000;
    x_47 = 'b000010000;
    x_48 = 'b000010101;
    x_49 = 'b000010000;
    x_50 = 'b000001111;
    x_51 = 'b000010011;
    x_52 = 'b000010010;
    x_53 = 'b000010010;
    x_54 = 'b000011110;
    x_55 = 'b000010001;
    x_56 = 'b000010111;
    x_57 = 'b000010001;
    x_58 = 'b000011101;
    x_59 = 'b000011100;
    x_60 = 'b000001001;
    x_61 = 'b000011010;
    x_62 = 'b000010001;
    x_63 = 'b000001000;

    h_0 = 'b111111010;
    h_1 = 'b000000110;
    h_2 = 'b000000001;
    h_3 = 'b000001001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000001001;
    x_1 = 'b000001001;
    x_2 = 'b111111110;
    x_3 = 'b000000001;
    x_4 = 'b111111000;
    x_5 = 'b111110111;
    x_6 = 'b111111100;
    x_7 = 'b000011000;
    x_8 = 'b000000110;
    x_9 = 'b000001001;
    x_10 = 'b000001001;
    x_11 = 'b111111011;
    x_12 = 'b111111101;
    x_13 = 'b111111001;
    x_14 = 'b000010011;
    x_15 = 'b000010001;
    x_16 = 'b000001100;
    x_17 = 'b000001111;
    x_18 = 'b000000000;
    x_19 = 'b111111111;
    x_20 = 'b000001010;
    x_21 = 'b000000101;
    x_22 = 'b000001010;
    x_23 = 'b000001110;
    x_24 = 'b000001011;
    x_25 = 'b000001011;
    x_26 = 'b111110111;
    x_27 = 'b111111010;
    x_28 = 'b000001000;
    x_29 = 'b000000010;
    x_30 = 'b000010101;
    x_31 = 'b111111010;
    x_32 = 'b111111010;
    x_33 = 'b111111001;
    x_34 = 'b111110010;
    x_35 = 'b111101100;
    x_36 = 'b111110110;
    x_37 = 'b111011100;
    x_38 = 'b000010000;
    x_39 = 'b111110110;
    x_40 = 'b000011010;
    x_41 = 'b111100100;
    x_42 = 'b000001111;
    x_43 = 'b000011000;
    x_44 = 'b000010110;
    x_45 = 'b000010000;
    x_46 = 'b000010110;
    x_47 = 'b000010100;
    x_48 = 'b000010101;
    x_49 = 'b000001111;
    x_50 = 'b000000101;
    x_51 = 'b000000011;
    x_52 = 'b111111110;
    x_53 = 'b111111101;
    x_54 = 'b000001010;
    x_55 = 'b000010110;
    x_56 = 'b000011001;
    x_57 = 'b000001001;
    x_58 = 'b000001001;
    x_59 = 'b000001000;
    x_60 = 'b000001010;
    x_61 = 'b000010110;
    x_62 = 'b000001010;
    x_63 = 'b000001001;

    h_0 = 'b000001001;
    h_1 = 'b000001001;
    h_2 = 'b111111110;
    h_3 = 'b000000001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000001010;
    x_1 = 'b000001010;
    x_2 = 'b111111011;
    x_3 = 'b111111101;
    x_4 = 'b111110000;
    x_5 = 'b111101001;
    x_6 = 'b111110000;
    x_7 = 'b000011011;
    x_8 = 'b000001101;
    x_9 = 'b000001000;
    x_10 = 'b000000011;
    x_11 = 'b111111010;
    x_12 = 'b111110000;
    x_13 = 'b111101010;
    x_14 = 'b000010110;
    x_15 = 'b000010000;
    x_16 = 'b000001011;
    x_17 = 'b000001010;
    x_18 = 'b111110111;
    x_19 = 'b111110010;
    x_20 = 'b111111001;
    x_21 = 'b000000001;
    x_22 = 'b000000111;
    x_23 = 'b000001001;
    x_24 = 'b000001001;
    x_25 = 'b000001001;
    x_26 = 'b111111010;
    x_27 = 'b111111000;
    x_28 = 'b000000011;
    x_29 = 'b000000111;
    x_30 = 'b000010011;
    x_31 = 'b111111111;
    x_32 = 'b111111111;
    x_33 = 'b000000000;
    x_34 = 'b111110111;
    x_35 = 'b111101111;
    x_36 = 'b111111000;
    x_37 = 'b111011100;
    x_38 = 'b000010011;
    x_39 = 'b111110111;
    x_40 = 'b000011101;
    x_41 = 'b000000101;
    x_42 = 'b000101100;
    x_43 = 'b111111010;
    x_44 = 'b000100101;
    x_45 = 'b000000100;
    x_46 = 'b000100010;
    x_47 = 'b000011011;
    x_48 = 'b000011010;
    x_49 = 'b000010011;
    x_50 = 'b000001010;
    x_51 = 'b000000000;
    x_52 = 'b111111100;
    x_53 = 'b111110111;
    x_54 = 'b000000001;
    x_55 = 'b000100001;
    x_56 = 'b000100001;
    x_57 = 'b000001010;
    x_58 = 'b111111110;
    x_59 = 'b000000000;
    x_60 = 'b000010010;
    x_61 = 'b000010110;
    x_62 = 'b000000001;
    x_63 = 'b000001100;

    h_0 = 'b000001010;
    h_1 = 'b000001010;
    h_2 = 'b111111011;
    h_3 = 'b111111101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000011000;
    x_1 = 'b000011100;
    x_2 = 'b000001101;
    x_3 = 'b000001111;
    x_4 = 'b000000111;
    x_5 = 'b111111101;
    x_6 = 'b000000110;
    x_7 = 'b000101101;
    x_8 = 'b000011101;
    x_9 = 'b000011001;
    x_10 = 'b000010101;
    x_11 = 'b000001001;
    x_12 = 'b000000000;
    x_13 = 'b000000111;
    x_14 = 'b000100001;
    x_15 = 'b000011100;
    x_16 = 'b000010110;
    x_17 = 'b000010111;
    x_18 = 'b000000100;
    x_19 = 'b111111010;
    x_20 = 'b000000010;
    x_21 = 'b000010011;
    x_22 = 'b000011001;
    x_23 = 'b000011000;
    x_24 = 'b000011100;
    x_25 = 'b000011100;
    x_26 = 'b000001110;
    x_27 = 'b000001011;
    x_28 = 'b000010100;
    x_29 = 'b000011110;
    x_30 = 'b000100011;
    x_31 = 'b000010001;
    x_32 = 'b000010010;
    x_33 = 'b000010100;
    x_34 = 'b000001100;
    x_35 = 'b000000011;
    x_36 = 'b000001010;
    x_37 = 'b111101011;
    x_38 = 'b000100100;
    x_39 = 'b000010001;
    x_40 = 'b000100101;
    x_41 = 'b000010001;
    x_42 = 'b000111101;
    x_43 = 'b111110101;
    x_44 = 'b000101111;
    x_45 = 'b111111011;
    x_46 = 'b000101100;
    x_47 = 'b000011111;
    x_48 = 'b000011011;
    x_49 = 'b000010010;
    x_50 = 'b000000100;
    x_51 = 'b111101110;
    x_52 = 'b111101010;
    x_53 = 'b111100001;
    x_54 = 'b111101100;
    x_55 = 'b000100100;
    x_56 = 'b000100000;
    x_57 = 'b111111011;
    x_58 = 'b111011011;
    x_59 = 'b111100110;
    x_60 = 'b000011000;
    x_61 = 'b000010010;
    x_62 = 'b111110000;
    x_63 = 'b000001101;

    h_0 = 'b000011000;
    h_1 = 'b000011100;
    h_2 = 'b000001101;
    h_3 = 'b000001111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000011111;
    x_1 = 'b000100000;
    x_2 = 'b000001110;
    x_3 = 'b000010111;
    x_4 = 'b000001011;
    x_5 = 'b000000000;
    x_6 = 'b000000000;
    x_7 = 'b000101001;
    x_8 = 'b000011001;
    x_9 = 'b000010110;
    x_10 = 'b000010010;
    x_11 = 'b111111111;
    x_12 = 'b111110111;
    x_13 = 'b111110010;
    x_14 = 'b000011110;
    x_15 = 'b000010011;
    x_16 = 'b000001100;
    x_17 = 'b000001001;
    x_18 = 'b111110101;
    x_19 = 'b111101000;
    x_20 = 'b111101001;
    x_21 = 'b000010100;
    x_22 = 'b000011010;
    x_23 = 'b000011011;
    x_24 = 'b000010111;
    x_25 = 'b000011000;
    x_26 = 'b000001100;
    x_27 = 'b000001010;
    x_28 = 'b000010011;
    x_29 = 'b000010111;
    x_30 = 'b000011001;
    x_31 = 'b000001010;
    x_32 = 'b000001101;
    x_33 = 'b000001110;
    x_34 = 'b000001000;
    x_35 = 'b111111110;
    x_36 = 'b000000100;
    x_37 = 'b111100010;
    x_38 = 'b000010100;
    x_39 = 'b111111111;
    x_40 = 'b000100010;
    x_41 = 'b111011000;
    x_42 = 'b000101001;
    x_43 = 'b000010100;
    x_44 = 'b000101010;
    x_45 = 'b111101011;
    x_46 = 'b000101000;
    x_47 = 'b000010010;
    x_48 = 'b000001000;
    x_49 = 'b000000001;
    x_50 = 'b111101111;
    x_51 = 'b111010101;
    x_52 = 'b111010000;
    x_53 = 'b111001100;
    x_54 = 'b111011111;
    x_55 = 'b000011011;
    x_56 = 'b000010101;
    x_57 = 'b111101010;
    x_58 = 'b111000011;
    x_59 = 'b111011000;
    x_60 = 'b000010101;
    x_61 = 'b000000101;
    x_62 = 'b111011010;
    x_63 = 'b000001101;

    h_0 = 'b000011111;
    h_1 = 'b000100000;
    h_2 = 'b000001110;
    h_3 = 'b000010111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000001100;
    x_1 = 'b000010101;
    x_2 = 'b111111110;
    x_3 = 'b000010010;
    x_4 = 'b000000110;
    x_5 = 'b111111000;
    x_6 = 'b111111011;
    x_7 = 'b000011101;
    x_8 = 'b000001110;
    x_9 = 'b000001101;
    x_10 = 'b000001001;
    x_11 = 'b111111011;
    x_12 = 'b111111000;
    x_13 = 'b111101101;
    x_14 = 'b000010110;
    x_15 = 'b000001011;
    x_16 = 'b000000010;
    x_17 = 'b111111111;
    x_18 = 'b111110001;
    x_19 = 'b111101100;
    x_20 = 'b111101111;
    x_21 = 'b000001000;
    x_22 = 'b000010000;
    x_23 = 'b000010011;
    x_24 = 'b000001110;
    x_25 = 'b000001110;
    x_26 = 'b000000101;
    x_27 = 'b000000010;
    x_28 = 'b000001101;
    x_29 = 'b000000101;
    x_30 = 'b000001111;
    x_31 = 'b000001000;
    x_32 = 'b000001010;
    x_33 = 'b000001110;
    x_34 = 'b000000101;
    x_35 = 'b111111000;
    x_36 = 'b000000011;
    x_37 = 'b111011100;
    x_38 = 'b111111111;
    x_39 = 'b000000110;
    x_40 = 'b000010011;
    x_41 = 'b111101100;
    x_42 = 'b000011010;
    x_43 = 'b111110000;
    x_44 = 'b000011000;
    x_45 = 'b111111101;
    x_46 = 'b000011000;
    x_47 = 'b000001101;
    x_48 = 'b000001000;
    x_49 = 'b111111010;
    x_50 = 'b111101110;
    x_51 = 'b111011011;
    x_52 = 'b111011001;
    x_53 = 'b111010101;
    x_54 = 'b111100011;
    x_55 = 'b000010110;
    x_56 = 'b000001111;
    x_57 = 'b111100101;
    x_58 = 'b111001001;
    x_59 = 'b111011001;
    x_60 = 'b000001111;
    x_61 = 'b111111000;
    x_62 = 'b111001110;
    x_63 = 'b000001011;

    h_0 = 'b000001100;
    h_1 = 'b000010101;
    h_2 = 'b111111110;
    h_3 = 'b000010010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111110101;
    x_1 = 'b111110101;
    x_2 = 'b111110000;
    x_3 = 'b111110001;
    x_4 = 'b111101100;
    x_5 = 'b111011100;
    x_6 = 'b111011000;
    x_7 = 'b111111101;
    x_8 = 'b111110001;
    x_9 = 'b111101101;
    x_10 = 'b111101100;
    x_11 = 'b111100101;
    x_12 = 'b111011101;
    x_13 = 'b111001000;
    x_14 = 'b111111101;
    x_15 = 'b111110011;
    x_16 = 'b111101110;
    x_17 = 'b111101001;
    x_18 = 'b111101001;
    x_19 = 'b111100101;
    x_20 = 'b111100001;
    x_21 = 'b111110110;
    x_22 = 'b111101010;
    x_23 = 'b111110001;
    x_24 = 'b111110101;
    x_25 = 'b111110110;
    x_26 = 'b111100110;
    x_27 = 'b111101010;
    x_28 = 'b111101010;
    x_29 = 'b111110111;
    x_30 = 'b111101001;
    x_31 = 'b111110110;
    x_32 = 'b111110001;
    x_33 = 'b111101001;
    x_34 = 'b111100011;
    x_35 = 'b111011110;
    x_36 = 'b111011100;
    x_37 = 'b111000011;
    x_38 = 'b111110001;
    x_39 = 'b111000111;
    x_40 = 'b111110000;
    x_41 = 'b111010101;
    x_42 = 'b111111100;
    x_43 = 'b111110110;
    x_44 = 'b111011100;
    x_45 = 'b111011000;
    x_46 = 'b111111110;
    x_47 = 'b111111000;
    x_48 = 'b111110011;
    x_49 = 'b111111010;
    x_50 = 'b111110001;
    x_51 = 'b111110010;
    x_52 = 'b111110010;
    x_53 = 'b111101000;
    x_54 = 'b111100100;
    x_55 = 'b111111000;
    x_56 = 'b111111110;
    x_57 = 'b111111110;
    x_58 = 'b000000010;
    x_59 = 'b000000001;
    x_60 = 'b111110110;
    x_61 = 'b111101110;
    x_62 = 'b111110100;
    x_63 = 'b111100001;

    h_0 = 'b111110101;
    h_1 = 'b111110101;
    h_2 = 'b111110000;
    h_3 = 'b111110001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111100100;
    x_1 = 'b111100100;
    x_2 = 'b111011111;
    x_3 = 'b111011101;
    x_4 = 'b111011011;
    x_5 = 'b111001111;
    x_6 = 'b111001111;
    x_7 = 'b111110101;
    x_8 = 'b111101000;
    x_9 = 'b111100010;
    x_10 = 'b111100010;
    x_11 = 'b111100000;
    x_12 = 'b111011110;
    x_13 = 'b111010001;
    x_14 = 'b111110110;
    x_15 = 'b111101110;
    x_16 = 'b111101001;
    x_17 = 'b111100101;
    x_18 = 'b111101010;
    x_19 = 'b111101101;
    x_20 = 'b111101010;
    x_21 = 'b111101010;
    x_22 = 'b111011111;
    x_23 = 'b111100110;
    x_24 = 'b111101011;
    x_25 = 'b111101011;
    x_26 = 'b111010110;
    x_27 = 'b111011011;
    x_28 = 'b111011110;
    x_29 = 'b111101000;
    x_30 = 'b111011010;
    x_31 = 'b111101000;
    x_32 = 'b111100000;
    x_33 = 'b111011000;
    x_34 = 'b111010011;
    x_35 = 'b111001101;
    x_36 = 'b111001111;
    x_37 = 'b111000100;
    x_38 = 'b111100011;
    x_39 = 'b111001100;
    x_40 = 'b111100100;
    x_41 = 'b111100110;
    x_42 = 'b111100001;
    x_43 = 'b111001010;
    x_44 = 'b111001111;
    x_45 = 'b111101001;
    x_46 = 'b111110010;
    x_47 = 'b111111000;
    x_48 = 'b111111001;
    x_49 = 'b000000100;
    x_50 = 'b111111001;
    x_51 = 'b111111111;
    x_52 = 'b000000000;
    x_53 = 'b111110111;
    x_54 = 'b111110101;
    x_55 = 'b111111110;
    x_56 = 'b000000110;
    x_57 = 'b000001011;
    x_58 = 'b000001111;
    x_59 = 'b000010000;
    x_60 = 'b111111010;
    x_61 = 'b111110111;
    x_62 = 'b000000001;
    x_63 = 'b111101101;

    h_0 = 'b111100100;
    h_1 = 'b111100100;
    h_2 = 'b111011111;
    h_3 = 'b111011101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111100010;
    x_1 = 'b111100001;
    x_2 = 'b111011011;
    x_3 = 'b111011101;
    x_4 = 'b111011011;
    x_5 = 'b111010011;
    x_6 = 'b111001110;
    x_7 = 'b111110001;
    x_8 = 'b111101000;
    x_9 = 'b111100111;
    x_10 = 'b111101101;
    x_11 = 'b111101111;
    x_12 = 'b111101010;
    x_13 = 'b111100010;
    x_14 = 'b111101110;
    x_15 = 'b111110001;
    x_16 = 'b111110001;
    x_17 = 'b111101111;
    x_18 = 'b111110101;
    x_19 = 'b111111010;
    x_20 = 'b111111000;
    x_21 = 'b111100111;
    x_22 = 'b111011011;
    x_23 = 'b111100011;
    x_24 = 'b111101000;
    x_25 = 'b111101001;
    x_26 = 'b111011000;
    x_27 = 'b111011011;
    x_28 = 'b111011001;
    x_29 = 'b111100111;
    x_30 = 'b111011010;
    x_31 = 'b111101111;
    x_32 = 'b111101000;
    x_33 = 'b111100010;
    x_34 = 'b111011100;
    x_35 = 'b111010110;
    x_36 = 'b111011000;
    x_37 = 'b111000110;
    x_38 = 'b111101010;
    x_39 = 'b111011011;
    x_40 = 'b111110011;
    x_41 = 'b111111110;
    x_42 = 'b111110101;
    x_43 = 'b110111011;
    x_44 = 'b111011011;
    x_45 = 'b111110001;
    x_46 = 'b000000000;
    x_47 = 'b000000101;
    x_48 = 'b000000111;
    x_49 = 'b000010101;
    x_50 = 'b000001001;
    x_51 = 'b000001011;
    x_52 = 'b000001010;
    x_53 = 'b000000011;
    x_54 = 'b000000100;
    x_55 = 'b000001111;
    x_56 = 'b000011000;
    x_57 = 'b000011011;
    x_58 = 'b000010111;
    x_59 = 'b000011100;
    x_60 = 'b000001010;
    x_61 = 'b000001000;
    x_62 = 'b000010001;
    x_63 = 'b000000011;

    h_0 = 'b111100010;
    h_1 = 'b111100001;
    h_2 = 'b111011011;
    h_3 = 'b111011101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111101101;
    x_1 = 'b111110101;
    x_2 = 'b111110011;
    x_3 = 'b111110100;
    x_4 = 'b111110011;
    x_5 = 'b111101100;
    x_6 = 'b111100111;
    x_7 = 'b000000101;
    x_8 = 'b111111110;
    x_9 = 'b111111110;
    x_10 = 'b000000100;
    x_11 = 'b000000110;
    x_12 = 'b111111111;
    x_13 = 'b111110011;
    x_14 = 'b000001000;
    x_15 = 'b000001000;
    x_16 = 'b000001000;
    x_17 = 'b000000101;
    x_18 = 'b000001010;
    x_19 = 'b000001100;
    x_20 = 'b000001001;
    x_21 = 'b111110011;
    x_22 = 'b111100111;
    x_23 = 'b111101100;
    x_24 = 'b111110011;
    x_25 = 'b111110100;
    x_26 = 'b111101100;
    x_27 = 'b111101101;
    x_28 = 'b111100110;
    x_29 = 'b111110010;
    x_30 = 'b111101000;
    x_31 = 'b000000010;
    x_32 = 'b111111111;
    x_33 = 'b111111000;
    x_34 = 'b111110000;
    x_35 = 'b111101110;
    x_36 = 'b111101111;
    x_37 = 'b111010011;
    x_38 = 'b111111111;
    x_39 = 'b111101000;
    x_40 = 'b000000110;
    x_41 = 'b111111100;
    x_42 = 'b000001010;
    x_43 = 'b111110110;
    x_44 = 'b111110010;
    x_45 = 'b111111101;
    x_46 = 'b000011000;
    x_47 = 'b000011101;
    x_48 = 'b000011100;
    x_49 = 'b000101001;
    x_50 = 'b000011111;
    x_51 = 'b000011011;
    x_52 = 'b000010111;
    x_53 = 'b000001110;
    x_54 = 'b000010011;
    x_55 = 'b000100100;
    x_56 = 'b000101100;
    x_57 = 'b000101111;
    x_58 = 'b000100010;
    x_59 = 'b000100011;
    x_60 = 'b000100011;
    x_61 = 'b000100001;
    x_62 = 'b000100001;
    x_63 = 'b000011110;

    h_0 = 'b111101101;
    h_1 = 'b111110101;
    h_2 = 'b111110011;
    h_3 = 'b111110100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111111100;
    x_1 = 'b000000110;
    x_2 = 'b111111111;
    x_3 = 'b111111100;
    x_4 = 'b111111000;
    x_5 = 'b111110001;
    x_6 = 'b111101111;
    x_7 = 'b000011000;
    x_8 = 'b000001011;
    x_9 = 'b000001000;
    x_10 = 'b000001010;
    x_11 = 'b000000010;
    x_12 = 'b111111101;
    x_13 = 'b111100111;
    x_14 = 'b000010111;
    x_15 = 'b000010011;
    x_16 = 'b000010000;
    x_17 = 'b000001011;
    x_18 = 'b000001101;
    x_19 = 'b000001010;
    x_20 = 'b000000001;
    x_21 = 'b111110011;
    x_22 = 'b111101011;
    x_23 = 'b111101110;
    x_24 = 'b111110100;
    x_25 = 'b111110110;
    x_26 = 'b111101101;
    x_27 = 'b111110000;
    x_28 = 'b111101010;
    x_29 = 'b111111111;
    x_30 = 'b111100001;
    x_31 = 'b000000100;
    x_32 = 'b111111110;
    x_33 = 'b111110100;
    x_34 = 'b111101101;
    x_35 = 'b111101011;
    x_36 = 'b111110000;
    x_37 = 'b111010100;
    x_38 = 'b000000100;
    x_39 = 'b111100011;
    x_40 = 'b000001110;
    x_41 = 'b111101010;
    x_42 = 'b000000111;
    x_43 = 'b111100011;
    x_44 = 'b111110111;
    x_45 = 'b111110101;
    x_46 = 'b000011111;
    x_47 = 'b000100010;
    x_48 = 'b000100010;
    x_49 = 'b000101010;
    x_50 = 'b000100000;
    x_51 = 'b000011010;
    x_52 = 'b000010100;
    x_53 = 'b000000111;
    x_54 = 'b000000100;
    x_55 = 'b000101100;
    x_56 = 'b000110010;
    x_57 = 'b000110110;
    x_58 = 'b000100000;
    x_59 = 'b000011011;
    x_60 = 'b000110111;
    x_61 = 'b000110001;
    x_62 = 'b000100111;
    x_63 = 'b000101100;

    h_0 = 'b111111100;
    h_1 = 'b000000110;
    h_2 = 'b111111111;
    h_3 = 'b111111100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000000010;
    x_1 = 'b000000010;
    x_2 = 'b111111001;
    x_3 = 'b111110010;
    x_4 = 'b111101110;
    x_5 = 'b111101000;
    x_6 = 'b111101001;
    x_7 = 'b000011001;
    x_8 = 'b000001010;
    x_9 = 'b000000011;
    x_10 = 'b111111111;
    x_11 = 'b111110011;
    x_12 = 'b111110011;
    x_13 = 'b111100011;
    x_14 = 'b000011100;
    x_15 = 'b000010101;
    x_16 = 'b000001110;
    x_17 = 'b000001000;
    x_18 = 'b000001000;
    x_19 = 'b000000100;
    x_20 = 'b111111111;
    x_21 = 'b111110101;
    x_22 = 'b111101101;
    x_23 = 'b111110001;
    x_24 = 'b111111000;
    x_25 = 'b111111010;
    x_26 = 'b111101101;
    x_27 = 'b111110010;
    x_28 = 'b111101110;
    x_29 = 'b000000111;
    x_30 = 'b111101101;
    x_31 = 'b000000100;
    x_32 = 'b000000000;
    x_33 = 'b111110111;
    x_34 = 'b111101111;
    x_35 = 'b111101110;
    x_36 = 'b111110001;
    x_37 = 'b111010110;
    x_38 = 'b000011000;
    x_39 = 'b111101100;
    x_40 = 'b000011101;
    x_41 = 'b000000110;
    x_42 = 'b000011000;
    x_43 = 'b111010100;
    x_44 = 'b000000001;
    x_45 = 'b111110100;
    x_46 = 'b000101110;
    x_47 = 'b000101110;
    x_48 = 'b000101100;
    x_49 = 'b000110011;
    x_50 = 'b000100101;
    x_51 = 'b000011110;
    x_52 = 'b000011001;
    x_53 = 'b000001011;
    x_54 = 'b000000100;
    x_55 = 'b000111001;
    x_56 = 'b000111100;
    x_57 = 'b000111110;
    x_58 = 'b000100011;
    x_59 = 'b000011110;
    x_60 = 'b001000011;
    x_61 = 'b000111001;
    x_62 = 'b000100110;
    x_63 = 'b000101110;

    h_0 = 'b000000010;
    h_1 = 'b000000010;
    h_2 = 'b111111001;
    h_3 = 'b111110010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000010011;
    x_1 = 'b000010010;
    x_2 = 'b000000110;
    x_3 = 'b111111101;
    x_4 = 'b111111000;
    x_5 = 'b111101111;
    x_6 = 'b111101110;
    x_7 = 'b000101101;
    x_8 = 'b000011101;
    x_9 = 'b000010011;
    x_10 = 'b000001011;
    x_11 = 'b111111101;
    x_12 = 'b111111011;
    x_13 = 'b111101110;
    x_14 = 'b000110000;
    x_15 = 'b000101000;
    x_16 = 'b000011101;
    x_17 = 'b000010100;
    x_18 = 'b000010010;
    x_19 = 'b000001110;
    x_20 = 'b000001001;
    x_21 = 'b111111100;
    x_22 = 'b111110001;
    x_23 = 'b111110100;
    x_24 = 'b111111110;
    x_25 = 'b111111111;
    x_26 = 'b111110011;
    x_27 = 'b111110101;
    x_28 = 'b111101101;
    x_29 = 'b000001101;
    x_30 = 'b111111001;
    x_31 = 'b000001001;
    x_32 = 'b000001000;
    x_33 = 'b111111110;
    x_34 = 'b111110110;
    x_35 = 'b111110011;
    x_36 = 'b111101101;
    x_37 = 'b111010001;
    x_38 = 'b000011100;
    x_39 = 'b111100101;
    x_40 = 'b000011100;
    x_41 = 'b111110011;
    x_42 = 'b000001110;
    x_43 = 'b111011011;
    x_44 = 'b000001111;
    x_45 = 'b111111000;
    x_46 = 'b000110110;
    x_47 = 'b000110111;
    x_48 = 'b000110101;
    x_49 = 'b000111100;
    x_50 = 'b000101101;
    x_51 = 'b000100101;
    x_52 = 'b000100000;
    x_53 = 'b000010011;
    x_54 = 'b000001101;
    x_55 = 'b000111101;
    x_56 = 'b001000000;
    x_57 = 'b001000001;
    x_58 = 'b000101000;
    x_59 = 'b000100101;
    x_60 = 'b001001000;
    x_61 = 'b000111110;
    x_62 = 'b000101001;
    x_63 = 'b000110011;

    h_0 = 'b000010011;
    h_1 = 'b000010010;
    h_2 = 'b000000110;
    h_3 = 'b111111101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000001111;
    x_1 = 'b000010011;
    x_2 = 'b000000110;
    x_3 = 'b000000001;
    x_4 = 'b111111011;
    x_5 = 'b111110000;
    x_6 = 'b111110000;
    x_7 = 'b000101001;
    x_8 = 'b000100000;
    x_9 = 'b000010110;
    x_10 = 'b000010100;
    x_11 = 'b000000110;
    x_12 = 'b000000011;
    x_13 = 'b111110011;
    x_14 = 'b000101011;
    x_15 = 'b000101010;
    x_16 = 'b000100011;
    x_17 = 'b000011001;
    x_18 = 'b000010111;
    x_19 = 'b000010010;
    x_20 = 'b000001100;
    x_21 = 'b111110111;
    x_22 = 'b111101011;
    x_23 = 'b111101110;
    x_24 = 'b111110111;
    x_25 = 'b111111001;
    x_26 = 'b111101010;
    x_27 = 'b111101101;
    x_28 = 'b111100110;
    x_29 = 'b000000011;
    x_30 = 'b111110011;
    x_31 = 'b000000010;
    x_32 = 'b111111101;
    x_33 = 'b111110011;
    x_34 = 'b111101101;
    x_35 = 'b111100111;
    x_36 = 'b111100110;
    x_37 = 'b111001110;
    x_38 = 'b000001111;
    x_39 = 'b111100000;
    x_40 = 'b000001100;
    x_41 = 'b111110101;
    x_42 = 'b000010100;
    x_43 = 'b111000110;
    x_44 = 'b000001110;
    x_45 = 'b111110001;
    x_46 = 'b000101000;
    x_47 = 'b000101110;
    x_48 = 'b000101111;
    x_49 = 'b000111000;
    x_50 = 'b000101001;
    x_51 = 'b000011111;
    x_52 = 'b000011010;
    x_53 = 'b000001100;
    x_54 = 'b000001100;
    x_55 = 'b000110111;
    x_56 = 'b000111011;
    x_57 = 'b000111011;
    x_58 = 'b000100010;
    x_59 = 'b000011111;
    x_60 = 'b001001000;
    x_61 = 'b000111111;
    x_62 = 'b000101111;
    x_63 = 'b000111010;

    h_0 = 'b000001111;
    h_1 = 'b000010011;
    h_2 = 'b000000110;
    h_3 = 'b000000001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000000011;
    x_1 = 'b000001001;
    x_2 = 'b000000010;
    x_3 = 'b111111101;
    x_4 = 'b111111001;
    x_5 = 'b111101101;
    x_6 = 'b111101011;
    x_7 = 'b000011011;
    x_8 = 'b000011001;
    x_9 = 'b000010100;
    x_10 = 'b000010101;
    x_11 = 'b000001001;
    x_12 = 'b111111110;
    x_13 = 'b111100100;
    x_14 = 'b000100101;
    x_15 = 'b000100110;
    x_16 = 'b000100000;
    x_17 = 'b000010101;
    x_18 = 'b000010011;
    x_19 = 'b000001010;
    x_20 = 'b111111100;
    x_21 = 'b111111000;
    x_22 = 'b111101101;
    x_23 = 'b111101111;
    x_24 = 'b111111001;
    x_25 = 'b111111011;
    x_26 = 'b111101101;
    x_27 = 'b111110000;
    x_28 = 'b111101011;
    x_29 = 'b000000110;
    x_30 = 'b111110111;
    x_31 = 'b000000111;
    x_32 = 'b000000101;
    x_33 = 'b111111100;
    x_34 = 'b111110100;
    x_35 = 'b111110001;
    x_36 = 'b111101101;
    x_37 = 'b111011011;
    x_38 = 'b000010000;
    x_39 = 'b111100111;
    x_40 = 'b000010100;
    x_41 = 'b111101001;
    x_42 = 'b000011011;
    x_43 = 'b111101000;
    x_44 = 'b000001101;
    x_45 = 'b111101110;
    x_46 = 'b000100110;
    x_47 = 'b000101101;
    x_48 = 'b000101110;
    x_49 = 'b000110100;
    x_50 = 'b000101000;
    x_51 = 'b000011010;
    x_52 = 'b000010011;
    x_53 = 'b000000011;
    x_54 = 'b000000100;
    x_55 = 'b000111001;
    x_56 = 'b000111100;
    x_57 = 'b000111000;
    x_58 = 'b000011011;
    x_59 = 'b000011001;
    x_60 = 'b001000011;
    x_61 = 'b000111001;
    x_62 = 'b000101110;
    x_63 = 'b000110011;

    h_0 = 'b000000011;
    h_1 = 'b000001001;
    h_2 = 'b000000010;
    h_3 = 'b111111101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000010001;
    x_1 = 'b000011101;
    x_2 = 'b000010111;
    x_3 = 'b000010011;
    x_4 = 'b000001011;
    x_5 = 'b111111011;
    x_6 = 'b111101111;
    x_7 = 'b000110010;
    x_8 = 'b000101100;
    x_9 = 'b000100111;
    x_10 = 'b000100010;
    x_11 = 'b000010111;
    x_12 = 'b000000110;
    x_13 = 'b111100011;
    x_14 = 'b000111100;
    x_15 = 'b000110100;
    x_16 = 'b000101101;
    x_17 = 'b000100001;
    x_18 = 'b000011101;
    x_19 = 'b000010010;
    x_20 = 'b000000001;
    x_21 = 'b111111001;
    x_22 = 'b111110000;
    x_23 = 'b111110100;
    x_24 = 'b111111110;
    x_25 = 'b000000000;
    x_26 = 'b111111010;
    x_27 = 'b111111010;
    x_28 = 'b111110010;
    x_29 = 'b000001110;
    x_30 = 'b000000000;
    x_31 = 'b000010110;
    x_32 = 'b000010011;
    x_33 = 'b000001011;
    x_34 = 'b000000011;
    x_35 = 'b111111101;
    x_36 = 'b111110110;
    x_37 = 'b111100000;
    x_38 = 'b000010101;
    x_39 = 'b111101011;
    x_40 = 'b000010011;
    x_41 = 'b111100111;
    x_42 = 'b000011111;
    x_43 = 'b111110010;
    x_44 = 'b000011100;
    x_45 = 'b000000001;
    x_46 = 'b000110111;
    x_47 = 'b000111100;
    x_48 = 'b000110111;
    x_49 = 'b001000000;
    x_50 = 'b000110011;
    x_51 = 'b000100111;
    x_52 = 'b000100010;
    x_53 = 'b000010001;
    x_54 = 'b000010001;
    x_55 = 'b001000011;
    x_56 = 'b001000110;
    x_57 = 'b001000001;
    x_58 = 'b000100011;
    x_59 = 'b000100000;
    x_60 = 'b001000011;
    x_61 = 'b000111000;
    x_62 = 'b000110000;
    x_63 = 'b000110100;

    h_0 = 'b000010001;
    h_1 = 'b000011101;
    h_2 = 'b000010111;
    h_3 = 'b000010011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000010110;
    x_1 = 'b000011011;
    x_2 = 'b000010101;
    x_3 = 'b000010101;
    x_4 = 'b000001110;
    x_5 = 'b000000001;
    x_6 = 'b111111100;
    x_7 = 'b000100111;
    x_8 = 'b000100011;
    x_9 = 'b000100000;
    x_10 = 'b000011111;
    x_11 = 'b000011001;
    x_12 = 'b000001101;
    x_13 = 'b111111000;
    x_14 = 'b000101100;
    x_15 = 'b000101001;
    x_16 = 'b000100111;
    x_17 = 'b000011101;
    x_18 = 'b000100001;
    x_19 = 'b000011100;
    x_20 = 'b000010010;
    x_21 = 'b111110110;
    x_22 = 'b111101100;
    x_23 = 'b111110010;
    x_24 = 'b111111001;
    x_25 = 'b111111011;
    x_26 = 'b111110011;
    x_27 = 'b111110111;
    x_28 = 'b111110001;
    x_29 = 'b000001110;
    x_30 = 'b111111101;
    x_31 = 'b000001111;
    x_32 = 'b000000111;
    x_33 = 'b000000010;
    x_34 = 'b111111100;
    x_35 = 'b111110110;
    x_36 = 'b111110011;
    x_37 = 'b111100001;
    x_38 = 'b000011100;
    x_39 = 'b111111000;
    x_40 = 'b000101001;
    x_41 = 'b000011011;
    x_42 = 'b000101101;
    x_43 = 'b111110101;
    x_44 = 'b000011110;
    x_45 = 'b000001101;
    x_46 = 'b000101100;
    x_47 = 'b000101101;
    x_48 = 'b000100110;
    x_49 = 'b000110101;
    x_50 = 'b000101000;
    x_51 = 'b000100010;
    x_52 = 'b000100001;
    x_53 = 'b000010101;
    x_54 = 'b000010110;
    x_55 = 'b000110100;
    x_56 = 'b000111001;
    x_57 = 'b000110111;
    x_58 = 'b000100001;
    x_59 = 'b000100000;
    x_60 = 'b001000010;
    x_61 = 'b000111001;
    x_62 = 'b000110001;
    x_63 = 'b000110101;

    h_0 = 'b000010110;
    h_1 = 'b000011011;
    h_2 = 'b000010101;
    h_3 = 'b000010101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000010100;
    x_1 = 'b000010101;
    x_2 = 'b000001110;
    x_3 = 'b000001111;
    x_4 = 'b000001001;
    x_5 = 'b000000000;
    x_6 = 'b000001000;
    x_7 = 'b000011110;
    x_8 = 'b000011010;
    x_9 = 'b000010111;
    x_10 = 'b000011001;
    x_11 = 'b000011010;
    x_12 = 'b000010010;
    x_13 = 'b000001101;
    x_14 = 'b000011111;
    x_15 = 'b000011111;
    x_16 = 'b000011110;
    x_17 = 'b000011001;
    x_18 = 'b000100001;
    x_19 = 'b000100000;
    x_20 = 'b000100010;
    x_21 = 'b111111010;
    x_22 = 'b111110000;
    x_23 = 'b111110100;
    x_24 = 'b111111111;
    x_25 = 'b000000000;
    x_26 = 'b111111001;
    x_27 = 'b111111010;
    x_28 = 'b111110010;
    x_29 = 'b000010100;
    x_30 = 'b000000011;
    x_31 = 'b000010100;
    x_32 = 'b000001111;
    x_33 = 'b000001001;
    x_34 = 'b000000011;
    x_35 = 'b111111111;
    x_36 = 'b111111100;
    x_37 = 'b111101001;
    x_38 = 'b000011110;
    x_39 = 'b000001010;
    x_40 = 'b000100100;
    x_41 = 'b000101011;
    x_42 = 'b000101101;
    x_43 = 'b000000110;
    x_44 = 'b000010010;
    x_45 = 'b000011011;
    x_46 = 'b000100111;
    x_47 = 'b000101010;
    x_48 = 'b000100101;
    x_49 = 'b000110011;
    x_50 = 'b000101001;
    x_51 = 'b000100110;
    x_52 = 'b000101001;
    x_53 = 'b000100001;
    x_54 = 'b000100011;
    x_55 = 'b000101111;
    x_56 = 'b000110011;
    x_57 = 'b000110100;
    x_58 = 'b000100101;
    x_59 = 'b000100110;
    x_60 = 'b000111011;
    x_61 = 'b000110101;
    x_62 = 'b000110011;
    x_63 = 'b000110000;

    h_0 = 'b000010100;
    h_1 = 'b000010101;
    h_2 = 'b000001110;
    h_3 = 'b000001111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000011100;
    x_1 = 'b000100000;
    x_2 = 'b000011100;
    x_3 = 'b000011010;
    x_4 = 'b000010011;
    x_5 = 'b000001100;
    x_6 = 'b000010010;
    x_7 = 'b000101001;
    x_8 = 'b000100110;
    x_9 = 'b000100001;
    x_10 = 'b000100001;
    x_11 = 'b000011111;
    x_12 = 'b000011100;
    x_13 = 'b000010000;
    x_14 = 'b000101000;
    x_15 = 'b000100100;
    x_16 = 'b000100001;
    x_17 = 'b000011101;
    x_18 = 'b000100010;
    x_19 = 'b000100010;
    x_20 = 'b000100100;
    x_21 = 'b111111011;
    x_22 = 'b111101111;
    x_23 = 'b111110001;
    x_24 = 'b111111110;
    x_25 = 'b000000001;
    x_26 = 'b111111100;
    x_27 = 'b111111101;
    x_28 = 'b111110001;
    x_29 = 'b000001111;
    x_30 = 'b000000110;
    x_31 = 'b000011011;
    x_32 = 'b000010010;
    x_33 = 'b000001011;
    x_34 = 'b000000110;
    x_35 = 'b000000010;
    x_36 = 'b000000010;
    x_37 = 'b111110011;
    x_38 = 'b000100010;
    x_39 = 'b000000111;
    x_40 = 'b000101010;
    x_41 = 'b000010101;
    x_42 = 'b000011100;
    x_43 = 'b000010110;
    x_44 = 'b000010001;
    x_45 = 'b000011100;
    x_46 = 'b000100011;
    x_47 = 'b000100011;
    x_48 = 'b000011110;
    x_49 = 'b000101001;
    x_50 = 'b000100000;
    x_51 = 'b000011100;
    x_52 = 'b000011110;
    x_53 = 'b000010111;
    x_54 = 'b000011001;
    x_55 = 'b000100001;
    x_56 = 'b000100101;
    x_57 = 'b000100011;
    x_58 = 'b000011000;
    x_59 = 'b000010101;
    x_60 = 'b000101010;
    x_61 = 'b000011111;
    x_62 = 'b000100100;
    x_63 = 'b000010111;

    h_0 = 'b000011100;
    h_1 = 'b000100000;
    h_2 = 'b000011100;
    h_3 = 'b000011010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000011010;
    x_1 = 'b000100001;
    x_2 = 'b000011010;
    x_3 = 'b000010111;
    x_4 = 'b000010000;
    x_5 = 'b000001010;
    x_6 = 'b000001110;
    x_7 = 'b000101101;
    x_8 = 'b000100111;
    x_9 = 'b000100011;
    x_10 = 'b000100011;
    x_11 = 'b000011011;
    x_12 = 'b000011010;
    x_13 = 'b000001100;
    x_14 = 'b000110000;
    x_15 = 'b000101000;
    x_16 = 'b000100011;
    x_17 = 'b000011110;
    x_18 = 'b000100010;
    x_19 = 'b000100001;
    x_20 = 'b000100001;
    x_21 = 'b111111011;
    x_22 = 'b111110001;
    x_23 = 'b111110000;
    x_24 = 'b111111110;
    x_25 = 'b000000001;
    x_26 = 'b111111101;
    x_27 = 'b111111111;
    x_28 = 'b111110011;
    x_29 = 'b000001110;
    x_30 = 'b000001011;
    x_31 = 'b000011011;
    x_32 = 'b000010110;
    x_33 = 'b000001101;
    x_34 = 'b000000110;
    x_35 = 'b000000011;
    x_36 = 'b000000000;
    x_37 = 'b111110101;
    x_38 = 'b000101001;
    x_39 = 'b000000101;
    x_40 = 'b000100101;
    x_41 = 'b000001100;
    x_42 = 'b000011111;
    x_43 = 'b000100011;
    x_44 = 'b000010110;
    x_45 = 'b000101011;
    x_46 = 'b000101010;
    x_47 = 'b000101010;
    x_48 = 'b000100100;
    x_49 = 'b000110000;
    x_50 = 'b000101001;
    x_51 = 'b000101000;
    x_52 = 'b000101001;
    x_53 = 'b000100011;
    x_54 = 'b000101000;
    x_55 = 'b000100011;
    x_56 = 'b000101000;
    x_57 = 'b000101010;
    x_58 = 'b000100011;
    x_59 = 'b000100000;
    x_60 = 'b000100000;
    x_61 = 'b000010011;
    x_62 = 'b000011100;
    x_63 = 'b000001101;

    h_0 = 'b000011010;
    h_1 = 'b000100001;
    h_2 = 'b000011010;
    h_3 = 'b000010111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000100110;
    x_1 = 'b000101100;
    x_2 = 'b000100011;
    x_3 = 'b000100100;
    x_4 = 'b000011010;
    x_5 = 'b000001110;
    x_6 = 'b000001101;
    x_7 = 'b000110100;
    x_8 = 'b000101101;
    x_9 = 'b000110001;
    x_10 = 'b000110000;
    x_11 = 'b000101011;
    x_12 = 'b000100010;
    x_13 = 'b000010001;
    x_14 = 'b000101011;
    x_15 = 'b000101101;
    x_16 = 'b000101101;
    x_17 = 'b000101010;
    x_18 = 'b000110000;
    x_19 = 'b000101101;
    x_20 = 'b000100111;
    x_21 = 'b111111011;
    x_22 = 'b111110011;
    x_23 = 'b111110011;
    x_24 = 'b111111110;
    x_25 = 'b000000001;
    x_26 = 'b000000010;
    x_27 = 'b000000000;
    x_28 = 'b111110101;
    x_29 = 'b000010111;
    x_30 = 'b000000011;
    x_31 = 'b000011010;
    x_32 = 'b000011000;
    x_33 = 'b000010000;
    x_34 = 'b000001000;
    x_35 = 'b000000010;
    x_36 = 'b111111101;
    x_37 = 'b111101110;
    x_38 = 'b000011011;
    x_39 = 'b000000011;
    x_40 = 'b000001001;
    x_41 = 'b000010100;
    x_42 = 'b000101110;
    x_43 = 'b000100000;
    x_44 = 'b000010010;
    x_45 = 'b000100110;
    x_46 = 'b000100001;
    x_47 = 'b000100010;
    x_48 = 'b000011111;
    x_49 = 'b000101001;
    x_50 = 'b000101000;
    x_51 = 'b000101001;
    x_52 = 'b000101001;
    x_53 = 'b000100001;
    x_54 = 'b000100010;
    x_55 = 'b000011011;
    x_56 = 'b000100100;
    x_57 = 'b000101000;
    x_58 = 'b000100101;
    x_59 = 'b000100001;
    x_60 = 'b000011100;
    x_61 = 'b000010011;
    x_62 = 'b000011110;
    x_63 = 'b000010011;

    h_0 = 'b000100110;
    h_1 = 'b000101100;
    h_2 = 'b000100011;
    h_3 = 'b000100100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000010101;
    x_1 = 'b000011100;
    x_2 = 'b000011001;
    x_3 = 'b000100000;
    x_4 = 'b000011001;
    x_5 = 'b000001100;
    x_6 = 'b000001111;
    x_7 = 'b000010111;
    x_8 = 'b000100000;
    x_9 = 'b000100100;
    x_10 = 'b000100110;
    x_11 = 'b000100010;
    x_12 = 'b000100001;
    x_13 = 'b000010000;
    x_14 = 'b000011101;
    x_15 = 'b000100010;
    x_16 = 'b000100100;
    x_17 = 'b000100001;
    x_18 = 'b000101011;
    x_19 = 'b000101000;
    x_20 = 'b000100011;
    x_21 = 'b111111010;
    x_22 = 'b111110010;
    x_23 = 'b111110011;
    x_24 = 'b111111100;
    x_25 = 'b111111110;
    x_26 = 'b111111111;
    x_27 = 'b000000000;
    x_28 = 'b111110100;
    x_29 = 'b000010011;
    x_30 = 'b111111111;
    x_31 = 'b000011001;
    x_32 = 'b000010000;
    x_33 = 'b000001011;
    x_34 = 'b000000110;
    x_35 = 'b111111111;
    x_36 = 'b111111111;
    x_37 = 'b111110100;
    x_38 = 'b000010111;
    x_39 = 'b000001000;
    x_40 = 'b000011100;
    x_41 = 'b000100000;
    x_42 = 'b000110001;
    x_43 = 'b111110101;
    x_44 = 'b000011010;
    x_45 = 'b000100111;
    x_46 = 'b000011011;
    x_47 = 'b000100010;
    x_48 = 'b000011111;
    x_49 = 'b000101010;
    x_50 = 'b000101001;
    x_51 = 'b000101111;
    x_52 = 'b000101101;
    x_53 = 'b000100111;
    x_54 = 'b000101000;
    x_55 = 'b000011101;
    x_56 = 'b000100111;
    x_57 = 'b000110000;
    x_58 = 'b000110000;
    x_59 = 'b000101101;
    x_60 = 'b000011110;
    x_61 = 'b000011101;
    x_62 = 'b000101011;
    x_63 = 'b000100011;

    h_0 = 'b000010101;
    h_1 = 'b000011100;
    h_2 = 'b000011001;
    h_3 = 'b000100000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111100111;
    x_1 = 'b111011000;
    x_2 = 'b111000111;
    x_3 = 'b110111000;
    x_4 = 'b110111100;
    x_5 = 'b110111000;
    x_6 = 'b111000110;
    x_7 = 'b111101111;
    x_8 = 'b111000110;
    x_9 = 'b111000010;
    x_10 = 'b110111101;
    x_11 = 'b110110101;
    x_12 = 'b111000000;
    x_13 = 'b110110111;
    x_14 = 'b111010010;
    x_15 = 'b111001100;
    x_16 = 'b111000100;
    x_17 = 'b111000000;
    x_18 = 'b111001011;
    x_19 = 'b111001111;
    x_20 = 'b111001011;
    x_21 = 'b111101011;
    x_22 = 'b111011010;
    x_23 = 'b111011001;
    x_24 = 'b111111001;
    x_25 = 'b111110111;
    x_26 = 'b111000010;
    x_27 = 'b110111111;
    x_28 = 'b111010100;
    x_29 = 'b111101110;
    x_30 = 'b111100101;
    x_31 = 'b110111101;
    x_32 = 'b111000001;
    x_33 = 'b110111001;
    x_34 = 'b110110110;
    x_35 = 'b111000000;
    x_36 = 'b110111010;
    x_37 = 'b111101000;
    x_38 = 'b111011110;
    x_39 = 'b110110101;
    x_40 = 'b111001101;
    x_41 = 'b110110110;
    x_42 = 'b111010110;
    x_43 = 'b111100011;
    x_44 = 'b111011010;
    x_45 = 'b111100001;
    x_46 = 'b111011001;
    x_47 = 'b111010101;
    x_48 = 'b111010010;
    x_49 = 'b111001111;
    x_50 = 'b111001001;
    x_51 = 'b111011010;
    x_52 = 'b111100000;
    x_53 = 'b111101010;
    x_54 = 'b111100000;
    x_55 = 'b111110100;
    x_56 = 'b111100010;
    x_57 = 'b111100101;
    x_58 = 'b111110010;
    x_59 = 'b111110100;
    x_60 = 'b000000111;
    x_61 = 'b111110110;
    x_62 = 'b000000100;
    x_63 = 'b000001001;

    h_0 = 'b111100111;
    h_1 = 'b111011000;
    h_2 = 'b111000111;
    h_3 = 'b110111000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111010111;
    x_1 = 'b111001010;
    x_2 = 'b110110101;
    x_3 = 'b110100100;
    x_4 = 'b110100100;
    x_5 = 'b110011100;
    x_6 = 'b110110011;
    x_7 = 'b111100000;
    x_8 = 'b110111001;
    x_9 = 'b110110100;
    x_10 = 'b110101110;
    x_11 = 'b110101001;
    x_12 = 'b110101001;
    x_13 = 'b110101011;
    x_14 = 'b111001001;
    x_15 = 'b111000001;
    x_16 = 'b110111010;
    x_17 = 'b110110110;
    x_18 = 'b110111110;
    x_19 = 'b110111111;
    x_20 = 'b110111110;
    x_21 = 'b111100110;
    x_22 = 'b111010111;
    x_23 = 'b111010111;
    x_24 = 'b111110111;
    x_25 = 'b111110110;
    x_26 = 'b110111001;
    x_27 = 'b110110111;
    x_28 = 'b111010010;
    x_29 = 'b111101110;
    x_30 = 'b111100100;
    x_31 = 'b110110011;
    x_32 = 'b110111000;
    x_33 = 'b110101110;
    x_34 = 'b110101011;
    x_35 = 'b110110101;
    x_36 = 'b110110000;
    x_37 = 'b111100101;
    x_38 = 'b111100000;
    x_39 = 'b110110001;
    x_40 = 'b111010001;
    x_41 = 'b110101000;
    x_42 = 'b111101110;
    x_43 = 'b111000011;
    x_44 = 'b111100100;
    x_45 = 'b111011101;
    x_46 = 'b111100010;
    x_47 = 'b111011001;
    x_48 = 'b111010101;
    x_49 = 'b111010101;
    x_50 = 'b111001111;
    x_51 = 'b111011111;
    x_52 = 'b111100010;
    x_53 = 'b111101010;
    x_54 = 'b111100011;
    x_55 = 'b111110111;
    x_56 = 'b111100110;
    x_57 = 'b111110000;
    x_58 = 'b111110011;
    x_59 = 'b111110010;
    x_60 = 'b111111100;
    x_61 = 'b111101111;
    x_62 = 'b111111001;
    x_63 = 'b111110011;

    h_0 = 'b111010111;
    h_1 = 'b111001010;
    h_2 = 'b110110101;
    h_3 = 'b110100100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111011001;
    x_1 = 'b111001001;
    x_2 = 'b110111001;
    x_3 = 'b110101010;
    x_4 = 'b110101001;
    x_5 = 'b110100110;
    x_6 = 'b110111010;
    x_7 = 'b111100101;
    x_8 = 'b111000100;
    x_9 = 'b110111111;
    x_10 = 'b110111100;
    x_11 = 'b110110111;
    x_12 = 'b110110000;
    x_13 = 'b110110010;
    x_14 = 'b111011000;
    x_15 = 'b111001111;
    x_16 = 'b111001010;
    x_17 = 'b111000110;
    x_18 = 'b111001100;
    x_19 = 'b111001011;
    x_20 = 'b111000101;
    x_21 = 'b111101010;
    x_22 = 'b111011011;
    x_23 = 'b111011011;
    x_24 = 'b111111100;
    x_25 = 'b111111011;
    x_26 = 'b111000010;
    x_27 = 'b110111111;
    x_28 = 'b111010101;
    x_29 = 'b111110110;
    x_30 = 'b111101101;
    x_31 = 'b111000001;
    x_32 = 'b111000100;
    x_33 = 'b110111001;
    x_34 = 'b110111000;
    x_35 = 'b111000011;
    x_36 = 'b110111101;
    x_37 = 'b111110011;
    x_38 = 'b111110011;
    x_39 = 'b111000111;
    x_40 = 'b111110111;
    x_41 = 'b111000001;
    x_42 = 'b111110101;
    x_43 = 'b111001101;
    x_44 = 'b111110111;
    x_45 = 'b111110100;
    x_46 = 'b111110010;
    x_47 = 'b111101010;
    x_48 = 'b111100111;
    x_49 = 'b111101010;
    x_50 = 'b111100111;
    x_51 = 'b111110010;
    x_52 = 'b111110010;
    x_53 = 'b111110111;
    x_54 = 'b111110010;
    x_55 = 'b111111010;
    x_56 = 'b111101110;
    x_57 = 'b000000000;
    x_58 = 'b111111101;
    x_59 = 'b111110101;
    x_60 = 'b111111000;
    x_61 = 'b111110001;
    x_62 = 'b111111001;
    x_63 = 'b111101111;

    h_0 = 'b111011001;
    h_1 = 'b111001001;
    h_2 = 'b110111001;
    h_3 = 'b110101010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111101101;
    x_1 = 'b111100001;
    x_2 = 'b111010000;
    x_3 = 'b111000000;
    x_4 = 'b111000000;
    x_5 = 'b110111110;
    x_6 = 'b111010110;
    x_7 = 'b000000110;
    x_8 = 'b111011111;
    x_9 = 'b111011110;
    x_10 = 'b111011010;
    x_11 = 'b111001100;
    x_12 = 'b111001011;
    x_13 = 'b111001001;
    x_14 = 'b111110110;
    x_15 = 'b111101011;
    x_16 = 'b111100101;
    x_17 = 'b111100011;
    x_18 = 'b111100101;
    x_19 = 'b111100010;
    x_20 = 'b111010111;
    x_21 = 'b111110000;
    x_22 = 'b111100010;
    x_23 = 'b111100001;
    x_24 = 'b000000011;
    x_25 = 'b000000010;
    x_26 = 'b111001010;
    x_27 = 'b111001000;
    x_28 = 'b111011011;
    x_29 = 'b111111111;
    x_30 = 'b111110101;
    x_31 = 'b111001011;
    x_32 = 'b111010011;
    x_33 = 'b111001000;
    x_34 = 'b111000101;
    x_35 = 'b111010001;
    x_36 = 'b111001110;
    x_37 = 'b111111110;
    x_38 = 'b000000010;
    x_39 = 'b111010110;
    x_40 = 'b111111000;
    x_41 = 'b111100000;
    x_42 = 'b111110111;
    x_43 = 'b000000000;
    x_44 = 'b111111110;
    x_45 = 'b111111000;
    x_46 = 'b111101101;
    x_47 = 'b111101110;
    x_48 = 'b111101101;
    x_49 = 'b111110000;
    x_50 = 'b111110011;
    x_51 = 'b111111000;
    x_52 = 'b111110111;
    x_53 = 'b111111000;
    x_54 = 'b111101111;
    x_55 = 'b111110100;
    x_56 = 'b111101011;
    x_57 = 'b000000001;
    x_58 = 'b111111001;
    x_59 = 'b111101010;
    x_60 = 'b111110101;
    x_61 = 'b111110001;
    x_62 = 'b111111011;
    x_63 = 'b111101110;

    h_0 = 'b111101101;
    h_1 = 'b111100001;
    h_2 = 'b111010000;
    h_3 = 'b111000000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111111101;
    x_1 = 'b111110000;
    x_2 = 'b111100001;
    x_3 = 'b111010110;
    x_4 = 'b111010110;
    x_5 = 'b111010010;
    x_6 = 'b111101001;
    x_7 = 'b000001101;
    x_8 = 'b111100110;
    x_9 = 'b111101100;
    x_10 = 'b111101100;
    x_11 = 'b111011011;
    x_12 = 'b111011101;
    x_13 = 'b111011001;
    x_14 = 'b111101110;
    x_15 = 'b111101101;
    x_16 = 'b111101101;
    x_17 = 'b111101100;
    x_18 = 'b111101101;
    x_19 = 'b111101001;
    x_20 = 'b111011111;
    x_21 = 'b111110100;
    x_22 = 'b111101000;
    x_23 = 'b111101001;
    x_24 = 'b000000110;
    x_25 = 'b000000101;
    x_26 = 'b111010100;
    x_27 = 'b111010011;
    x_28 = 'b111100101;
    x_29 = 'b000000010;
    x_30 = 'b111111110;
    x_31 = 'b111011001;
    x_32 = 'b111011100;
    x_33 = 'b111010100;
    x_34 = 'b111010001;
    x_35 = 'b111011100;
    x_36 = 'b111011100;
    x_37 = 'b000000111;
    x_38 = 'b000000001;
    x_39 = 'b111100001;
    x_40 = 'b111110011;
    x_41 = 'b111011101;
    x_42 = 'b000001111;
    x_43 = 'b111111011;
    x_44 = 'b000000101;
    x_45 = 'b111101111;
    x_46 = 'b111101101;
    x_47 = 'b111101010;
    x_48 = 'b111101001;
    x_49 = 'b111101110;
    x_50 = 'b111110011;
    x_51 = 'b111110110;
    x_52 = 'b111110011;
    x_53 = 'b111110011;
    x_54 = 'b111100000;
    x_55 = 'b111101100;
    x_56 = 'b111100011;
    x_57 = 'b111111010;
    x_58 = 'b111101101;
    x_59 = 'b111011110;
    x_60 = 'b111101101;
    x_61 = 'b111101001;
    x_62 = 'b111110001;
    x_63 = 'b111100111;

    h_0 = 'b111111101;
    h_1 = 'b111110000;
    h_2 = 'b111100001;
    h_3 = 'b111010110;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111111011;
    x_1 = 'b111101111;
    x_2 = 'b111100010;
    x_3 = 'b111011010;
    x_4 = 'b111011001;
    x_5 = 'b111010100;
    x_6 = 'b111100110;
    x_7 = 'b000001000;
    x_8 = 'b111100100;
    x_9 = 'b111101000;
    x_10 = 'b111100110;
    x_11 = 'b111010110;
    x_12 = 'b111011011;
    x_13 = 'b111011100;
    x_14 = 'b111101101;
    x_15 = 'b111101001;
    x_16 = 'b111101001;
    x_17 = 'b111100101;
    x_18 = 'b111100101;
    x_19 = 'b111100001;
    x_20 = 'b111011000;
    x_21 = 'b111110101;
    x_22 = 'b111101001;
    x_23 = 'b111101100;
    x_24 = 'b000000110;
    x_25 = 'b000000101;
    x_26 = 'b111010100;
    x_27 = 'b111010111;
    x_28 = 'b111101000;
    x_29 = 'b000000011;
    x_30 = 'b111111111;
    x_31 = 'b111011010;
    x_32 = 'b111011011;
    x_33 = 'b111010010;
    x_34 = 'b111010001;
    x_35 = 'b111011101;
    x_36 = 'b111011100;
    x_37 = 'b000001101;
    x_38 = 'b111111111;
    x_39 = 'b111100010;
    x_40 = 'b000001011;
    x_41 = 'b111011000;
    x_42 = 'b000001001;
    x_43 = 'b111001011;
    x_44 = 'b000010100;
    x_45 = 'b111011001;
    x_46 = 'b111110001;
    x_47 = 'b111101011;
    x_48 = 'b111100111;
    x_49 = 'b111101000;
    x_50 = 'b111100111;
    x_51 = 'b111100101;
    x_52 = 'b111100001;
    x_53 = 'b111100000;
    x_54 = 'b111010001;
    x_55 = 'b111100110;
    x_56 = 'b111011101;
    x_57 = 'b111101110;
    x_58 = 'b111011000;
    x_59 = 'b111001111;
    x_60 = 'b111100010;
    x_61 = 'b111011010;
    x_62 = 'b111011011;
    x_63 = 'b111011110;

    h_0 = 'b111111011;
    h_1 = 'b111101111;
    h_2 = 'b111100010;
    h_3 = 'b111011010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111111010;
    x_1 = 'b111101100;
    x_2 = 'b111011100;
    x_3 = 'b111010001;
    x_4 = 'b111010001;
    x_5 = 'b111001101;
    x_6 = 'b111011101;
    x_7 = 'b000000111;
    x_8 = 'b111100110;
    x_9 = 'b111100010;
    x_10 = 'b111011100;
    x_11 = 'b111001010;
    x_12 = 'b111010100;
    x_13 = 'b111010000;
    x_14 = 'b111111000;
    x_15 = 'b111101000;
    x_16 = 'b111100010;
    x_17 = 'b111011010;
    x_18 = 'b111011011;
    x_19 = 'b111010111;
    x_20 = 'b111001111;
    x_21 = 'b111110100;
    x_22 = 'b111100111;
    x_23 = 'b111100111;
    x_24 = 'b000000110;
    x_25 = 'b000000101;
    x_26 = 'b111010000;
    x_27 = 'b111010001;
    x_28 = 'b111100011;
    x_29 = 'b000000100;
    x_30 = 'b111111010;
    x_31 = 'b111010010;
    x_32 = 'b111010111;
    x_33 = 'b111001100;
    x_34 = 'b111001010;
    x_35 = 'b111010111;
    x_36 = 'b111010001;
    x_37 = 'b000000001;
    x_38 = 'b000001001;
    x_39 = 'b111001110;
    x_40 = 'b000010110;
    x_41 = 'b110100110;
    x_42 = 'b000010001;
    x_43 = 'b111110111;
    x_44 = 'b000010011;
    x_45 = 'b111100100;
    x_46 = 'b111101111;
    x_47 = 'b111101001;
    x_48 = 'b111100011;
    x_49 = 'b111100000;
    x_50 = 'b111011101;
    x_51 = 'b111011000;
    x_52 = 'b111011000;
    x_53 = 'b111011100;
    x_54 = 'b111010111;
    x_55 = 'b111100010;
    x_56 = 'b111011010;
    x_57 = 'b111100011;
    x_58 = 'b111010000;
    x_59 = 'b111001111;
    x_60 = 'b111011001;
    x_61 = 'b111001111;
    x_62 = 'b111001001;
    x_63 = 'b111011010;

    h_0 = 'b111111010;
    h_1 = 'b111101100;
    h_2 = 'b111011100;
    h_3 = 'b111010001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111110111;
    x_1 = 'b111100111;
    x_2 = 'b111010110;
    x_3 = 'b111001110;
    x_4 = 'b111001101;
    x_5 = 'b111001010;
    x_6 = 'b111010011;
    x_7 = 'b000000001;
    x_8 = 'b111100000;
    x_9 = 'b111011011;
    x_10 = 'b111011000;
    x_11 = 'b111001001;
    x_12 = 'b111010000;
    x_13 = 'b111000000;
    x_14 = 'b111110010;
    x_15 = 'b111100011;
    x_16 = 'b111011100;
    x_17 = 'b111010100;
    x_18 = 'b111011000;
    x_19 = 'b111010100;
    x_20 = 'b111001101;
    x_21 = 'b111110000;
    x_22 = 'b111100011;
    x_23 = 'b111100010;
    x_24 = 'b000000100;
    x_25 = 'b000000100;
    x_26 = 'b111001110;
    x_27 = 'b111001101;
    x_28 = 'b111100001;
    x_29 = 'b000000100;
    x_30 = 'b111111011;
    x_31 = 'b111010001;
    x_32 = 'b111010001;
    x_33 = 'b111001001;
    x_34 = 'b111000111;
    x_35 = 'b111010011;
    x_36 = 'b111001110;
    x_37 = 'b111111010;
    x_38 = 'b000000001;
    x_39 = 'b111001011;
    x_40 = 'b000001001;
    x_41 = 'b111000100;
    x_42 = 'b000001100;
    x_43 = 'b111110101;
    x_44 = 'b000000101;
    x_45 = 'b111110010;
    x_46 = 'b111110101;
    x_47 = 'b111101010;
    x_48 = 'b111100010;
    x_49 = 'b111011110;
    x_50 = 'b111011100;
    x_51 = 'b111011011;
    x_52 = 'b111011111;
    x_53 = 'b111100111;
    x_54 = 'b111101001;
    x_55 = 'b111100011;
    x_56 = 'b111011100;
    x_57 = 'b111100110;
    x_58 = 'b111100001;
    x_59 = 'b111100110;
    x_60 = 'b111010111;
    x_61 = 'b111010001;
    x_62 = 'b111001011;
    x_63 = 'b111100011;

    h_0 = 'b111110111;
    h_1 = 'b111100111;
    h_2 = 'b111010110;
    h_3 = 'b111001110;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111110110;
    x_1 = 'b111011111;
    x_2 = 'b111010000;
    x_3 = 'b111000111;
    x_4 = 'b111001000;
    x_5 = 'b111001010;
    x_6 = 'b111011001;
    x_7 = 'b000000000;
    x_8 = 'b111011010;
    x_9 = 'b111011000;
    x_10 = 'b111010101;
    x_11 = 'b111001001;
    x_12 = 'b111010010;
    x_13 = 'b111001100;
    x_14 = 'b111110001;
    x_15 = 'b111100100;
    x_16 = 'b111011100;
    x_17 = 'b111010101;
    x_18 = 'b111011011;
    x_19 = 'b111011001;
    x_20 = 'b111010011;
    x_21 = 'b111101100;
    x_22 = 'b111100001;
    x_23 = 'b111100000;
    x_24 = 'b000000001;
    x_25 = 'b000000000;
    x_26 = 'b111001100;
    x_27 = 'b111001100;
    x_28 = 'b111011111;
    x_29 = 'b000000011;
    x_30 = 'b111110110;
    x_31 = 'b111001111;
    x_32 = 'b111001101;
    x_33 = 'b111001000;
    x_34 = 'b111000111;
    x_35 = 'b111010010;
    x_36 = 'b111010011;
    x_37 = 'b111111001;
    x_38 = 'b111111011;
    x_39 = 'b111011001;
    x_40 = 'b111111101;
    x_41 = 'b111011111;
    x_42 = 'b111110101;
    x_43 = 'b111011101;
    x_44 = 'b000000010;
    x_45 = 'b111101001;
    x_46 = 'b111110011;
    x_47 = 'b111110000;
    x_48 = 'b111100111;
    x_49 = 'b111101001;
    x_50 = 'b111100011;
    x_51 = 'b111101100;
    x_52 = 'b111110000;
    x_53 = 'b111111011;
    x_54 = 'b111111100;
    x_55 = 'b111110000;
    x_56 = 'b111101010;
    x_57 = 'b111110101;
    x_58 = 'b111111111;
    x_59 = 'b000001100;
    x_60 = 'b111100100;
    x_61 = 'b111100110;
    x_62 = 'b111101001;
    x_63 = 'b111111001;

    h_0 = 'b111110110;
    h_1 = 'b111011111;
    h_2 = 'b111010000;
    h_3 = 'b111000111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111101111;
    x_1 = 'b111011011;
    x_2 = 'b111001101;
    x_3 = 'b111000011;
    x_4 = 'b111001000;
    x_5 = 'b111001001;
    x_6 = 'b111011000;
    x_7 = 'b111111011;
    x_8 = 'b111011010;
    x_9 = 'b111011000;
    x_10 = 'b111010111;
    x_11 = 'b111001011;
    x_12 = 'b111010101;
    x_13 = 'b111010000;
    x_14 = 'b111110000;
    x_15 = 'b111101000;
    x_16 = 'b111100010;
    x_17 = 'b111010111;
    x_18 = 'b111100011;
    x_19 = 'b111100001;
    x_20 = 'b111011010;
    x_21 = 'b111101010;
    x_22 = 'b111011100;
    x_23 = 'b111011011;
    x_24 = 'b111111011;
    x_25 = 'b111111011;
    x_26 = 'b111000101;
    x_27 = 'b111000101;
    x_28 = 'b111011001;
    x_29 = 'b111110111;
    x_30 = 'b111101110;
    x_31 = 'b111000111;
    x_32 = 'b111001000;
    x_33 = 'b111000010;
    x_34 = 'b111000010;
    x_35 = 'b111001011;
    x_36 = 'b111001010;
    x_37 = 'b111101110;
    x_38 = 'b111111010;
    x_39 = 'b111001011;
    x_40 = 'b111110011;
    x_41 = 'b110110111;
    x_42 = 'b111111000;
    x_43 = 'b111101010;
    x_44 = 'b000000001;
    x_45 = 'b111111010;
    x_46 = 'b111110010;
    x_47 = 'b111110101;
    x_48 = 'b111110000;
    x_49 = 'b111110010;
    x_50 = 'b111101010;
    x_51 = 'b111111101;
    x_52 = 'b000000010;
    x_53 = 'b000010010;
    x_54 = 'b000011001;
    x_55 = 'b111111110;
    x_56 = 'b111110111;
    x_57 = 'b000000011;
    x_58 = 'b000011111;
    x_59 = 'b000110100;
    x_60 = 'b111111001;
    x_61 = 'b000000111;
    x_62 = 'b000011000;
    x_63 = 'b000010100;

    h_0 = 'b111101111;
    h_1 = 'b111011011;
    h_2 = 'b111001101;
    h_3 = 'b111000011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111101110;
    x_1 = 'b111100000;
    x_2 = 'b111001101;
    x_3 = 'b111000011;
    x_4 = 'b111000110;
    x_5 = 'b111000101;
    x_6 = 'b111001101;
    x_7 = 'b111111010;
    x_8 = 'b111011111;
    x_9 = 'b111011011;
    x_10 = 'b111011010;
    x_11 = 'b111001110;
    x_12 = 'b111010011;
    x_13 = 'b111000101;
    x_14 = 'b111110100;
    x_15 = 'b111101100;
    x_16 = 'b111100111;
    x_17 = 'b111011010;
    x_18 = 'b111100111;
    x_19 = 'b111100111;
    x_20 = 'b111100000;
    x_21 = 'b111101111;
    x_22 = 'b111100001;
    x_23 = 'b111100001;
    x_24 = 'b000000001;
    x_25 = 'b000000000;
    x_26 = 'b111001101;
    x_27 = 'b111001011;
    x_28 = 'b111011101;
    x_29 = 'b000000000;
    x_30 = 'b111110101;
    x_31 = 'b111010000;
    x_32 = 'b111010001;
    x_33 = 'b111000111;
    x_34 = 'b111000110;
    x_35 = 'b111010010;
    x_36 = 'b111001010;
    x_37 = 'b111101011;
    x_38 = 'b000000100;
    x_39 = 'b111000110;
    x_40 = 'b000000101;
    x_41 = 'b110111000;
    x_42 = 'b000010101;
    x_43 = 'b111100001;
    x_44 = 'b000010101;
    x_45 = 'b000010000;
    x_46 = 'b000000011;
    x_47 = 'b000000001;
    x_48 = 'b111111001;
    x_49 = 'b111110100;
    x_50 = 'b111101011;
    x_51 = 'b000000001;
    x_52 = 'b000001010;
    x_53 = 'b000011110;
    x_54 = 'b000101000;
    x_55 = 'b000001111;
    x_56 = 'b000000010;
    x_57 = 'b000000011;
    x_58 = 'b000101001;
    x_59 = 'b001000100;
    x_60 = 'b000001110;
    x_61 = 'b000100000;
    x_62 = 'b000111101;
    x_63 = 'b000101001;

    h_0 = 'b111101110;
    h_1 = 'b111100000;
    h_2 = 'b111001101;
    h_3 = 'b111000011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111111101;
    x_1 = 'b111110000;
    x_2 = 'b111011010;
    x_3 = 'b111001111;
    x_4 = 'b111001011;
    x_5 = 'b111001001;
    x_6 = 'b111010010;
    x_7 = 'b000001000;
    x_8 = 'b111101010;
    x_9 = 'b111100010;
    x_10 = 'b111011111;
    x_11 = 'b111010001;
    x_12 = 'b111011001;
    x_13 = 'b111001111;
    x_14 = 'b000000000;
    x_15 = 'b111110000;
    x_16 = 'b111101001;
    x_17 = 'b111011101;
    x_18 = 'b111101001;
    x_19 = 'b111101100;
    x_20 = 'b111101010;
    x_21 = 'b111110001;
    x_22 = 'b111100000;
    x_23 = 'b111011111;
    x_24 = 'b000000100;
    x_25 = 'b000000010;
    x_26 = 'b111010000;
    x_27 = 'b111001000;
    x_28 = 'b111011000;
    x_29 = 'b000000101;
    x_30 = 'b111111011;
    x_31 = 'b111001110;
    x_32 = 'b111010111;
    x_33 = 'b111001100;
    x_34 = 'b111000110;
    x_35 = 'b111010010;
    x_36 = 'b111000100;
    x_37 = 'b111101000;
    x_38 = 'b000000110;
    x_39 = 'b111000111;
    x_40 = 'b000010011;
    x_41 = 'b111001001;
    x_42 = 'b000010010;
    x_43 = 'b111011111;
    x_44 = 'b000010110;
    x_45 = 'b111111100;
    x_46 = 'b000001010;
    x_47 = 'b000000011;
    x_48 = 'b111111000;
    x_49 = 'b111110010;
    x_50 = 'b111101000;
    x_51 = 'b000000001;
    x_52 = 'b000001011;
    x_53 = 'b000011110;
    x_54 = 'b000100101;
    x_55 = 'b000010101;
    x_56 = 'b000000100;
    x_57 = 'b000000010;
    x_58 = 'b000101011;
    x_59 = 'b001000111;
    x_60 = 'b000011011;
    x_61 = 'b000100111;
    x_62 = 'b001001010;
    x_63 = 'b000101011;

    h_0 = 'b111111101;
    h_1 = 'b111110000;
    h_2 = 'b111011010;
    h_3 = 'b111001111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111111101;
    x_1 = 'b111101011;
    x_2 = 'b111010111;
    x_3 = 'b111001010;
    x_4 = 'b111000101;
    x_5 = 'b111000010;
    x_6 = 'b111001000;
    x_7 = 'b000000110;
    x_8 = 'b111100110;
    x_9 = 'b111100000;
    x_10 = 'b111011111;
    x_11 = 'b111001101;
    x_12 = 'b111010111;
    x_13 = 'b111010000;
    x_14 = 'b000000001;
    x_15 = 'b111101101;
    x_16 = 'b111101000;
    x_17 = 'b111011111;
    x_18 = 'b111101101;
    x_19 = 'b111110000;
    x_20 = 'b111110000;
    x_21 = 'b111101000;
    x_22 = 'b111010110;
    x_23 = 'b111010100;
    x_24 = 'b111111101;
    x_25 = 'b111111011;
    x_26 = 'b111000101;
    x_27 = 'b110111011;
    x_28 = 'b111001110;
    x_29 = 'b000001010;
    x_30 = 'b111110010;
    x_31 = 'b111000111;
    x_32 = 'b111001111;
    x_33 = 'b111000011;
    x_34 = 'b110111011;
    x_35 = 'b111000110;
    x_36 = 'b110111100;
    x_37 = 'b111100111;
    x_38 = 'b000001100;
    x_39 = 'b110111111;
    x_40 = 'b000010101;
    x_41 = 'b111000110;
    x_42 = 'b000001110;
    x_43 = 'b000010000;
    x_44 = 'b000100000;
    x_45 = 'b000001110;
    x_46 = 'b000011011;
    x_47 = 'b000010010;
    x_48 = 'b000000100;
    x_49 = 'b111111111;
    x_50 = 'b111110110;
    x_51 = 'b000001111;
    x_52 = 'b000011000;
    x_53 = 'b000101100;
    x_54 = 'b000110011;
    x_55 = 'b000101001;
    x_56 = 'b000010110;
    x_57 = 'b000001111;
    x_58 = 'b000110101;
    x_59 = 'b001001011;
    x_60 = 'b000100110;
    x_61 = 'b000101000;
    x_62 = 'b001001001;
    x_63 = 'b000101101;

    h_0 = 'b111111101;
    h_1 = 'b111101011;
    h_2 = 'b111010111;
    h_3 = 'b111001010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000000101;
    x_1 = 'b111110010;
    x_2 = 'b111011100;
    x_3 = 'b111000110;
    x_4 = 'b111000100;
    x_5 = 'b111000010;
    x_6 = 'b111001111;
    x_7 = 'b000010101;
    x_8 = 'b111110011;
    x_9 = 'b111101101;
    x_10 = 'b111101010;
    x_11 = 'b111010100;
    x_12 = 'b111011011;
    x_13 = 'b111011101;
    x_14 = 'b000010011;
    x_15 = 'b000000010;
    x_16 = 'b111111010;
    x_17 = 'b111101110;
    x_18 = 'b111111010;
    x_19 = 'b111111100;
    x_20 = 'b111111110;
    x_21 = 'b111101011;
    x_22 = 'b111011000;
    x_23 = 'b111011000;
    x_24 = 'b111111111;
    x_25 = 'b111111101;
    x_26 = 'b111000110;
    x_27 = 'b110111100;
    x_28 = 'b111010011;
    x_29 = 'b000001001;
    x_30 = 'b111110110;
    x_31 = 'b111000111;
    x_32 = 'b111010010;
    x_33 = 'b111000010;
    x_34 = 'b110111010;
    x_35 = 'b111000110;
    x_36 = 'b111000000;
    x_37 = 'b111110000;
    x_38 = 'b000010001;
    x_39 = 'b111001001;
    x_40 = 'b000001111;
    x_41 = 'b111001001;
    x_42 = 'b000100100;
    x_43 = 'b111110110;
    x_44 = 'b000110110;
    x_45 = 'b000011011;
    x_46 = 'b000110101;
    x_47 = 'b000100010;
    x_48 = 'b000001111;
    x_49 = 'b000001010;
    x_50 = 'b111111111;
    x_51 = 'b000010001;
    x_52 = 'b000010110;
    x_53 = 'b000101000;
    x_54 = 'b000101110;
    x_55 = 'b000111000;
    x_56 = 'b000100001;
    x_57 = 'b000010101;
    x_58 = 'b000101111;
    x_59 = 'b001000001;
    x_60 = 'b000110010;
    x_61 = 'b000101011;
    x_62 = 'b001000011;
    x_63 = 'b000111000;

    h_0 = 'b000000101;
    h_1 = 'b111110010;
    h_2 = 'b111011100;
    h_3 = 'b111000110;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000000001;
    x_1 = 'b111110111;
    x_2 = 'b111100001;
    x_3 = 'b111001011;
    x_4 = 'b111000001;
    x_5 = 'b110111010;
    x_6 = 'b111001010;
    x_7 = 'b000010100;
    x_8 = 'b111110101;
    x_9 = 'b111110010;
    x_10 = 'b111101011;
    x_11 = 'b111001100;
    x_12 = 'b111001011;
    x_13 = 'b111010000;
    x_14 = 'b000011100;
    x_15 = 'b000000101;
    x_16 = 'b111111100;
    x_17 = 'b111101111;
    x_18 = 'b111110101;
    x_19 = 'b111110001;
    x_20 = 'b111101101;
    x_21 = 'b111101111;
    x_22 = 'b111011100;
    x_23 = 'b111011011;
    x_24 = 'b000000100;
    x_25 = 'b000000010;
    x_26 = 'b111001010;
    x_27 = 'b110111110;
    x_28 = 'b111001111;
    x_29 = 'b000001111;
    x_30 = 'b111111010;
    x_31 = 'b111001010;
    x_32 = 'b111011001;
    x_33 = 'b111001010;
    x_34 = 'b111000000;
    x_35 = 'b111001011;
    x_36 = 'b111000001;
    x_37 = 'b111110000;
    x_38 = 'b000010010;
    x_39 = 'b111001010;
    x_40 = 'b000011011;
    x_41 = 'b111011100;
    x_42 = 'b000101100;
    x_43 = 'b111101011;
    x_44 = 'b000110110;
    x_45 = 'b000000101;
    x_46 = 'b000110000;
    x_47 = 'b000100001;
    x_48 = 'b000001101;
    x_49 = 'b000001001;
    x_50 = 'b111111011;
    x_51 = 'b000000111;
    x_52 = 'b000001011;
    x_53 = 'b000010111;
    x_54 = 'b000011100;
    x_55 = 'b000110111;
    x_56 = 'b000100000;
    x_57 = 'b000010001;
    x_58 = 'b000011110;
    x_59 = 'b000100011;
    x_60 = 'b000110110;
    x_61 = 'b000100011;
    x_62 = 'b000110100;
    x_63 = 'b000110100;

    h_0 = 'b000000001;
    h_1 = 'b111110111;
    h_2 = 'b111100001;
    h_3 = 'b111001011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000000111;
    x_1 = 'b111111011;
    x_2 = 'b111100100;
    x_3 = 'b111001111;
    x_4 = 'b111000111;
    x_5 = 'b110111101;
    x_6 = 'b111001011;
    x_7 = 'b000010111;
    x_8 = 'b111110110;
    x_9 = 'b111110001;
    x_10 = 'b111100101;
    x_11 = 'b111001100;
    x_12 = 'b111000111;
    x_13 = 'b111010000;
    x_14 = 'b000010111;
    x_15 = 'b000000011;
    x_16 = 'b111111001;
    x_17 = 'b111101101;
    x_18 = 'b111110001;
    x_19 = 'b111101001;
    x_20 = 'b111100101;
    x_21 = 'b111110101;
    x_22 = 'b111100011;
    x_23 = 'b111100011;
    x_24 = 'b000001000;
    x_25 = 'b000000111;
    x_26 = 'b111010001;
    x_27 = 'b111000111;
    x_28 = 'b111011101;
    x_29 = 'b000010100;
    x_30 = 'b111111011;
    x_31 = 'b111010100;
    x_32 = 'b111011010;
    x_33 = 'b111001101;
    x_34 = 'b111000111;
    x_35 = 'b111010000;
    x_36 = 'b111000111;
    x_37 = 'b111110100;
    x_38 = 'b000011000;
    x_39 = 'b111010101;
    x_40 = 'b000101010;
    x_41 = 'b111101011;
    x_42 = 'b000101110;
    x_43 = 'b111100100;
    x_44 = 'b000110110;
    x_45 = 'b111111110;
    x_46 = 'b000101010;
    x_47 = 'b000011011;
    x_48 = 'b000001010;
    x_49 = 'b000001000;
    x_50 = 'b111111101;
    x_51 = 'b000000101;
    x_52 = 'b000000110;
    x_53 = 'b000001100;
    x_54 = 'b000001101;
    x_55 = 'b000110000;
    x_56 = 'b000011011;
    x_57 = 'b000010000;
    x_58 = 'b000010110;
    x_59 = 'b000010001;
    x_60 = 'b000101111;
    x_61 = 'b000010110;
    x_62 = 'b000100010;
    x_63 = 'b000101011;

    h_0 = 'b000000111;
    h_1 = 'b111111011;
    h_2 = 'b111100100;
    h_3 = 'b111001111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111001010;
    x_1 = 'b111011110;
    x_2 = 'b111100001;
    x_3 = 'b111110101;
    x_4 = 'b111111001;
    x_5 = 'b111111000;
    x_6 = 'b111101000;
    x_7 = 'b111011011;
    x_8 = 'b111101100;
    x_9 = 'b111110011;
    x_10 = 'b111111011;
    x_11 = 'b000000000;
    x_12 = 'b000000011;
    x_13 = 'b111111001;
    x_14 = 'b111101100;
    x_15 = 'b111110100;
    x_16 = 'b111111000;
    x_17 = 'b000000100;
    x_18 = 'b000000101;
    x_19 = 'b000001001;
    x_20 = 'b000001100;
    x_21 = 'b111001100;
    x_22 = 'b111001001;
    x_23 = 'b111010010;
    x_24 = 'b111001000;
    x_25 = 'b111001001;
    x_26 = 'b111010110;
    x_27 = 'b111011001;
    x_28 = 'b111010110;
    x_29 = 'b111000101;
    x_30 = 'b111010011;
    x_31 = 'b111011011;
    x_32 = 'b111011101;
    x_33 = 'b111100011;
    x_34 = 'b111101010;
    x_35 = 'b111101001;
    x_36 = 'b111101000;
    x_37 = 'b111101010;
    x_38 = 'b111001010;
    x_39 = 'b111101011;
    x_40 = 'b111001110;
    x_41 = 'b000000000;
    x_42 = 'b110111110;
    x_43 = 'b000000110;
    x_44 = 'b111100001;
    x_45 = 'b111111100;
    x_46 = 'b111111101;
    x_47 = 'b111111100;
    x_48 = 'b000000011;
    x_49 = 'b000000101;
    x_50 = 'b000000110;
    x_51 = 'b000010010;
    x_52 = 'b000001011;
    x_53 = 'b000010001;
    x_54 = 'b000001011;
    x_55 = 'b000001101;
    x_56 = 'b000001101;
    x_57 = 'b000011100;
    x_58 = 'b000011100;
    x_59 = 'b000010110;
    x_60 = 'b000011101;
    x_61 = 'b000100111;
    x_62 = 'b000001011;
    x_63 = 'b000011010;

    h_0 = 'b111001010;
    h_1 = 'b111011110;
    h_2 = 'b111100001;
    h_3 = 'b111110101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111001110;
    x_1 = 'b111100100;
    x_2 = 'b111100111;
    x_3 = 'b111110101;
    x_4 = 'b111111011;
    x_5 = 'b111111110;
    x_6 = 'b111111000;
    x_7 = 'b111100010;
    x_8 = 'b111110001;
    x_9 = 'b111110100;
    x_10 = 'b111110110;
    x_11 = 'b111111111;
    x_12 = 'b000000101;
    x_13 = 'b000000101;
    x_14 = 'b111101011;
    x_15 = 'b111110011;
    x_16 = 'b111110110;
    x_17 = 'b111111100;
    x_18 = 'b111111000;
    x_19 = 'b111111111;
    x_20 = 'b000000101;
    x_21 = 'b111001001;
    x_22 = 'b111001100;
    x_23 = 'b111010111;
    x_24 = 'b111000111;
    x_25 = 'b111001000;
    x_26 = 'b111010111;
    x_27 = 'b111011111;
    x_28 = 'b111011101;
    x_29 = 'b111000111;
    x_30 = 'b111011001;
    x_31 = 'b111011111;
    x_32 = 'b111011101;
    x_33 = 'b111100100;
    x_34 = 'b111101100;
    x_35 = 'b111101011;
    x_36 = 'b111110010;
    x_37 = 'b111110000;
    x_38 = 'b111001100;
    x_39 = 'b111111100;
    x_40 = 'b111010000;
    x_41 = 'b000101001;
    x_42 = 'b110111111;
    x_43 = 'b111011111;
    x_44 = 'b111011000;
    x_45 = 'b111101011;
    x_46 = 'b111110011;
    x_47 = 'b111111001;
    x_48 = 'b000000011;
    x_49 = 'b000000001;
    x_50 = 'b111111110;
    x_51 = 'b000001000;
    x_52 = 'b000000010;
    x_53 = 'b000001011;
    x_54 = 'b000000110;
    x_55 = 'b000001100;
    x_56 = 'b000001011;
    x_57 = 'b000011001;
    x_58 = 'b000011000;
    x_59 = 'b000010101;
    x_60 = 'b000011001;
    x_61 = 'b000100011;
    x_62 = 'b000000101;
    x_63 = 'b000010111;

    h_0 = 'b111001110;
    h_1 = 'b111100100;
    h_2 = 'b111100111;
    h_3 = 'b111110101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111010101;
    x_1 = 'b111101011;
    x_2 = 'b111101011;
    x_3 = 'b111110100;
    x_4 = 'b111111001;
    x_5 = 'b111111110;
    x_6 = 'b000000000;
    x_7 = 'b111101011;
    x_8 = 'b111110111;
    x_9 = 'b111110010;
    x_10 = 'b111101111;
    x_11 = 'b111111000;
    x_12 = 'b000000010;
    x_13 = 'b000001010;
    x_14 = 'b111110000;
    x_15 = 'b111110111;
    x_16 = 'b111110100;
    x_17 = 'b111111000;
    x_18 = 'b111110000;
    x_19 = 'b111111000;
    x_20 = 'b000000110;
    x_21 = 'b111010001;
    x_22 = 'b111010001;
    x_23 = 'b111011010;
    x_24 = 'b111001111;
    x_25 = 'b111001111;
    x_26 = 'b111011011;
    x_27 = 'b111100001;
    x_28 = 'b111011101;
    x_29 = 'b111010001;
    x_30 = 'b111011010;
    x_31 = 'b111100011;
    x_32 = 'b111100011;
    x_33 = 'b111100111;
    x_34 = 'b111101110;
    x_35 = 'b111101110;
    x_36 = 'b111110010;
    x_37 = 'b111101110;
    x_38 = 'b111011011;
    x_39 = 'b111111000;
    x_40 = 'b111100000;
    x_41 = 'b000010011;
    x_42 = 'b110111100;
    x_43 = 'b000000110;
    x_44 = 'b111100100;
    x_45 = 'b111111000;
    x_46 = 'b111111111;
    x_47 = 'b000000001;
    x_48 = 'b000001001;
    x_49 = 'b000000100;
    x_50 = 'b111111111;
    x_51 = 'b000000101;
    x_52 = 'b000000000;
    x_53 = 'b000001110;
    x_54 = 'b000010000;
    x_55 = 'b000001110;
    x_56 = 'b000001101;
    x_57 = 'b000011001;
    x_58 = 'b000011011;
    x_59 = 'b000011001;
    x_60 = 'b000010111;
    x_61 = 'b000100001;
    x_62 = 'b000000101;
    x_63 = 'b000011000;

    h_0 = 'b111010101;
    h_1 = 'b111101011;
    h_2 = 'b111101011;
    h_3 = 'b111110100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111100010;
    x_1 = 'b111110010;
    x_2 = 'b111101111;
    x_3 = 'b111110101;
    x_4 = 'b111111000;
    x_5 = 'b111111010;
    x_6 = 'b111111000;
    x_7 = 'b111110101;
    x_8 = 'b111111011;
    x_9 = 'b111110101;
    x_10 = 'b111110100;
    x_11 = 'b111110100;
    x_12 = 'b111111000;
    x_13 = 'b111110011;
    x_14 = 'b111111001;
    x_15 = 'b111111010;
    x_16 = 'b111111000;
    x_17 = 'b111111000;
    x_18 = 'b111101011;
    x_19 = 'b111101111;
    x_20 = 'b111111000;
    x_21 = 'b111010001;
    x_22 = 'b111010000;
    x_23 = 'b111011001;
    x_24 = 'b111010000;
    x_25 = 'b111010001;
    x_26 = 'b111011100;
    x_27 = 'b111100001;
    x_28 = 'b111011101;
    x_29 = 'b111010100;
    x_30 = 'b111011111;
    x_31 = 'b111100010;
    x_32 = 'b111100100;
    x_33 = 'b111100111;
    x_34 = 'b111101111;
    x_35 = 'b111110000;
    x_36 = 'b111101100;
    x_37 = 'b111101101;
    x_38 = 'b111011000;
    x_39 = 'b111100101;
    x_40 = 'b111010111;
    x_41 = 'b111010000;
    x_42 = 'b111000100;
    x_43 = 'b111100111;
    x_44 = 'b111100001;
    x_45 = 'b111101100;
    x_46 = 'b111110110;
    x_47 = 'b111110110;
    x_48 = 'b111111101;
    x_49 = 'b111111011;
    x_50 = 'b111111100;
    x_51 = 'b111111110;
    x_52 = 'b111111001;
    x_53 = 'b000000010;
    x_54 = 'b000000011;
    x_55 = 'b111111001;
    x_56 = 'b111111011;
    x_57 = 'b000001110;
    x_58 = 'b000001110;
    x_59 = 'b000001101;
    x_60 = 'b000001100;
    x_61 = 'b000010111;
    x_62 = 'b111111110;
    x_63 = 'b000001100;

    h_0 = 'b111100010;
    h_1 = 'b111110010;
    h_2 = 'b111101111;
    h_3 = 'b111110101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111011111;
    x_1 = 'b111101111;
    x_2 = 'b111101110;
    x_3 = 'b111110101;
    x_4 = 'b111110111;
    x_5 = 'b111110111;
    x_6 = 'b111101110;
    x_7 = 'b111101100;
    x_8 = 'b111110111;
    x_9 = 'b111110111;
    x_10 = 'b111111001;
    x_11 = 'b111111100;
    x_12 = 'b111110110;
    x_13 = 'b111101111;
    x_14 = 'b111101010;
    x_15 = 'b111110011;
    x_16 = 'b111111001;
    x_17 = 'b111111100;
    x_18 = 'b111110101;
    x_19 = 'b111110110;
    x_20 = 'b111111100;
    x_21 = 'b111001011;
    x_22 = 'b111001001;
    x_23 = 'b111010001;
    x_24 = 'b111001001;
    x_25 = 'b111001011;
    x_26 = 'b111011001;
    x_27 = 'b111011011;
    x_28 = 'b111010111;
    x_29 = 'b111001110;
    x_30 = 'b111100110;
    x_31 = 'b111100100;
    x_32 = 'b111100011;
    x_33 = 'b111101000;
    x_34 = 'b111101111;
    x_35 = 'b111101110;
    x_36 = 'b111101000;
    x_37 = 'b111110000;
    x_38 = 'b111011010;
    x_39 = 'b111101110;
    x_40 = 'b111100101;
    x_41 = 'b000010001;
    x_42 = 'b111000011;
    x_43 = 'b111101000;
    x_44 = 'b111100010;
    x_45 = 'b111110011;
    x_46 = 'b111101101;
    x_47 = 'b111110001;
    x_48 = 'b000000000;
    x_49 = 'b000000001;
    x_50 = 'b000000110;
    x_51 = 'b000001101;
    x_52 = 'b000001010;
    x_53 = 'b000001110;
    x_54 = 'b000001110;
    x_55 = 'b111110100;
    x_56 = 'b111111010;
    x_57 = 'b000010001;
    x_58 = 'b000010111;
    x_59 = 'b000010101;
    x_60 = 'b000000000;
    x_61 = 'b000001100;
    x_62 = 'b111111001;
    x_63 = 'b111111110;

    h_0 = 'b111011111;
    h_1 = 'b111101111;
    h_2 = 'b111101110;
    h_3 = 'b111110101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111100000;
    x_1 = 'b111110000;
    x_2 = 'b111110100;
    x_3 = 'b111111110;
    x_4 = 'b000000010;
    x_5 = 'b000000100;
    x_6 = 'b111111101;
    x_7 = 'b111110010;
    x_8 = 'b111111100;
    x_9 = 'b111111110;
    x_10 = 'b000000000;
    x_11 = 'b000000100;
    x_12 = 'b000001000;
    x_13 = 'b000000101;
    x_14 = 'b111101000;
    x_15 = 'b111110110;
    x_16 = 'b111111101;
    x_17 = 'b000000100;
    x_18 = 'b000000101;
    x_19 = 'b000000110;
    x_20 = 'b000000110;
    x_21 = 'b111001110;
    x_22 = 'b111001111;
    x_23 = 'b111010110;
    x_24 = 'b111001011;
    x_25 = 'b111001100;
    x_26 = 'b111011100;
    x_27 = 'b111011111;
    x_28 = 'b111011010;
    x_29 = 'b111010101;
    x_30 = 'b111011111;
    x_31 = 'b111100011;
    x_32 = 'b111100100;
    x_33 = 'b111101000;
    x_34 = 'b111110010;
    x_35 = 'b111101110;
    x_36 = 'b111101011;
    x_37 = 'b111110011;
    x_38 = 'b111011000;
    x_39 = 'b111101101;
    x_40 = 'b111010000;
    x_41 = 'b111100110;
    x_42 = 'b110111101;
    x_43 = 'b000000100;
    x_44 = 'b111011011;
    x_45 = 'b111100111;
    x_46 = 'b111100110;
    x_47 = 'b111101000;
    x_48 = 'b111110111;
    x_49 = 'b111111000;
    x_50 = 'b000000000;
    x_51 = 'b000001100;
    x_52 = 'b000001000;
    x_53 = 'b000001001;
    x_54 = 'b000000110;
    x_55 = 'b111101110;
    x_56 = 'b111110011;
    x_57 = 'b000001011;
    x_58 = 'b000010000;
    x_59 = 'b000001101;
    x_60 = 'b111110111;
    x_61 = 'b000000101;
    x_62 = 'b111110101;
    x_63 = 'b111110010;

    h_0 = 'b111100000;
    h_1 = 'b111110000;
    h_2 = 'b111110100;
    h_3 = 'b111111110;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111010001;
    x_1 = 'b111100100;
    x_2 = 'b111100111;
    x_3 = 'b111110111;
    x_4 = 'b111111011;
    x_5 = 'b111111100;
    x_6 = 'b111110010;
    x_7 = 'b111011111;
    x_8 = 'b111101110;
    x_9 = 'b111101111;
    x_10 = 'b111110100;
    x_11 = 'b111111111;
    x_12 = 'b000000101;
    x_13 = 'b111111001;
    x_14 = 'b111011111;
    x_15 = 'b111101000;
    x_16 = 'b111110001;
    x_17 = 'b111111100;
    x_18 = 'b000000010;
    x_19 = 'b000000110;
    x_20 = 'b000000010;
    x_21 = 'b111001010;
    x_22 = 'b111001100;
    x_23 = 'b111010110;
    x_24 = 'b111001000;
    x_25 = 'b111001001;
    x_26 = 'b111010111;
    x_27 = 'b111011111;
    x_28 = 'b111011011;
    x_29 = 'b111001110;
    x_30 = 'b111011110;
    x_31 = 'b111100000;
    x_32 = 'b111011110;
    x_33 = 'b111100011;
    x_34 = 'b111101111;
    x_35 = 'b111101110;
    x_36 = 'b111101110;
    x_37 = 'b111110010;
    x_38 = 'b111001100;
    x_39 = 'b111110011;
    x_40 = 'b111000101;
    x_41 = 'b111100111;
    x_42 = 'b111000010;
    x_43 = 'b111111011;
    x_44 = 'b111011100;
    x_45 = 'b111110001;
    x_46 = 'b111101101;
    x_47 = 'b111101101;
    x_48 = 'b111111000;
    x_49 = 'b111111010;
    x_50 = 'b000000110;
    x_51 = 'b000010101;
    x_52 = 'b000010001;
    x_53 = 'b000010011;
    x_54 = 'b000001111;
    x_55 = 'b111111001;
    x_56 = 'b111111100;
    x_57 = 'b000010110;
    x_58 = 'b000011000;
    x_59 = 'b000010100;
    x_60 = 'b111111000;
    x_61 = 'b000000101;
    x_62 = 'b111110111;
    x_63 = 'b111110001;

    h_0 = 'b111010001;
    h_1 = 'b111100100;
    h_2 = 'b111100111;
    h_3 = 'b111110111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111010101;
    x_1 = 'b111101010;
    x_2 = 'b111101010;
    x_3 = 'b111111011;
    x_4 = 'b000000100;
    x_5 = 'b000001001;
    x_6 = 'b111111010;
    x_7 = 'b111101011;
    x_8 = 'b111110010;
    x_9 = 'b111110100;
    x_10 = 'b111111100;
    x_11 = 'b000001011;
    x_12 = 'b000010011;
    x_13 = 'b000001001;
    x_14 = 'b111101000;
    x_15 = 'b111101011;
    x_16 = 'b111110101;
    x_17 = 'b000000100;
    x_18 = 'b000010001;
    x_19 = 'b000010101;
    x_20 = 'b000010011;
    x_21 = 'b111010001;
    x_22 = 'b111010100;
    x_23 = 'b111011010;
    x_24 = 'b111001110;
    x_25 = 'b111001111;
    x_26 = 'b111100000;
    x_27 = 'b111100111;
    x_28 = 'b111011111;
    x_29 = 'b111010100;
    x_30 = 'b111101010;
    x_31 = 'b111101011;
    x_32 = 'b111100100;
    x_33 = 'b111101010;
    x_34 = 'b111110111;
    x_35 = 'b111110111;
    x_36 = 'b111110111;
    x_37 = 'b111110010;
    x_38 = 'b111011101;
    x_39 = 'b111111011;
    x_40 = 'b111101000;
    x_41 = 'b111110101;
    x_42 = 'b111000111;
    x_43 = 'b000000101;
    x_44 = 'b111100101;
    x_45 = 'b000000001;
    x_46 = 'b111110110;
    x_47 = 'b111110011;
    x_48 = 'b111111010;
    x_49 = 'b000000010;
    x_50 = 'b000001110;
    x_51 = 'b000011110;
    x_52 = 'b000011000;
    x_53 = 'b000011010;
    x_54 = 'b000010110;
    x_55 = 'b000000001;
    x_56 = 'b000000011;
    x_57 = 'b000011011;
    x_58 = 'b000011110;
    x_59 = 'b000011001;
    x_60 = 'b000000010;
    x_61 = 'b000010001;
    x_62 = 'b000000010;
    x_63 = 'b111111110;

    h_0 = 'b111010101;
    h_1 = 'b111101010;
    h_2 = 'b111101010;
    h_3 = 'b111111011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111100100;
    x_1 = 'b111110010;
    x_2 = 'b111110000;
    x_3 = 'b000000000;
    x_4 = 'b000000110;
    x_5 = 'b000000111;
    x_6 = 'b111111100;
    x_7 = 'b111101110;
    x_8 = 'b111110010;
    x_9 = 'b111110111;
    x_10 = 'b111111111;
    x_11 = 'b000001001;
    x_12 = 'b000001110;
    x_13 = 'b000000001;
    x_14 = 'b111100001;
    x_15 = 'b111101010;
    x_16 = 'b111111000;
    x_17 = 'b000000101;
    x_18 = 'b000001101;
    x_19 = 'b000001110;
    x_20 = 'b000001010;
    x_21 = 'b111011000;
    x_22 = 'b111011001;
    x_23 = 'b111011101;
    x_24 = 'b111010101;
    x_25 = 'b111010110;
    x_26 = 'b111100110;
    x_27 = 'b111100111;
    x_28 = 'b111011101;
    x_29 = 'b111011011;
    x_30 = 'b111110011;
    x_31 = 'b111101011;
    x_32 = 'b111101011;
    x_33 = 'b111101110;
    x_34 = 'b111110111;
    x_35 = 'b111111000;
    x_36 = 'b111110001;
    x_37 = 'b111110010;
    x_38 = 'b111100101;
    x_39 = 'b111110011;
    x_40 = 'b111011110;
    x_41 = 'b000001011;
    x_42 = 'b111000110;
    x_43 = 'b111101110;
    x_44 = 'b111100111;
    x_45 = 'b111101001;
    x_46 = 'b111111000;
    x_47 = 'b111110001;
    x_48 = 'b111111010;
    x_49 = 'b111111101;
    x_50 = 'b000000111;
    x_51 = 'b000001100;
    x_52 = 'b000000101;
    x_53 = 'b000000101;
    x_54 = 'b111111100;
    x_55 = 'b111111101;
    x_56 = 'b111111110;
    x_57 = 'b000001110;
    x_58 = 'b000001001;
    x_59 = 'b000000010;
    x_60 = 'b000000111;
    x_61 = 'b000010000;
    x_62 = 'b111111111;
    x_63 = 'b111111011;

    h_0 = 'b111100100;
    h_1 = 'b111110010;
    h_2 = 'b111110000;
    h_3 = 'b000000000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111100111;
    x_1 = 'b111111000;
    x_2 = 'b111110011;
    x_3 = 'b000000010;
    x_4 = 'b000000010;
    x_5 = 'b000000001;
    x_6 = 'b111111000;
    x_7 = 'b111110011;
    x_8 = 'b111110111;
    x_9 = 'b111111100;
    x_10 = 'b000000010;
    x_11 = 'b000001001;
    x_12 = 'b000001001;
    x_13 = 'b111111111;
    x_14 = 'b111101100;
    x_15 = 'b111110100;
    x_16 = 'b111111110;
    x_17 = 'b000001001;
    x_18 = 'b000000110;
    x_19 = 'b000000110;
    x_20 = 'b000000101;
    x_21 = 'b111011010;
    x_22 = 'b111011010;
    x_23 = 'b111100000;
    x_24 = 'b111011000;
    x_25 = 'b111011000;
    x_26 = 'b111101010;
    x_27 = 'b111101010;
    x_28 = 'b111100010;
    x_29 = 'b111011010;
    x_30 = 'b111110100;
    x_31 = 'b111101111;
    x_32 = 'b111101111;
    x_33 = 'b111110010;
    x_34 = 'b111111010;
    x_35 = 'b111111010;
    x_36 = 'b111110100;
    x_37 = 'b111111100;
    x_38 = 'b111011011;
    x_39 = 'b111111011;
    x_40 = 'b111011001;
    x_41 = 'b000011000;
    x_42 = 'b111001111;
    x_43 = 'b111100111;
    x_44 = 'b111101100;
    x_45 = 'b111110010;
    x_46 = 'b111111110;
    x_47 = 'b111111111;
    x_48 = 'b000001001;
    x_49 = 'b000001000;
    x_50 = 'b000001100;
    x_51 = 'b000001101;
    x_52 = 'b000000111;
    x_53 = 'b000000111;
    x_54 = 'b000000101;
    x_55 = 'b000001101;
    x_56 = 'b000001011;
    x_57 = 'b000010101;
    x_58 = 'b000001001;
    x_59 = 'b000000101;
    x_60 = 'b000001100;
    x_61 = 'b000001100;
    x_62 = 'b111111001;
    x_63 = 'b111111010;

    h_0 = 'b111100111;
    h_1 = 'b111111000;
    h_2 = 'b111110011;
    h_3 = 'b000000010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111100100;
    x_1 = 'b111111010;
    x_2 = 'b111110100;
    x_3 = 'b000000010;
    x_4 = 'b000000001;
    x_5 = 'b000000100;
    x_6 = 'b111111010;
    x_7 = 'b111111100;
    x_8 = 'b000000000;
    x_9 = 'b111111110;
    x_10 = 'b111111111;
    x_11 = 'b000001001;
    x_12 = 'b000000110;
    x_13 = 'b000000001;
    x_14 = 'b111110111;
    x_15 = 'b111111101;
    x_16 = 'b000000000;
    x_17 = 'b000000100;
    x_18 = 'b000000000;
    x_19 = 'b111111111;
    x_20 = 'b000000010;
    x_21 = 'b111011011;
    x_22 = 'b111011101;
    x_23 = 'b111100010;
    x_24 = 'b111010101;
    x_25 = 'b111010110;
    x_26 = 'b111101010;
    x_27 = 'b111101011;
    x_28 = 'b111100101;
    x_29 = 'b111010110;
    x_30 = 'b111101100;
    x_31 = 'b111101010;
    x_32 = 'b111101001;
    x_33 = 'b111101100;
    x_34 = 'b111110101;
    x_35 = 'b111110011;
    x_36 = 'b111110001;
    x_37 = 'b111110101;
    x_38 = 'b111011111;
    x_39 = 'b111101111;
    x_40 = 'b111100111;
    x_41 = 'b111101100;
    x_42 = 'b111010111;
    x_43 = 'b111011011;
    x_44 = 'b111101110;
    x_45 = 'b111100100;
    x_46 = 'b111111110;
    x_47 = 'b111111100;
    x_48 = 'b000000011;
    x_49 = 'b111111101;
    x_50 = 'b111111010;
    x_51 = 'b111111010;
    x_52 = 'b111110001;
    x_53 = 'b111110111;
    x_54 = 'b111110110;
    x_55 = 'b000000111;
    x_56 = 'b000000011;
    x_57 = 'b000000101;
    x_58 = 'b111110111;
    x_59 = 'b111111100;
    x_60 = 'b000001101;
    x_61 = 'b000000111;
    x_62 = 'b111110101;
    x_63 = 'b111111101;

    h_0 = 'b111100100;
    h_1 = 'b111111010;
    h_2 = 'b111110100;
    h_3 = 'b000000010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111011101;
    x_1 = 'b111101000;
    x_2 = 'b111100111;
    x_3 = 'b111110111;
    x_4 = 'b111110110;
    x_5 = 'b111110011;
    x_6 = 'b111101011;
    x_7 = 'b111101100;
    x_8 = 'b111110001;
    x_9 = 'b111101110;
    x_10 = 'b111101111;
    x_11 = 'b111111010;
    x_12 = 'b111110011;
    x_13 = 'b111101001;
    x_14 = 'b111101110;
    x_15 = 'b111110000;
    x_16 = 'b111110001;
    x_17 = 'b111110001;
    x_18 = 'b111101101;
    x_19 = 'b111101110;
    x_20 = 'b111110000;
    x_21 = 'b111011011;
    x_22 = 'b111011100;
    x_23 = 'b111100001;
    x_24 = 'b111010110;
    x_25 = 'b111010110;
    x_26 = 'b111101010;
    x_27 = 'b111101000;
    x_28 = 'b111100010;
    x_29 = 'b111011001;
    x_30 = 'b111101100;
    x_31 = 'b111100110;
    x_32 = 'b111101010;
    x_33 = 'b111101111;
    x_34 = 'b111110110;
    x_35 = 'b111110011;
    x_36 = 'b111101100;
    x_37 = 'b111110001;
    x_38 = 'b111101101;
    x_39 = 'b111101010;
    x_40 = 'b111110100;
    x_41 = 'b111100010;
    x_42 = 'b111101010;
    x_43 = 'b111100111;
    x_44 = 'b111110000;
    x_45 = 'b111101100;
    x_46 = 'b000000001;
    x_47 = 'b111111110;
    x_48 = 'b000000010;
    x_49 = 'b111111010;
    x_50 = 'b111110110;
    x_51 = 'b111110110;
    x_52 = 'b111110010;
    x_53 = 'b111111101;
    x_54 = 'b000000000;
    x_55 = 'b000001100;
    x_56 = 'b000001000;
    x_57 = 'b000000100;
    x_58 = 'b111111010;
    x_59 = 'b000000110;
    x_60 = 'b000001100;
    x_61 = 'b000000110;
    x_62 = 'b111110111;
    x_63 = 'b000000111;

    h_0 = 'b111011101;
    h_1 = 'b111101000;
    h_2 = 'b111100111;
    h_3 = 'b111110111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111110001;
    x_1 = 'b111111011;
    x_2 = 'b111111000;
    x_3 = 'b000000111;
    x_4 = 'b000000110;
    x_5 = 'b000000001;
    x_6 = 'b111110101;
    x_7 = 'b000001011;
    x_8 = 'b000000110;
    x_9 = 'b000000000;
    x_10 = 'b000000001;
    x_11 = 'b000001101;
    x_12 = 'b000000100;
    x_13 = 'b111111001;
    x_14 = 'b000000011;
    x_15 = 'b000000101;
    x_16 = 'b000000010;
    x_17 = 'b000000010;
    x_18 = 'b111111100;
    x_19 = 'b111111111;
    x_20 = 'b000000100;
    x_21 = 'b111100011;
    x_22 = 'b111100101;
    x_23 = 'b111100111;
    x_24 = 'b111100010;
    x_25 = 'b111100010;
    x_26 = 'b111110101;
    x_27 = 'b111110010;
    x_28 = 'b111100111;
    x_29 = 'b111101001;
    x_30 = 'b000000000;
    x_31 = 'b111110110;
    x_32 = 'b111110111;
    x_33 = 'b111111010;
    x_34 = 'b000000011;
    x_35 = 'b111111111;
    x_36 = 'b111110111;
    x_37 = 'b111111001;
    x_38 = 'b111111100;
    x_39 = 'b111101101;
    x_40 = 'b000000010;
    x_41 = 'b111110000;
    x_42 = 'b111101000;
    x_43 = 'b111111101;
    x_44 = 'b000000000;
    x_45 = 'b111110010;
    x_46 = 'b000001011;
    x_47 = 'b000001000;
    x_48 = 'b000001100;
    x_49 = 'b000000001;
    x_50 = 'b111111010;
    x_51 = 'b111111000;
    x_52 = 'b111110010;
    x_53 = 'b111111011;
    x_54 = 'b111111101;
    x_55 = 'b000001110;
    x_56 = 'b000001010;
    x_57 = 'b000000010;
    x_58 = 'b111110110;
    x_59 = 'b111111010;
    x_60 = 'b000001110;
    x_61 = 'b000001010;
    x_62 = 'b111110111;
    x_63 = 'b000010010;

    h_0 = 'b111110001;
    h_1 = 'b111111011;
    h_2 = 'b111111000;
    h_3 = 'b000000111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111110101;
    x_1 = 'b111111011;
    x_2 = 'b111110100;
    x_3 = 'b111111111;
    x_4 = 'b111111101;
    x_5 = 'b111111001;
    x_6 = 'b111101110;
    x_7 = 'b000000100;
    x_8 = 'b111111111;
    x_9 = 'b111111001;
    x_10 = 'b111110111;
    x_11 = 'b111111101;
    x_12 = 'b111110001;
    x_13 = 'b111101001;
    x_14 = 'b111110100;
    x_15 = 'b111111000;
    x_16 = 'b111110101;
    x_17 = 'b111110101;
    x_18 = 'b111101011;
    x_19 = 'b111101001;
    x_20 = 'b111101010;
    x_21 = 'b111011110;
    x_22 = 'b111011111;
    x_23 = 'b111100000;
    x_24 = 'b111011011;
    x_25 = 'b111011100;
    x_26 = 'b111101010;
    x_27 = 'b111101001;
    x_28 = 'b111100000;
    x_29 = 'b111011001;
    x_30 = 'b111111101;
    x_31 = 'b111101000;
    x_32 = 'b111101000;
    x_33 = 'b111101001;
    x_34 = 'b111110011;
    x_35 = 'b111110000;
    x_36 = 'b111101001;
    x_37 = 'b111101011;
    x_38 = 'b111100100;
    x_39 = 'b111011110;
    x_40 = 'b111100100;
    x_41 = 'b111101100;
    x_42 = 'b111001011;
    x_43 = 'b111011101;
    x_44 = 'b111101001;
    x_45 = 'b111001100;
    x_46 = 'b111110010;
    x_47 = 'b111101110;
    x_48 = 'b111110000;
    x_49 = 'b111100111;
    x_50 = 'b111100011;
    x_51 = 'b111100000;
    x_52 = 'b111011001;
    x_53 = 'b111011111;
    x_54 = 'b111011100;
    x_55 = 'b111111001;
    x_56 = 'b111110110;
    x_57 = 'b111101110;
    x_58 = 'b111100011;
    x_59 = 'b111100101;
    x_60 = 'b000000111;
    x_61 = 'b111111111;
    x_62 = 'b111100110;
    x_63 = 'b000000110;

    h_0 = 'b111110101;
    h_1 = 'b111111011;
    h_2 = 'b111110100;
    h_3 = 'b111111111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111101001;
    x_1 = 'b111110010;
    x_2 = 'b111101101;
    x_3 = 'b111110100;
    x_4 = 'b111110101;
    x_5 = 'b111110011;
    x_6 = 'b111101110;
    x_7 = 'b111110000;
    x_8 = 'b111110001;
    x_9 = 'b111101111;
    x_10 = 'b111101101;
    x_11 = 'b111110111;
    x_12 = 'b111101100;
    x_13 = 'b111101001;
    x_14 = 'b111100111;
    x_15 = 'b111101001;
    x_16 = 'b111101010;
    x_17 = 'b111101011;
    x_18 = 'b111100111;
    x_19 = 'b111100111;
    x_20 = 'b111101001;
    x_21 = 'b111011111;
    x_22 = 'b111100000;
    x_23 = 'b111100001;
    x_24 = 'b111011110;
    x_25 = 'b111011101;
    x_26 = 'b111101111;
    x_27 = 'b111101100;
    x_28 = 'b111100000;
    x_29 = 'b111100000;
    x_30 = 'b111111010;
    x_31 = 'b111101011;
    x_32 = 'b111110000;
    x_33 = 'b111110010;
    x_34 = 'b111111001;
    x_35 = 'b111110110;
    x_36 = 'b111101111;
    x_37 = 'b111110001;
    x_38 = 'b111101011;
    x_39 = 'b111110100;
    x_40 = 'b111110011;
    x_41 = 'b000001100;
    x_42 = 'b111010010;
    x_43 = 'b111010000;
    x_44 = 'b111101011;
    x_45 = 'b111011001;
    x_46 = 'b111110101;
    x_47 = 'b111101110;
    x_48 = 'b111110001;
    x_49 = 'b111101100;
    x_50 = 'b111101011;
    x_51 = 'b111110000;
    x_52 = 'b111101001;
    x_53 = 'b111101110;
    x_54 = 'b111101011;
    x_55 = 'b111111100;
    x_56 = 'b111111001;
    x_57 = 'b111111001;
    x_58 = 'b111110110;
    x_59 = 'b111110110;
    x_60 = 'b111111111;
    x_61 = 'b111110111;
    x_62 = 'b111011111;
    x_63 = 'b111111011;

    h_0 = 'b111101001;
    h_1 = 'b111110010;
    h_2 = 'b111101101;
    h_3 = 'b111110100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111101011;
    x_1 = 'b111110110;
    x_2 = 'b111110100;
    x_3 = 'b111111101;
    x_4 = 'b111111111;
    x_5 = 'b000000000;
    x_6 = 'b111110101;
    x_7 = 'b111111000;
    x_8 = 'b111110101;
    x_9 = 'b111110100;
    x_10 = 'b111110101;
    x_11 = 'b000000001;
    x_12 = 'b111111011;
    x_13 = 'b111111000;
    x_14 = 'b111101011;
    x_15 = 'b111101101;
    x_16 = 'b111110010;
    x_17 = 'b111110010;
    x_18 = 'b111110101;
    x_19 = 'b111111000;
    x_20 = 'b111111000;
    x_21 = 'b111100000;
    x_22 = 'b111011110;
    x_23 = 'b111100000;
    x_24 = 'b111011110;
    x_25 = 'b111011111;
    x_26 = 'b111101101;
    x_27 = 'b111101010;
    x_28 = 'b111011111;
    x_29 = 'b111100011;
    x_30 = 'b111110101;
    x_31 = 'b111101110;
    x_32 = 'b111101111;
    x_33 = 'b111110011;
    x_34 = 'b111111001;
    x_35 = 'b111110100;
    x_36 = 'b111101110;
    x_37 = 'b111110001;
    x_38 = 'b111101100;
    x_39 = 'b111110111;
    x_40 = 'b111011010;
    x_41 = 'b111111010;
    x_42 = 'b111001111;
    x_43 = 'b111110111;
    x_44 = 'b111101001;
    x_45 = 'b111101101;
    x_46 = 'b111110001;
    x_47 = 'b111101110;
    x_48 = 'b111110001;
    x_49 = 'b111110011;
    x_50 = 'b111110101;
    x_51 = 'b111111110;
    x_52 = 'b111111010;
    x_53 = 'b111111110;
    x_54 = 'b111111011;
    x_55 = 'b111111000;
    x_56 = 'b111110101;
    x_57 = 'b000000001;
    x_58 = 'b000000100;
    x_59 = 'b000000100;
    x_60 = 'b111111100;
    x_61 = 'b111111010;
    x_62 = 'b111101011;
    x_63 = 'b111111110;

    h_0 = 'b111101011;
    h_1 = 'b111110110;
    h_2 = 'b111110100;
    h_3 = 'b111111101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000001110;
    x_1 = 'b000001110;
    x_2 = 'b000000110;
    x_3 = 'b000001100;
    x_4 = 'b000010000;
    x_5 = 'b000000111;
    x_6 = 'b000000111;
    x_7 = 'b000000011;
    x_8 = 'b000001010;
    x_9 = 'b000001100;
    x_10 = 'b000010001;
    x_11 = 'b000000010;
    x_12 = 'b000001011;
    x_13 = 'b000010000;
    x_14 = 'b000001011;
    x_15 = 'b000001100;
    x_16 = 'b000001101;
    x_17 = 'b000001011;
    x_18 = 'b000001011;
    x_19 = 'b000010000;
    x_20 = 'b000001000;
    x_21 = 'b000000100;
    x_22 = 'b000000110;
    x_23 = 'b111111100;
    x_24 = 'b111111011;
    x_25 = 'b111111100;
    x_26 = 'b111111100;
    x_27 = 'b111111101;
    x_28 = 'b000000100;
    x_29 = 'b000000110;
    x_30 = 'b111111100;
    x_31 = 'b111110110;
    x_32 = 'b111111101;
    x_33 = 'b111111011;
    x_34 = 'b111111000;
    x_35 = 'b111111011;
    x_36 = 'b111111011;
    x_37 = 'b000001000;
    x_38 = 'b111111100;
    x_39 = 'b000001100;
    x_40 = 'b111111111;
    x_41 = 'b111110000;
    x_42 = 'b111111011;
    x_43 = 'b000011110;
    x_44 = 'b111110001;
    x_45 = 'b000010101;
    x_46 = 'b000001000;
    x_47 = 'b000000111;
    x_48 = 'b000001001;
    x_49 = 'b000001000;
    x_50 = 'b000001101;
    x_51 = 'b000001111;
    x_52 = 'b000001101;
    x_53 = 'b000001011;
    x_54 = 'b000000111;
    x_55 = 'b000001010;
    x_56 = 'b000000111;
    x_57 = 'b000010010;
    x_58 = 'b000010101;
    x_59 = 'b000010111;
    x_60 = 'b000010111;
    x_61 = 'b000100101;
    x_62 = 'b000010010;
    x_63 = 'b000001111;

    h_0 = 'b000001110;
    h_1 = 'b000001110;
    h_2 = 'b000000110;
    h_3 = 'b000001100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000000101;
    x_1 = 'b000000110;
    x_2 = 'b000000001;
    x_3 = 'b000001010;
    x_4 = 'b000001101;
    x_5 = 'b000000000;
    x_6 = 'b111111110;
    x_7 = 'b111111011;
    x_8 = 'b000000011;
    x_9 = 'b000001001;
    x_10 = 'b000001101;
    x_11 = 'b000000011;
    x_12 = 'b000000110;
    x_13 = 'b000000111;
    x_14 = 'b000000110;
    x_15 = 'b000000100;
    x_16 = 'b000000110;
    x_17 = 'b000000110;
    x_18 = 'b000001000;
    x_19 = 'b000001011;
    x_20 = 'b000000010;
    x_21 = 'b000000111;
    x_22 = 'b000001001;
    x_23 = 'b000000000;
    x_24 = 'b111111100;
    x_25 = 'b111111101;
    x_26 = 'b000000000;
    x_27 = 'b000000001;
    x_28 = 'b000000110;
    x_29 = 'b000000011;
    x_30 = 'b111111100;
    x_31 = 'b111111000;
    x_32 = 'b000000001;
    x_33 = 'b000000001;
    x_34 = 'b111111101;
    x_35 = 'b111111101;
    x_36 = 'b111111000;
    x_37 = 'b000000110;
    x_38 = 'b111111001;
    x_39 = 'b000000000;
    x_40 = 'b000000000;
    x_41 = 'b111011010;
    x_42 = 'b111101101;
    x_43 = 'b000010000;
    x_44 = 'b111101100;
    x_45 = 'b000100001;
    x_46 = 'b000000011;
    x_47 = 'b000000011;
    x_48 = 'b000000111;
    x_49 = 'b000001000;
    x_50 = 'b000001011;
    x_51 = 'b000001111;
    x_52 = 'b000001100;
    x_53 = 'b000001100;
    x_54 = 'b000001101;
    x_55 = 'b000001001;
    x_56 = 'b000000110;
    x_57 = 'b000010001;
    x_58 = 'b000010010;
    x_59 = 'b000011000;
    x_60 = 'b000010111;
    x_61 = 'b000100000;
    x_62 = 'b000001010;
    x_63 = 'b000010010;

    h_0 = 'b000000101;
    h_1 = 'b000000110;
    h_2 = 'b000000001;
    h_3 = 'b000001010;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111111011;
    x_1 = 'b000000000;
    x_2 = 'b000000000;
    x_3 = 'b000001100;
    x_4 = 'b000001110;
    x_5 = 'b000000000;
    x_6 = 'b111111010;
    x_7 = 'b111101111;
    x_8 = 'b111111010;
    x_9 = 'b000000101;
    x_10 = 'b000001111;
    x_11 = 'b000000000;
    x_12 = 'b000000011;
    x_13 = 'b000000110;
    x_14 = 'b111110111;
    x_15 = 'b111111110;
    x_16 = 'b000000010;
    x_17 = 'b000000100;
    x_18 = 'b000000100;
    x_19 = 'b000000101;
    x_20 = 'b111111111;
    x_21 = 'b111111101;
    x_22 = 'b111111110;
    x_23 = 'b111111000;
    x_24 = 'b111101101;
    x_25 = 'b111101110;
    x_26 = 'b111110100;
    x_27 = 'b111110101;
    x_28 = 'b111111110;
    x_29 = 'b111110010;
    x_30 = 'b111101001;
    x_31 = 'b111101110;
    x_32 = 'b111110011;
    x_33 = 'b111110101;
    x_34 = 'b111110000;
    x_35 = 'b111101110;
    x_36 = 'b111101000;
    x_37 = 'b111111000;
    x_38 = 'b111100111;
    x_39 = 'b111111010;
    x_40 = 'b111100101;
    x_41 = 'b111100100;
    x_42 = 'b111100010;
    x_43 = 'b111111110;
    x_44 = 'b111100000;
    x_45 = 'b000011111;
    x_46 = 'b111111000;
    x_47 = 'b111111100;
    x_48 = 'b000000000;
    x_49 = 'b000000010;
    x_50 = 'b000000011;
    x_51 = 'b000000101;
    x_52 = 'b000000010;
    x_53 = 'b000000101;
    x_54 = 'b000001101;
    x_55 = 'b000001010;
    x_56 = 'b000000011;
    x_57 = 'b000001001;
    x_58 = 'b000001011;
    x_59 = 'b000011000;
    x_60 = 'b000010101;
    x_61 = 'b000011100;
    x_62 = 'b000000010;
    x_63 = 'b000010001;

    h_0 = 'b111111011;
    h_1 = 'b000000000;
    h_2 = 'b000000000;
    h_3 = 'b000001100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111101101;
    x_1 = 'b111110011;
    x_2 = 'b111110010;
    x_3 = 'b111111100;
    x_4 = 'b111111110;
    x_5 = 'b111110000;
    x_6 = 'b111101001;
    x_7 = 'b111100001;
    x_8 = 'b111110000;
    x_9 = 'b111111010;
    x_10 = 'b000000100;
    x_11 = 'b111101110;
    x_12 = 'b111110101;
    x_13 = 'b111111110;
    x_14 = 'b111110111;
    x_15 = 'b111111101;
    x_16 = 'b111111011;
    x_17 = 'b111111010;
    x_18 = 'b111110110;
    x_19 = 'b111111000;
    x_20 = 'b111110011;
    x_21 = 'b111111010;
    x_22 = 'b111111000;
    x_23 = 'b111110001;
    x_24 = 'b111101100;
    x_25 = 'b111101100;
    x_26 = 'b111101111;
    x_27 = 'b111101101;
    x_28 = 'b111110101;
    x_29 = 'b111110100;
    x_30 = 'b111101011;
    x_31 = 'b111100101;
    x_32 = 'b111110000;
    x_33 = 'b111101110;
    x_34 = 'b111101001;
    x_35 = 'b111101011;
    x_36 = 'b111100010;
    x_37 = 'b111110010;
    x_38 = 'b111110000;
    x_39 = 'b000000011;
    x_40 = 'b111111011;
    x_41 = 'b111111101;
    x_42 = 'b111110010;
    x_43 = 'b111101100;
    x_44 = 'b111101010;
    x_45 = 'b000001110;
    x_46 = 'b000000010;
    x_47 = 'b000000001;
    x_48 = 'b111111100;
    x_49 = 'b111111111;
    x_50 = 'b111111001;
    x_51 = 'b111111000;
    x_52 = 'b111110100;
    x_53 = 'b111110111;
    x_54 = 'b000000111;
    x_55 = 'b000001110;
    x_56 = 'b000000010;
    x_57 = 'b111111111;
    x_58 = 'b000000011;
    x_59 = 'b000011000;
    x_60 = 'b000010101;
    x_61 = 'b000011010;
    x_62 = 'b000000000;
    x_63 = 'b000010001;

    h_0 = 'b111101101;
    h_1 = 'b111110011;
    h_2 = 'b111110010;
    h_3 = 'b111111100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111110101;
    x_1 = 'b111111010;
    x_2 = 'b111110000;
    x_3 = 'b111110110;
    x_4 = 'b111110110;
    x_5 = 'b111101011;
    x_6 = 'b111101011;
    x_7 = 'b111101100;
    x_8 = 'b111110101;
    x_9 = 'b111110111;
    x_10 = 'b111111100;
    x_11 = 'b111101000;
    x_12 = 'b111101011;
    x_13 = 'b111111001;
    x_14 = 'b111111011;
    x_15 = 'b111111101;
    x_16 = 'b111110111;
    x_17 = 'b111110001;
    x_18 = 'b111101001;
    x_19 = 'b111101010;
    x_20 = 'b111100101;
    x_21 = 'b111110110;
    x_22 = 'b111110011;
    x_23 = 'b111101101;
    x_24 = 'b111101000;
    x_25 = 'b111101000;
    x_26 = 'b111101000;
    x_27 = 'b111101001;
    x_28 = 'b111110011;
    x_29 = 'b111101011;
    x_30 = 'b111100110;
    x_31 = 'b111100100;
    x_32 = 'b111101101;
    x_33 = 'b111101000;
    x_34 = 'b111100011;
    x_35 = 'b111100101;
    x_36 = 'b111100000;
    x_37 = 'b111101110;
    x_38 = 'b111101010;
    x_39 = 'b111110111;
    x_40 = 'b111101101;
    x_41 = 'b111100100;
    x_42 = 'b111100111;
    x_43 = 'b000010000;
    x_44 = 'b111101011;
    x_45 = 'b000001001;
    x_46 = 'b000000010;
    x_47 = 'b000000000;
    x_48 = 'b111111000;
    x_49 = 'b111111011;
    x_50 = 'b111110001;
    x_51 = 'b111110000;
    x_52 = 'b111101100;
    x_53 = 'b111110100;
    x_54 = 'b000000101;
    x_55 = 'b000000111;
    x_56 = 'b111111101;
    x_57 = 'b111110110;
    x_58 = 'b111111110;
    x_59 = 'b000011010;
    x_60 = 'b000010011;
    x_61 = 'b000010111;
    x_62 = 'b000000100;
    x_63 = 'b000010001;

    h_0 = 'b111110101;
    h_1 = 'b111111010;
    h_2 = 'b111110000;
    h_3 = 'b111110110;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111110101;
    x_1 = 'b111111010;
    x_2 = 'b111110011;
    x_3 = 'b111110101;
    x_4 = 'b111111010;
    x_5 = 'b111110000;
    x_6 = 'b111101101;
    x_7 = 'b111110011;
    x_8 = 'b111111010;
    x_9 = 'b111111100;
    x_10 = 'b111111110;
    x_11 = 'b111101101;
    x_12 = 'b111110000;
    x_13 = 'b111111001;
    x_14 = 'b000000010;
    x_15 = 'b000000100;
    x_16 = 'b111111011;
    x_17 = 'b111110100;
    x_18 = 'b111101100;
    x_19 = 'b111101101;
    x_20 = 'b111101000;
    x_21 = 'b111111100;
    x_22 = 'b111110110;
    x_23 = 'b111101110;
    x_24 = 'b111101110;
    x_25 = 'b111101110;
    x_26 = 'b111101111;
    x_27 = 'b111101110;
    x_28 = 'b111110011;
    x_29 = 'b111110110;
    x_30 = 'b111101111;
    x_31 = 'b111101110;
    x_32 = 'b111110110;
    x_33 = 'b111110010;
    x_34 = 'b111101101;
    x_35 = 'b111110000;
    x_36 = 'b111101011;
    x_37 = 'b111110100;
    x_38 = 'b111110101;
    x_39 = 'b000000000;
    x_40 = 'b111111110;
    x_41 = 'b111011111;
    x_42 = 'b111111110;
    x_43 = 'b000010000;
    x_44 = 'b111111010;
    x_45 = 'b000010010;
    x_46 = 'b000001001;
    x_47 = 'b000000101;
    x_48 = 'b111111101;
    x_49 = 'b111111101;
    x_50 = 'b111110010;
    x_51 = 'b111110001;
    x_52 = 'b111101110;
    x_53 = 'b111110111;
    x_54 = 'b000000010;
    x_55 = 'b000000110;
    x_56 = 'b111111100;
    x_57 = 'b111110011;
    x_58 = 'b111111100;
    x_59 = 'b000010011;
    x_60 = 'b000010000;
    x_61 = 'b000010010;
    x_62 = 'b000000101;
    x_63 = 'b000001101;

    h_0 = 'b111110101;
    h_1 = 'b111111010;
    h_2 = 'b111110011;
    h_3 = 'b111110101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000000001;
    x_1 = 'b000000011;
    x_2 = 'b111111010;
    x_3 = 'b111111011;
    x_4 = 'b000000010;
    x_5 = 'b111111110;
    x_6 = 'b111111111;
    x_7 = 'b111111011;
    x_8 = 'b000000000;
    x_9 = 'b000000010;
    x_10 = 'b000000100;
    x_11 = 'b111110100;
    x_12 = 'b111111111;
    x_13 = 'b000001001;
    x_14 = 'b000001001;
    x_15 = 'b000000111;
    x_16 = 'b000000000;
    x_17 = 'b111111001;
    x_18 = 'b111110110;
    x_19 = 'b111111001;
    x_20 = 'b111110101;
    x_21 = 'b000000111;
    x_22 = 'b000000011;
    x_23 = 'b111111010;
    x_24 = 'b111111010;
    x_25 = 'b111111001;
    x_26 = 'b111110110;
    x_27 = 'b111111011;
    x_28 = 'b111111111;
    x_29 = 'b000000101;
    x_30 = 'b111111011;
    x_31 = 'b111110011;
    x_32 = 'b111111010;
    x_33 = 'b111110101;
    x_34 = 'b111110011;
    x_35 = 'b111111000;
    x_36 = 'b111111000;
    x_37 = 'b111111111;
    x_38 = 'b000000001;
    x_39 = 'b000010110;
    x_40 = 'b000010000;
    x_41 = 'b000000101;
    x_42 = 'b000000111;
    x_43 = 'b000010001;
    x_44 = 'b111111110;
    x_45 = 'b000011001;
    x_46 = 'b000001101;
    x_47 = 'b000001011;
    x_48 = 'b000000010;
    x_49 = 'b111111111;
    x_50 = 'b111110111;
    x_51 = 'b111110010;
    x_52 = 'b111110010;
    x_53 = 'b111111010;
    x_54 = 'b111111111;
    x_55 = 'b000001001;
    x_56 = 'b000000010;
    x_57 = 'b111110101;
    x_58 = 'b111110110;
    x_59 = 'b000000110;
    x_60 = 'b000001001;
    x_61 = 'b000000101;
    x_62 = 'b111111001;
    x_63 = 'b111111111;

    h_0 = 'b000000001;
    h_1 = 'b000000011;
    h_2 = 'b111111010;
    h_3 = 'b111111011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000001000;
    x_1 = 'b000001000;
    x_2 = 'b111111111;
    x_3 = 'b000000000;
    x_4 = 'b000000100;
    x_5 = 'b000000000;
    x_6 = 'b000000000;
    x_7 = 'b000000100;
    x_8 = 'b000000111;
    x_9 = 'b000001010;
    x_10 = 'b000010001;
    x_11 = 'b111111011;
    x_12 = 'b000000111;
    x_13 = 'b000001110;
    x_14 = 'b000010101;
    x_15 = 'b000010000;
    x_16 = 'b000001000;
    x_17 = 'b000000010;
    x_18 = 'b111111110;
    x_19 = 'b000000010;
    x_20 = 'b111111110;
    x_21 = 'b111111111;
    x_22 = 'b000000000;
    x_23 = 'b111111000;
    x_24 = 'b111110110;
    x_25 = 'b111110101;
    x_26 = 'b111110001;
    x_27 = 'b111111000;
    x_28 = 'b000000000;
    x_29 = 'b000000000;
    x_30 = 'b111110101;
    x_31 = 'b111110001;
    x_32 = 'b111111000;
    x_33 = 'b111110010;
    x_34 = 'b111101101;
    x_35 = 'b111110001;
    x_36 = 'b111110000;
    x_37 = 'b111110010;
    x_38 = 'b000000000;
    x_39 = 'b000001011;
    x_40 = 'b000011000;
    x_41 = 'b111101110;
    x_42 = 'b111110001;
    x_43 = 'b000011110;
    x_44 = 'b000000101;
    x_45 = 'b000011011;
    x_46 = 'b000011101;
    x_47 = 'b000011010;
    x_48 = 'b000001101;
    x_49 = 'b000001101;
    x_50 = 'b000000010;
    x_51 = 'b111110101;
    x_52 = 'b111110100;
    x_53 = 'b111111010;
    x_54 = 'b111111011;
    x_55 = 'b000010010;
    x_56 = 'b000010000;
    x_57 = 'b111111010;
    x_58 = 'b111101101;
    x_59 = 'b111111000;
    x_60 = 'b000001001;
    x_61 = 'b111111001;
    x_62 = 'b111100101;
    x_63 = 'b111110110;

    h_0 = 'b000001000;
    h_1 = 'b000001000;
    h_2 = 'b111111111;
    h_3 = 'b000000000;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000001011;
    x_1 = 'b000001001;
    x_2 = 'b000000001;
    x_3 = 'b000000110;
    x_4 = 'b000001001;
    x_5 = 'b000000000;
    x_6 = 'b111110101;
    x_7 = 'b000001000;
    x_8 = 'b000000111;
    x_9 = 'b000001100;
    x_10 = 'b000010101;
    x_11 = 'b000000000;
    x_12 = 'b000001011;
    x_13 = 'b000001111;
    x_14 = 'b000010110;
    x_15 = 'b000001111;
    x_16 = 'b000001100;
    x_17 = 'b000001001;
    x_18 = 'b000000010;
    x_19 = 'b000000011;
    x_20 = 'b111111111;
    x_21 = 'b111111011;
    x_22 = 'b111111101;
    x_23 = 'b111110101;
    x_24 = 'b111110101;
    x_25 = 'b111110100;
    x_26 = 'b111110011;
    x_27 = 'b111110100;
    x_28 = 'b111111010;
    x_29 = 'b000000000;
    x_30 = 'b111110011;
    x_31 = 'b111110010;
    x_32 = 'b111111110;
    x_33 = 'b111111000;
    x_34 = 'b111110001;
    x_35 = 'b111110111;
    x_36 = 'b111101110;
    x_37 = 'b111101100;
    x_38 = 'b000000100;
    x_39 = 'b000000001;
    x_40 = 'b000001010;
    x_41 = 'b111011010;
    x_42 = 'b111110011;
    x_43 = 'b000010000;
    x_44 = 'b111110111;
    x_45 = 'b000001101;
    x_46 = 'b000001010;
    x_47 = 'b000001110;
    x_48 = 'b000000110;
    x_49 = 'b000001001;
    x_50 = 'b111111110;
    x_51 = 'b111101011;
    x_52 = 'b111101010;
    x_53 = 'b111100111;
    x_54 = 'b111100101;
    x_55 = 'b000000011;
    x_56 = 'b000000110;
    x_57 = 'b111101110;
    x_58 = 'b111010100;
    x_59 = 'b111010011;
    x_60 = 'b000000000;
    x_61 = 'b111100111;
    x_62 = 'b111000110;
    x_63 = 'b111100011;

    h_0 = 'b000001011;
    h_1 = 'b000001001;
    h_2 = 'b000000001;
    h_3 = 'b000000110;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000001110;
    x_1 = 'b000001110;
    x_2 = 'b000001001;
    x_3 = 'b000001111;
    x_4 = 'b000010101;
    x_5 = 'b000001011;
    x_6 = 'b000000000;
    x_7 = 'b000000000;
    x_8 = 'b000000101;
    x_9 = 'b000001111;
    x_10 = 'b000011100;
    x_11 = 'b000001101;
    x_12 = 'b000001110;
    x_13 = 'b000001110;
    x_14 = 'b000000100;
    x_15 = 'b000000111;
    x_16 = 'b000001010;
    x_17 = 'b000001010;
    x_18 = 'b000000011;
    x_19 = 'b111111111;
    x_20 = 'b111111000;
    x_21 = 'b000000011;
    x_22 = 'b000000101;
    x_23 = 'b111111110;
    x_24 = 'b111111001;
    x_25 = 'b111111000;
    x_26 = 'b000000000;
    x_27 = 'b000000010;
    x_28 = 'b000000110;
    x_29 = 'b111111011;
    x_30 = 'b111111010;
    x_31 = 'b111111111;
    x_32 = 'b000001000;
    x_33 = 'b000001000;
    x_34 = 'b000000000;
    x_35 = 'b000000011;
    x_36 = 'b000000010;
    x_37 = 'b000000100;
    x_38 = 'b111111110;
    x_39 = 'b000011000;
    x_40 = 'b111111110;
    x_41 = 'b111100011;
    x_42 = 'b111100111;
    x_43 = 'b000000001;
    x_44 = 'b111100111;
    x_45 = 'b000000101;
    x_46 = 'b111110011;
    x_47 = 'b111111010;
    x_48 = 'b111110111;
    x_49 = 'b111111111;
    x_50 = 'b111111001;
    x_51 = 'b111100001;
    x_52 = 'b111011111;
    x_53 = 'b111010110;
    x_54 = 'b111010000;
    x_55 = 'b111101111;
    x_56 = 'b111110010;
    x_57 = 'b111100001;
    x_58 = 'b111000011;
    x_59 = 'b110110100;
    x_60 = 'b111101011;
    x_61 = 'b111001100;
    x_62 = 'b110100011;
    x_63 = 'b111000110;

    h_0 = 'b000001110;
    h_1 = 'b000001110;
    h_2 = 'b000001001;
    h_3 = 'b000001111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000001001;
    x_1 = 'b000010010;
    x_2 = 'b000010101;
    x_3 = 'b000011101;
    x_4 = 'b000011101;
    x_5 = 'b000010001;
    x_6 = 'b000001011;
    x_7 = 'b000000000;
    x_8 = 'b000001000;
    x_9 = 'b000011000;
    x_10 = 'b000100110;
    x_11 = 'b000001111;
    x_12 = 'b000001100;
    x_13 = 'b000001010;
    x_14 = 'b111111011;
    x_15 = 'b000001000;
    x_16 = 'b000001100;
    x_17 = 'b000001100;
    x_18 = 'b000000100;
    x_19 = 'b111111101;
    x_20 = 'b111110001;
    x_21 = 'b000000111;
    x_22 = 'b000001000;
    x_23 = 'b000000010;
    x_24 = 'b111111011;
    x_25 = 'b111111011;
    x_26 = 'b000000111;
    x_27 = 'b000000110;
    x_28 = 'b000001010;
    x_29 = 'b111111011;
    x_30 = 'b111111111;
    x_31 = 'b000000101;
    x_32 = 'b000010000;
    x_33 = 'b000010001;
    x_34 = 'b000001010;
    x_35 = 'b000001010;
    x_36 = 'b000000101;
    x_37 = 'b000000001;
    x_38 = 'b111111010;
    x_39 = 'b000011001;
    x_40 = 'b111110110;
    x_41 = 'b111111110;
    x_42 = 'b111110111;
    x_43 = 'b000011110;
    x_44 = 'b111110101;
    x_45 = 'b000000011;
    x_46 = 'b111110111;
    x_47 = 'b111111100;
    x_48 = 'b111111010;
    x_49 = 'b000000111;
    x_50 = 'b000000100;
    x_51 = 'b111101110;
    x_52 = 'b111101011;
    x_53 = 'b111100011;
    x_54 = 'b111011010;
    x_55 = 'b111110010;
    x_56 = 'b111110110;
    x_57 = 'b111101111;
    x_58 = 'b111010011;
    x_59 = 'b111000111;
    x_60 = 'b111011110;
    x_61 = 'b111000000;
    x_62 = 'b110010111;
    x_63 = 'b110111110;

    h_0 = 'b000001001;
    h_1 = 'b000010010;
    h_2 = 'b000010101;
    h_3 = 'b000011101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000001110;
    x_1 = 'b000011011;
    x_2 = 'b000011111;
    x_3 = 'b000100101;
    x_4 = 'b000100001;
    x_5 = 'b000010100;
    x_6 = 'b000001011;
    x_7 = 'b000000001;
    x_8 = 'b000010101;
    x_9 = 'b000100110;
    x_10 = 'b000110010;
    x_11 = 'b000010011;
    x_12 = 'b000010001;
    x_13 = 'b000010110;
    x_14 = 'b000000111;
    x_15 = 'b000010110;
    x_16 = 'b000011101;
    x_17 = 'b000011100;
    x_18 = 'b000010000;
    x_19 = 'b000000111;
    x_20 = 'b111111011;
    x_21 = 'b000001011;
    x_22 = 'b000001001;
    x_23 = 'b111111110;
    x_24 = 'b000000101;
    x_25 = 'b000000100;
    x_26 = 'b000000110;
    x_27 = 'b000000011;
    x_28 = 'b000000110;
    x_29 = 'b000010010;
    x_30 = 'b111111101;
    x_31 = 'b000000100;
    x_32 = 'b000010001;
    x_33 = 'b000001111;
    x_34 = 'b000001011;
    x_35 = 'b000001011;
    x_36 = 'b000000010;
    x_37 = 'b111110101;
    x_38 = 'b000001110;
    x_39 = 'b000011001;
    x_40 = 'b000010101;
    x_41 = 'b111111100;
    x_42 = 'b000010001;
    x_43 = 'b000001000;
    x_44 = 'b000000110;
    x_45 = 'b000000011;
    x_46 = 'b000000101;
    x_47 = 'b000001010;
    x_48 = 'b000000101;
    x_49 = 'b000010100;
    x_50 = 'b000010101;
    x_51 = 'b000000000;
    x_52 = 'b111111011;
    x_53 = 'b111110000;
    x_54 = 'b111100011;
    x_55 = 'b111111001;
    x_56 = 'b000000000;
    x_57 = 'b000000001;
    x_58 = 'b111101001;
    x_59 = 'b111011100;
    x_60 = 'b111100001;
    x_61 = 'b111001101;
    x_62 = 'b110100111;
    x_63 = 'b110111111;

    h_0 = 'b000001110;
    h_1 = 'b000011011;
    h_2 = 'b000011111;
    h_3 = 'b000100101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000011010;
    x_1 = 'b000100110;
    x_2 = 'b000100111;
    x_3 = 'b000101011;
    x_4 = 'b000100111;
    x_5 = 'b000011011;
    x_6 = 'b000010010;
    x_7 = 'b000010110;
    x_8 = 'b000100111;
    x_9 = 'b000110101;
    x_10 = 'b001000010;
    x_11 = 'b000100110;
    x_12 = 'b000011101;
    x_13 = 'b000011100;
    x_14 = 'b000100000;
    x_15 = 'b000101101;
    x_16 = 'b000110011;
    x_17 = 'b000110001;
    x_18 = 'b000100111;
    x_19 = 'b000011110;
    x_20 = 'b000001100;
    x_21 = 'b000010011;
    x_22 = 'b000010000;
    x_23 = 'b000000110;
    x_24 = 'b000001100;
    x_25 = 'b000001011;
    x_26 = 'b000001111;
    x_27 = 'b000001111;
    x_28 = 'b000001111;
    x_29 = 'b000011001;
    x_30 = 'b000000101;
    x_31 = 'b000010001;
    x_32 = 'b000011100;
    x_33 = 'b000011010;
    x_34 = 'b000010101;
    x_35 = 'b000010111;
    x_36 = 'b000010001;
    x_37 = 'b000000001;
    x_38 = 'b000011101;
    x_39 = 'b000100001;
    x_40 = 'b000101110;
    x_41 = 'b000000011;
    x_42 = 'b000010010;
    x_43 = 'b111111001;
    x_44 = 'b000011111;
    x_45 = 'b000011001;
    x_46 = 'b000011100;
    x_47 = 'b000100011;
    x_48 = 'b000011101;
    x_49 = 'b000101010;
    x_50 = 'b000101100;
    x_51 = 'b000100000;
    x_52 = 'b000011011;
    x_53 = 'b000001110;
    x_54 = 'b000000011;
    x_55 = 'b000001110;
    x_56 = 'b000010101;
    x_57 = 'b000011001;
    x_58 = 'b000001010;
    x_59 = 'b111111101;
    x_60 = 'b111110111;
    x_61 = 'b111101011;
    x_62 = 'b111001110;
    x_63 = 'b111001111;

    h_0 = 'b000011010;
    h_1 = 'b000100110;
    h_2 = 'b000100111;
    h_3 = 'b000101011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000100100;
    x_1 = 'b000101111;
    x_2 = 'b000101111;
    x_3 = 'b000110001;
    x_4 = 'b000101110;
    x_5 = 'b000100010;
    x_6 = 'b000011000;
    x_7 = 'b000100001;
    x_8 = 'b000110000;
    x_9 = 'b000111001;
    x_10 = 'b001000001;
    x_11 = 'b000101110;
    x_12 = 'b000101000;
    x_13 = 'b000100111;
    x_14 = 'b000101000;
    x_15 = 'b000110001;
    x_16 = 'b000110101;
    x_17 = 'b000110000;
    x_18 = 'b000101101;
    x_19 = 'b000101011;
    x_20 = 'b000011010;
    x_21 = 'b000001101;
    x_22 = 'b000001010;
    x_23 = 'b111111101;
    x_24 = 'b000000010;
    x_25 = 'b000000010;
    x_26 = 'b000000111;
    x_27 = 'b000000100;
    x_28 = 'b111111110;
    x_29 = 'b000001100;
    x_30 = 'b000000000;
    x_31 = 'b000000111;
    x_32 = 'b000010010;
    x_33 = 'b000001111;
    x_34 = 'b000001000;
    x_35 = 'b000001001;
    x_36 = 'b111111101;
    x_37 = 'b111110100;
    x_38 = 'b000010010;
    x_39 = 'b000010101;
    x_40 = 'b000011101;
    x_41 = 'b111111000;
    x_42 = 'b000000001;
    x_43 = 'b111011111;
    x_44 = 'b000001110;
    x_45 = 'b000010010;
    x_46 = 'b000010110;
    x_47 = 'b000011100;
    x_48 = 'b000010100;
    x_49 = 'b000100000;
    x_50 = 'b000011111;
    x_51 = 'b000011110;
    x_52 = 'b000011010;
    x_53 = 'b000010001;
    x_54 = 'b000000100;
    x_55 = 'b000001100;
    x_56 = 'b000001111;
    x_57 = 'b000011000;
    x_58 = 'b000010010;
    x_59 = 'b000001010;
    x_60 = 'b000001010;
    x_61 = 'b000000101;
    x_62 = 'b111110010;
    x_63 = 'b111100011;

    h_0 = 'b000100100;
    h_1 = 'b000101111;
    h_2 = 'b000101111;
    h_3 = 'b000110001;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000010010;
    x_1 = 'b000011010;
    x_2 = 'b000010110;
    x_3 = 'b000010101;
    x_4 = 'b000010001;
    x_5 = 'b000000011;
    x_6 = 'b111110100;
    x_7 = 'b000001111;
    x_8 = 'b000011101;
    x_9 = 'b000100000;
    x_10 = 'b000100111;
    x_11 = 'b000010110;
    x_12 = 'b000010100;
    x_13 = 'b000001101;
    x_14 = 'b000011000;
    x_15 = 'b000100001;
    x_16 = 'b000100011;
    x_17 = 'b000011110;
    x_18 = 'b000011111;
    x_19 = 'b000011111;
    x_20 = 'b000010001;
    x_21 = 'b111111011;
    x_22 = 'b111111010;
    x_23 = 'b111110001;
    x_24 = 'b111110010;
    x_25 = 'b111110010;
    x_26 = 'b111110010;
    x_27 = 'b111110001;
    x_28 = 'b111111100;
    x_29 = 'b111111100;
    x_30 = 'b111110010;
    x_31 = 'b111101111;
    x_32 = 'b111111111;
    x_33 = 'b111110111;
    x_34 = 'b111101111;
    x_35 = 'b111110011;
    x_36 = 'b111100111;
    x_37 = 'b111101010;
    x_38 = 'b000000000;
    x_39 = 'b000000000;
    x_40 = 'b000000111;
    x_41 = 'b111010111;
    x_42 = 'b000000001;
    x_43 = 'b000010110;
    x_44 = 'b000000111;
    x_45 = 'b000011010;
    x_46 = 'b000011011;
    x_47 = 'b000011100;
    x_48 = 'b000011000;
    x_49 = 'b000100101;
    x_50 = 'b000100011;
    x_51 = 'b000101000;
    x_52 = 'b000100101;
    x_53 = 'b000100000;
    x_54 = 'b000011001;
    x_55 = 'b000011001;
    x_56 = 'b000011101;
    x_57 = 'b000101000;
    x_58 = 'b000100111;
    x_59 = 'b000100101;
    x_60 = 'b000011011;
    x_61 = 'b000011110;
    x_62 = 'b000001101;
    x_63 = 'b111111110;

    h_0 = 'b000010010;
    h_1 = 'b000011010;
    h_2 = 'b000010110;
    h_3 = 'b000010101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000001001;
    x_1 = 'b000010000;
    x_2 = 'b000001011;
    x_3 = 'b000001011;
    x_4 = 'b000000110;
    x_5 = 'b111111001;
    x_6 = 'b111101110;
    x_7 = 'b000001001;
    x_8 = 'b000010100;
    x_9 = 'b000011010;
    x_10 = 'b000100100;
    x_11 = 'b000010011;
    x_12 = 'b000010010;
    x_13 = 'b000001010;
    x_14 = 'b000010101;
    x_15 = 'b000011110;
    x_16 = 'b000100000;
    x_17 = 'b000100001;
    x_18 = 'b000100011;
    x_19 = 'b000100100;
    x_20 = 'b000010111;
    x_21 = 'b111110111;
    x_22 = 'b111110100;
    x_23 = 'b111101100;
    x_24 = 'b111101111;
    x_25 = 'b111110000;
    x_26 = 'b111101011;
    x_27 = 'b111101100;
    x_28 = 'b111111011;
    x_29 = 'b111111101;
    x_30 = 'b111110001;
    x_31 = 'b111101110;
    x_32 = 'b111111010;
    x_33 = 'b111110100;
    x_34 = 'b111101011;
    x_35 = 'b111101101;
    x_36 = 'b111100110;
    x_37 = 'b111100111;
    x_38 = 'b111111111;
    x_39 = 'b111110111;
    x_40 = 'b000001000;
    x_41 = 'b111001111;
    x_42 = 'b000001000;
    x_43 = 'b000011110;
    x_44 = 'b111111101;
    x_45 = 'b000101001;
    x_46 = 'b000010010;
    x_47 = 'b000011001;
    x_48 = 'b000010110;
    x_49 = 'b000100110;
    x_50 = 'b000101000;
    x_51 = 'b000101101;
    x_52 = 'b000101001;
    x_53 = 'b000100111;
    x_54 = 'b000100110;
    x_55 = 'b000011101;
    x_56 = 'b000011110;
    x_57 = 'b000110000;
    x_58 = 'b000101110;
    x_59 = 'b000110000;
    x_60 = 'b000101001;
    x_61 = 'b000110011;
    x_62 = 'b000011111;
    x_63 = 'b000011001;

    h_0 = 'b000001001;
    h_1 = 'b000010000;
    h_2 = 'b000001011;
    h_3 = 'b000001011;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111111001;
    x_1 = 'b111111001;
    x_2 = 'b111101111;
    x_3 = 'b111110101;
    x_4 = 'b111111000;
    x_5 = 'b111110100;
    x_6 = 'b111111001;
    x_7 = 'b111111111;
    x_8 = 'b111110010;
    x_9 = 'b111101011;
    x_10 = 'b111101110;
    x_11 = 'b111101101;
    x_12 = 'b111111000;
    x_13 = 'b000000101;
    x_14 = 'b111110010;
    x_15 = 'b111110011;
    x_16 = 'b111101110;
    x_17 = 'b111101100;
    x_18 = 'b111110101;
    x_19 = 'b111110001;
    x_20 = 'b000000110;
    x_21 = 'b000001100;
    x_22 = 'b000001100;
    x_23 = 'b000000111;
    x_24 = 'b000000111;
    x_25 = 'b000000111;
    x_26 = 'b000000011;
    x_27 = 'b111111011;
    x_28 = 'b111110111;
    x_29 = 'b000000010;
    x_30 = 'b000001000;
    x_31 = 'b111111101;
    x_32 = 'b000000010;
    x_33 = 'b111111010;
    x_34 = 'b111111010;
    x_35 = 'b111111100;
    x_36 = 'b111111000;
    x_37 = 'b111111001;
    x_38 = 'b000000000;
    x_39 = 'b000010010;
    x_40 = 'b111111110;
    x_41 = 'b000110001;
    x_42 = 'b111111010;
    x_43 = 'b000010000;
    x_44 = 'b111110000;
    x_45 = 'b000010101;
    x_46 = 'b111101000;
    x_47 = 'b111110011;
    x_48 = 'b111110011;
    x_49 = 'b111110101;
    x_50 = 'b111110011;
    x_51 = 'b111110111;
    x_52 = 'b111110111;
    x_53 = 'b111111110;
    x_54 = 'b000000110;
    x_55 = 'b111101010;
    x_56 = 'b111110101;
    x_57 = 'b111111000;
    x_58 = 'b111111010;
    x_59 = 'b111111001;
    x_60 = 'b111111001;
    x_61 = 'b111110100;
    x_62 = 'b111110101;
    x_63 = 'b000000010;

    h_0 = 'b111111001;
    h_1 = 'b111111001;
    h_2 = 'b111101111;
    h_3 = 'b111110101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b000000001;
    x_1 = 'b000000000;
    x_2 = 'b111110101;
    x_3 = 'b111111101;
    x_4 = 'b111111100;
    x_5 = 'b111110111;
    x_6 = 'b111111010;
    x_7 = 'b000000011;
    x_8 = 'b111110100;
    x_9 = 'b111101110;
    x_10 = 'b111110011;
    x_11 = 'b111110011;
    x_12 = 'b111111010;
    x_13 = 'b000001011;
    x_14 = 'b111110011;
    x_15 = 'b111110000;
    x_16 = 'b111101110;
    x_17 = 'b111101110;
    x_18 = 'b111110101;
    x_19 = 'b111101111;
    x_20 = 'b000000011;
    x_21 = 'b000001101;
    x_22 = 'b000001011;
    x_23 = 'b000000110;
    x_24 = 'b000001000;
    x_25 = 'b000000111;
    x_26 = 'b000000010;
    x_27 = 'b111111100;
    x_28 = 'b111110101;
    x_29 = 'b000000010;
    x_30 = 'b000001000;
    x_31 = 'b111111110;
    x_32 = 'b000000010;
    x_33 = 'b111111001;
    x_34 = 'b111111001;
    x_35 = 'b111111001;
    x_36 = 'b111110111;
    x_37 = 'b111110100;
    x_38 = 'b111111111;
    x_39 = 'b000001001;
    x_40 = 'b111110111;
    x_41 = 'b000000101;
    x_42 = 'b111110011;
    x_43 = 'b000001001;
    x_44 = 'b111101000;
    x_45 = 'b000001010;
    x_46 = 'b111100001;
    x_47 = 'b111101010;
    x_48 = 'b111101011;
    x_49 = 'b111101110;
    x_50 = 'b111101101;
    x_51 = 'b111110000;
    x_52 = 'b111110000;
    x_53 = 'b111110100;
    x_54 = 'b111110111;
    x_55 = 'b111011111;
    x_56 = 'b111101010;
    x_57 = 'b111101111;
    x_58 = 'b111110011;
    x_59 = 'b111110100;
    x_60 = 'b111110010;
    x_61 = 'b111110000;
    x_62 = 'b111110100;
    x_63 = 'b111111101;

    h_0 = 'b000000001;
    h_1 = 'b000000000;
    h_2 = 'b111110101;
    h_3 = 'b111111101;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111110111;
    x_1 = 'b111110101;
    x_2 = 'b111101100;
    x_3 = 'b111110100;
    x_4 = 'b111110011;
    x_5 = 'b111101110;
    x_6 = 'b111101110;
    x_7 = 'b111110101;
    x_8 = 'b111100101;
    x_9 = 'b111100000;
    x_10 = 'b111100110;
    x_11 = 'b111100100;
    x_12 = 'b111101000;
    x_13 = 'b111110010;
    x_14 = 'b111100110;
    x_15 = 'b111011111;
    x_16 = 'b111011100;
    x_17 = 'b111011111;
    x_18 = 'b111100011;
    x_19 = 'b111011010;
    x_20 = 'b111100110;
    x_21 = 'b000001001;
    x_22 = 'b000000111;
    x_23 = 'b000000011;
    x_24 = 'b000000001;
    x_25 = 'b000000001;
    x_26 = 'b111111010;
    x_27 = 'b111110101;
    x_28 = 'b111110000;
    x_29 = 'b111111011;
    x_30 = 'b000000001;
    x_31 = 'b111110101;
    x_32 = 'b111110111;
    x_33 = 'b111101111;
    x_34 = 'b111110000;
    x_35 = 'b111110001;
    x_36 = 'b111101100;
    x_37 = 'b111101100;
    x_38 = 'b111111000;
    x_39 = 'b111110010;
    x_40 = 'b111110001;
    x_41 = 'b111100011;
    x_42 = 'b111101110;
    x_43 = 'b111110110;
    x_44 = 'b111100010;
    x_45 = 'b111100001;
    x_46 = 'b111011001;
    x_47 = 'b111011100;
    x_48 = 'b111011010;
    x_49 = 'b111011001;
    x_50 = 'b111011001;
    x_51 = 'b111011000;
    x_52 = 'b111010101;
    x_53 = 'b111010011;
    x_54 = 'b111001110;
    x_55 = 'b111010011;
    x_56 = 'b111011010;
    x_57 = 'b111011100;
    x_58 = 'b111011100;
    x_59 = 'b111011001;
    x_60 = 'b111100111;
    x_61 = 'b111100011;
    x_62 = 'b111101001;
    x_63 = 'b111110000;

    h_0 = 'b111110111;
    h_1 = 'b111110101;
    h_2 = 'b111101100;
    h_3 = 'b111110100;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    x_0 = 'b111110111;
    x_1 = 'b111110010;
    x_2 = 'b111100101;
    x_3 = 'b111101111;
    x_4 = 'b111101111;
    x_5 = 'b111101001;
    x_6 = 'b111101100;
    x_7 = 'b111111001;
    x_8 = 'b111011111;
    x_9 = 'b111011000;
    x_10 = 'b111011011;
    x_11 = 'b111011000;
    x_12 = 'b111011001;
    x_13 = 'b111100010;
    x_14 = 'b111100111;
    x_15 = 'b111011011;
    x_16 = 'b111010010;
    x_17 = 'b111010011;
    x_18 = 'b111011000;
    x_19 = 'b111001001;
    x_20 = 'b111010010;
    x_21 = 'b000010001;
    x_22 = 'b000010010;
    x_23 = 'b000001101;
    x_24 = 'b000001011;
    x_25 = 'b000001010;
    x_26 = 'b000000110;
    x_27 = 'b000000001;
    x_28 = 'b111111001;
    x_29 = 'b000001001;
    x_30 = 'b000001001;
    x_31 = 'b111111110;
    x_32 = 'b111111110;
    x_33 = 'b111111011;
    x_34 = 'b111111101;
    x_35 = 'b111111101;
    x_36 = 'b111111011;
    x_37 = 'b111111010;
    x_38 = 'b000000110;
    x_39 = 'b111111101;
    x_40 = 'b000000011;
    x_41 = 'b111111000;
    x_42 = 'b000000100;
    x_43 = 'b111011011;
    x_44 = 'b111101001;
    x_45 = 'b111000100;
    x_46 = 'b111011101;
    x_47 = 'b111011100;
    x_48 = 'b111010111;
    x_49 = 'b111010010;
    x_50 = 'b111010000;
    x_51 = 'b111001111;
    x_52 = 'b111001110;
    x_53 = 'b111001000;
    x_54 = 'b111000010;
    x_55 = 'b111001111;
    x_56 = 'b111010010;
    x_57 = 'b111010100;
    x_58 = 'b111010011;
    x_59 = 'b111010000;
    x_60 = 'b111011110;
    x_61 = 'b111011000;
    x_62 = 'b111011110;
    x_63 = 'b111101011;

    h_0 = 'b111110111;
    h_1 = 'b111110010;
    h_2 = 'b111100101;
    h_3 = 'b111101111;
    #20;
    $fdisplay(fd, "%09b %09b %09b %09b", y_0, y_1, y_2, y_3);

    $fclose(fd);    
$finish;
    end
endmodule