`timescale 1ns / 1ps

module gru_tb;

// Parameters
parameter int INT_WIDTH  = 6;
parameter int FRAC_WIDTH = 14;
parameter int WIDTH      = INT_WIDTH + FRAC_WIDTH;
parameter real CLK_PERIOD = 10.0;

// Clock and reset
logic clk;
logic reset;

// Inputs
logic signed [WIDTH-1:0] x_0 = 0;
logic signed [WIDTH-1:0] x_1 = 0;
logic signed [WIDTH-1:0] x_2 = 0;
logic signed [WIDTH-1:0] x_3 = 0;
logic signed [WIDTH-1:0] x_4 = 0;
logic signed [WIDTH-1:0] x_5 = 0;
logic signed [WIDTH-1:0] x_6 = 0;
logic signed [WIDTH-1:0] x_7 = 0;
logic signed [WIDTH-1:0] x_8 = 0;
logic signed [WIDTH-1:0] x_9 = 0;
logic signed [WIDTH-1:0] x_10 = 0;
logic signed [WIDTH-1:0] x_11 = 0;
logic signed [WIDTH-1:0] x_12 = 0;
logic signed [WIDTH-1:0] x_13 = 0;
logic signed [WIDTH-1:0] x_14 = 0;
logic signed [WIDTH-1:0] x_15 = 0;

logic signed [WIDTH-1:0] h_0 = 0;
logic signed [WIDTH-1:0] h_1 = 0;
logic signed [WIDTH-1:0] h_2 = 0;
logic signed [WIDTH-1:0] h_3 = 0;
logic signed [WIDTH-1:0] h_4 = 0;
logic signed [WIDTH-1:0] h_5 = 0;
logic signed [WIDTH-1:0] h_6 = 0;
logic signed [WIDTH-1:0] h_7 = 0;

// Input weights (h×d for each gate)
logic signed [WIDTH-1:0] w_ir_0_0 = 'b00000000010100101000;
logic signed [WIDTH-1:0] w_ir_0_1 = 'b00000000100111000110;
logic signed [WIDTH-1:0] w_ir_0_2 = 'b00000000011101110011;
logic signed [WIDTH-1:0] w_ir_0_3 = 'b00000000100011001100;
logic signed [WIDTH-1:0] w_ir_0_4 = 'b11111111101101001101;
logic signed [WIDTH-1:0] w_ir_0_5 = 'b11111111010101010000;
logic signed [WIDTH-1:0] w_ir_0_6 = 'b00000000011100110100;
logic signed [WIDTH-1:0] w_ir_0_7 = 'b00000000001111011100;
logic signed [WIDTH-1:0] w_ir_0_8 = 'b11111111001000001100;
logic signed [WIDTH-1:0] w_ir_0_9 = 'b00000000000101100110;
logic signed [WIDTH-1:0] w_ir_0_10 = 'b00000000111110110000;
logic signed [WIDTH-1:0] w_ir_0_11 = 'b11111111111111101011;
logic signed [WIDTH-1:0] w_ir_0_12 = 'b00000000100111111110;
logic signed [WIDTH-1:0] w_ir_0_13 = 'b00000000001011000000;
logic signed [WIDTH-1:0] w_ir_0_14 = 'b00000000001001110111;
logic signed [WIDTH-1:0] w_ir_0_15 = 'b00000000101110010111;
logic signed [WIDTH-1:0] w_ir_1_0 = 'b11111111111000000001;
logic signed [WIDTH-1:0] w_ir_1_1 = 'b00000000110111001110;
logic signed [WIDTH-1:0] w_ir_1_2 = 'b11111111111000110010;
logic signed [WIDTH-1:0] w_ir_1_3 = 'b00000000100100010011;
logic signed [WIDTH-1:0] w_ir_1_4 = 'b11111111111000011111;
logic signed [WIDTH-1:0] w_ir_1_5 = 'b00000000100001110010;
logic signed [WIDTH-1:0] w_ir_1_6 = 'b00000000011000100000;
logic signed [WIDTH-1:0] w_ir_1_7 = 'b00000000011000111000;
logic signed [WIDTH-1:0] w_ir_1_8 = 'b11111111010111101111;
logic signed [WIDTH-1:0] w_ir_1_9 = 'b00000000011110000011;
logic signed [WIDTH-1:0] w_ir_1_10 = 'b00000000100010111001;
logic signed [WIDTH-1:0] w_ir_1_11 = 'b00000000010110110101;
logic signed [WIDTH-1:0] w_ir_1_12 = 'b00000000111000101001;
logic signed [WIDTH-1:0] w_ir_1_13 = 'b11111111001011000011;
logic signed [WIDTH-1:0] w_ir_1_14 = 'b11111111101101011000;
logic signed [WIDTH-1:0] w_ir_1_15 = 'b00000000011001110000;
logic signed [WIDTH-1:0] w_ir_2_0 = 'b00000000001100011100;
logic signed [WIDTH-1:0] w_ir_2_1 = 'b00000000011110100011;
logic signed [WIDTH-1:0] w_ir_2_2 = 'b00000000011110100111;
logic signed [WIDTH-1:0] w_ir_2_3 = 'b00000000000110101111;
logic signed [WIDTH-1:0] w_ir_2_4 = 'b00000000111111101011;
logic signed [WIDTH-1:0] w_ir_2_5 = 'b00000000010100010000;
logic signed [WIDTH-1:0] w_ir_2_6 = 'b11111111101110110011;
logic signed [WIDTH-1:0] w_ir_2_7 = 'b00000000001111011001;
logic signed [WIDTH-1:0] w_ir_2_8 = 'b00000000100101011010;
logic signed [WIDTH-1:0] w_ir_2_9 = 'b11111111010000001111;
logic signed [WIDTH-1:0] w_ir_2_10 = 'b00000000001111001110;
logic signed [WIDTH-1:0] w_ir_2_11 = 'b11111111101000010011;
logic signed [WIDTH-1:0] w_ir_2_12 = 'b11111111111110010011;
logic signed [WIDTH-1:0] w_ir_2_13 = 'b11111111011100101001;
logic signed [WIDTH-1:0] w_ir_2_14 = 'b11111111001110100000;
logic signed [WIDTH-1:0] w_ir_2_15 = 'b00000000110111101100;
logic signed [WIDTH-1:0] w_ir_3_0 = 'b11111111110001010100;
logic signed [WIDTH-1:0] w_ir_3_1 = 'b11111111100111001000;
logic signed [WIDTH-1:0] w_ir_3_2 = 'b11111111111001100101;
logic signed [WIDTH-1:0] w_ir_3_3 = 'b00000000000000010010;
logic signed [WIDTH-1:0] w_ir_3_4 = 'b11111111000110110000;
logic signed [WIDTH-1:0] w_ir_3_5 = 'b11111111101010010011;
logic signed [WIDTH-1:0] w_ir_3_6 = 'b00000000010000110011;
logic signed [WIDTH-1:0] w_ir_3_7 = 'b11111111100111110000;
logic signed [WIDTH-1:0] w_ir_3_8 = 'b00000000100110010100;
logic signed [WIDTH-1:0] w_ir_3_9 = 'b11111111100101011001;
logic signed [WIDTH-1:0] w_ir_3_10 = 'b11111111101011011001;
logic signed [WIDTH-1:0] w_ir_3_11 = 'b00000000100010000000;
logic signed [WIDTH-1:0] w_ir_3_12 = 'b11111111010101000001;
logic signed [WIDTH-1:0] w_ir_3_13 = 'b11111111001101111100;
logic signed [WIDTH-1:0] w_ir_3_14 = 'b11111111001100011111;
logic signed [WIDTH-1:0] w_ir_3_15 = 'b00000000100001011101;
logic signed [WIDTH-1:0] w_ir_4_0 = 'b11111111100010111001;
logic signed [WIDTH-1:0] w_ir_4_1 = 'b11111111100110010111;
logic signed [WIDTH-1:0] w_ir_4_2 = 'b00000000101111110101;
logic signed [WIDTH-1:0] w_ir_4_3 = 'b00000000100101100100;
logic signed [WIDTH-1:0] w_ir_4_4 = 'b00000000000101000110;
logic signed [WIDTH-1:0] w_ir_4_5 = 'b00000000001111100011;
logic signed [WIDTH-1:0] w_ir_4_6 = 'b00000000001101001001;
logic signed [WIDTH-1:0] w_ir_4_7 = 'b00000000001000001111;
logic signed [WIDTH-1:0] w_ir_4_8 = 'b00000000001010000001;
logic signed [WIDTH-1:0] w_ir_4_9 = 'b00000000001001010001;
logic signed [WIDTH-1:0] w_ir_4_10 = 'b11111111111000011101;
logic signed [WIDTH-1:0] w_ir_4_11 = 'b11111111111111101100;
logic signed [WIDTH-1:0] w_ir_4_12 = 'b00000000001011101100;
logic signed [WIDTH-1:0] w_ir_4_13 = 'b00000000011100000001;
logic signed [WIDTH-1:0] w_ir_4_14 = 'b11111111010101101000;
logic signed [WIDTH-1:0] w_ir_4_15 = 'b00000000001000100001;
logic signed [WIDTH-1:0] w_ir_5_0 = 'b11111111111111110101;
logic signed [WIDTH-1:0] w_ir_5_1 = 'b11111111111111000111;
logic signed [WIDTH-1:0] w_ir_5_2 = 'b11111111111100100011;
logic signed [WIDTH-1:0] w_ir_5_3 = 'b11111111101011111101;
logic signed [WIDTH-1:0] w_ir_5_4 = 'b11111111111100000100;
logic signed [WIDTH-1:0] w_ir_5_5 = 'b00000000001011011011;
logic signed [WIDTH-1:0] w_ir_5_6 = 'b11111111110000000001;
logic signed [WIDTH-1:0] w_ir_5_7 = 'b11111111101000000001;
logic signed [WIDTH-1:0] w_ir_5_8 = 'b00000000000000010100;
logic signed [WIDTH-1:0] w_ir_5_9 = 'b00000000101110100100;
logic signed [WIDTH-1:0] w_ir_5_10 = 'b11111111001100101001;
logic signed [WIDTH-1:0] w_ir_5_11 = 'b11111111001110101000;
logic signed [WIDTH-1:0] w_ir_5_12 = 'b00000000110101101000;
logic signed [WIDTH-1:0] w_ir_5_13 = 'b00000000010000010100;
logic signed [WIDTH-1:0] w_ir_5_14 = 'b00000000000011101001;
logic signed [WIDTH-1:0] w_ir_5_15 = 'b11111111111111011010;
logic signed [WIDTH-1:0] w_ir_6_0 = 'b11111111100001010010;
logic signed [WIDTH-1:0] w_ir_6_1 = 'b11111111111101001000;
logic signed [WIDTH-1:0] w_ir_6_2 = 'b11111111111011010100;
logic signed [WIDTH-1:0] w_ir_6_3 = 'b00000000000011110001;
logic signed [WIDTH-1:0] w_ir_6_4 = 'b00000000001111101100;
logic signed [WIDTH-1:0] w_ir_6_5 = 'b00000000001001000101;
logic signed [WIDTH-1:0] w_ir_6_6 = 'b00000000001100100101;
logic signed [WIDTH-1:0] w_ir_6_7 = 'b00000000100000000101;
logic signed [WIDTH-1:0] w_ir_6_8 = 'b00000000010011010100;
logic signed [WIDTH-1:0] w_ir_6_9 = 'b00000000000000011001;
logic signed [WIDTH-1:0] w_ir_6_10 = 'b11111111111101010100;
logic signed [WIDTH-1:0] w_ir_6_11 = 'b00000000010000001101;
logic signed [WIDTH-1:0] w_ir_6_12 = 'b00000000000110001011;
logic signed [WIDTH-1:0] w_ir_6_13 = 'b00000000001100100111;
logic signed [WIDTH-1:0] w_ir_6_14 = 'b11111111111100111100;
logic signed [WIDTH-1:0] w_ir_6_15 = 'b11111111110111000110;
logic signed [WIDTH-1:0] w_ir_7_0 = 'b11111111110110110111;
logic signed [WIDTH-1:0] w_ir_7_1 = 'b11111111001010111010;
logic signed [WIDTH-1:0] w_ir_7_2 = 'b00000000011110100101;
logic signed [WIDTH-1:0] w_ir_7_3 = 'b00000000101010101011;
logic signed [WIDTH-1:0] w_ir_7_4 = 'b11111111110011100010;
logic signed [WIDTH-1:0] w_ir_7_5 = 'b11111111100111011010;
logic signed [WIDTH-1:0] w_ir_7_6 = 'b11111111101000000000;
logic signed [WIDTH-1:0] w_ir_7_7 = 'b11111111100100110111;
logic signed [WIDTH-1:0] w_ir_7_8 = 'b11111111110000011001;
logic signed [WIDTH-1:0] w_ir_7_9 = 'b00000000110010110111;
logic signed [WIDTH-1:0] w_ir_7_10 = 'b00000000011101110100;
logic signed [WIDTH-1:0] w_ir_7_11 = 'b11111111011111000110;
logic signed [WIDTH-1:0] w_ir_7_12 = 'b11111111110111100111;
logic signed [WIDTH-1:0] w_ir_7_13 = 'b11111111110010011010;
logic signed [WIDTH-1:0] w_ir_7_14 = 'b00000000101011000011;
logic signed [WIDTH-1:0] w_ir_7_15 = 'b11111111100111101111;

logic signed [WIDTH-1:0] w_iz_0_0 = 'b11111111101001001000;
logic signed [WIDTH-1:0] w_iz_0_1 = 'b11111111110000000111;
logic signed [WIDTH-1:0] w_iz_0_2 = 'b11111111001001100001;
logic signed [WIDTH-1:0] w_iz_0_3 = 'b11111111011110001110;
logic signed [WIDTH-1:0] w_iz_0_4 = 'b11111111101101011001;
logic signed [WIDTH-1:0] w_iz_0_5 = 'b11111111110111010111;
logic signed [WIDTH-1:0] w_iz_0_6 = 'b00000000000101111000;
logic signed [WIDTH-1:0] w_iz_0_7 = 'b11111111010111011001;
logic signed [WIDTH-1:0] w_iz_0_8 = 'b11111111110101000011;
logic signed [WIDTH-1:0] w_iz_0_9 = 'b11111111110101100001;
logic signed [WIDTH-1:0] w_iz_0_10 = 'b11111111110100000111;
logic signed [WIDTH-1:0] w_iz_0_11 = 'b11111111000101100111;
logic signed [WIDTH-1:0] w_iz_0_12 = 'b11111111110110101111;
logic signed [WIDTH-1:0] w_iz_0_13 = 'b00000000001101111001;
logic signed [WIDTH-1:0] w_iz_0_14 = 'b11111111110101000010;
logic signed [WIDTH-1:0] w_iz_0_15 = 'b00000000010101111110;
logic signed [WIDTH-1:0] w_iz_1_0 = 'b11111111010110100000;
logic signed [WIDTH-1:0] w_iz_1_1 = 'b00000000111001010110;
logic signed [WIDTH-1:0] w_iz_1_2 = 'b00000000000011000000;
logic signed [WIDTH-1:0] w_iz_1_3 = 'b00000000010010111101;
logic signed [WIDTH-1:0] w_iz_1_4 = 'b00000000001101111011;
logic signed [WIDTH-1:0] w_iz_1_5 = 'b11111111101101111110;
logic signed [WIDTH-1:0] w_iz_1_6 = 'b00000000011101111101;
logic signed [WIDTH-1:0] w_iz_1_7 = 'b00000000110100111111;
logic signed [WIDTH-1:0] w_iz_1_8 = 'b00000000011011000000;
logic signed [WIDTH-1:0] w_iz_1_9 = 'b00000000001000110101;
logic signed [WIDTH-1:0] w_iz_1_10 = 'b11111111111100000100;
logic signed [WIDTH-1:0] w_iz_1_11 = 'b11111111001011011011;
logic signed [WIDTH-1:0] w_iz_1_12 = 'b11111111110000111100;
logic signed [WIDTH-1:0] w_iz_1_13 = 'b00000000111100010101;
logic signed [WIDTH-1:0] w_iz_1_14 = 'b11111111100111111110;
logic signed [WIDTH-1:0] w_iz_1_15 = 'b11111111101000010000;
logic signed [WIDTH-1:0] w_iz_2_0 = 'b00000000000010101101;
logic signed [WIDTH-1:0] w_iz_2_1 = 'b00000000010110111101;
logic signed [WIDTH-1:0] w_iz_2_2 = 'b11111111110100010011;
logic signed [WIDTH-1:0] w_iz_2_3 = 'b11111111110010011110;
logic signed [WIDTH-1:0] w_iz_2_4 = 'b00000000000011000100;
logic signed [WIDTH-1:0] w_iz_2_5 = 'b00000000001010100110;
logic signed [WIDTH-1:0] w_iz_2_6 = 'b00000000100000000011;
logic signed [WIDTH-1:0] w_iz_2_7 = 'b11111111111111101010;
logic signed [WIDTH-1:0] w_iz_2_8 = 'b00000000011100011110;
logic signed [WIDTH-1:0] w_iz_2_9 = 'b11111111110010101011;
logic signed [WIDTH-1:0] w_iz_2_10 = 'b00000000011101100110;
logic signed [WIDTH-1:0] w_iz_2_11 = 'b11111111111100110010;
logic signed [WIDTH-1:0] w_iz_2_12 = 'b00000000001011010000;
logic signed [WIDTH-1:0] w_iz_2_13 = 'b00000000001111110101;
logic signed [WIDTH-1:0] w_iz_2_14 = 'b00000000001100011110;
logic signed [WIDTH-1:0] w_iz_2_15 = 'b00000000000110011111;
logic signed [WIDTH-1:0] w_iz_3_0 = 'b00000000001100111001;
logic signed [WIDTH-1:0] w_iz_3_1 = 'b00000000001010110101;
logic signed [WIDTH-1:0] w_iz_3_2 = 'b11111111100001100000;
logic signed [WIDTH-1:0] w_iz_3_3 = 'b00000000010101110000;
logic signed [WIDTH-1:0] w_iz_3_4 = 'b00000000010100100000;
logic signed [WIDTH-1:0] w_iz_3_5 = 'b00000000001110010001;
logic signed [WIDTH-1:0] w_iz_3_6 = 'b11111111001001010010;
logic signed [WIDTH-1:0] w_iz_3_7 = 'b00000000010010110010;
logic signed [WIDTH-1:0] w_iz_3_8 = 'b00000000001100100010;
logic signed [WIDTH-1:0] w_iz_3_9 = 'b11111111010111001110;
logic signed [WIDTH-1:0] w_iz_3_10 = 'b11111111100001111100;
logic signed [WIDTH-1:0] w_iz_3_11 = 'b11111111100101100101;
logic signed [WIDTH-1:0] w_iz_3_12 = 'b00000000100110010110;
logic signed [WIDTH-1:0] w_iz_3_13 = 'b00000000010001100011;
logic signed [WIDTH-1:0] w_iz_3_14 = 'b00000000100111110010;
logic signed [WIDTH-1:0] w_iz_3_15 = 'b00000001000110100101;
logic signed [WIDTH-1:0] w_iz_4_0 = 'b11111111111101110111;
logic signed [WIDTH-1:0] w_iz_4_1 = 'b00000000111111011000;
logic signed [WIDTH-1:0] w_iz_4_2 = 'b00000000000000001000;
logic signed [WIDTH-1:0] w_iz_4_3 = 'b00000000110010101000;
logic signed [WIDTH-1:0] w_iz_4_4 = 'b11111111010010000001;
logic signed [WIDTH-1:0] w_iz_4_5 = 'b00000000001010010110;
logic signed [WIDTH-1:0] w_iz_4_6 = 'b00000000000111101000;
logic signed [WIDTH-1:0] w_iz_4_7 = 'b11111111101100110101;
logic signed [WIDTH-1:0] w_iz_4_8 = 'b11111111111000110011;
logic signed [WIDTH-1:0] w_iz_4_9 = 'b00000000101001101011;
logic signed [WIDTH-1:0] w_iz_4_10 = 'b11111111100010011010;
logic signed [WIDTH-1:0] w_iz_4_11 = 'b11111111111010011111;
logic signed [WIDTH-1:0] w_iz_4_12 = 'b11111111011111101010;
logic signed [WIDTH-1:0] w_iz_4_13 = 'b11111111110101001010;
logic signed [WIDTH-1:0] w_iz_4_14 = 'b11111111110001111011;
logic signed [WIDTH-1:0] w_iz_4_15 = 'b11111111111000110001;
logic signed [WIDTH-1:0] w_iz_5_0 = 'b00000000000010011011;
logic signed [WIDTH-1:0] w_iz_5_1 = 'b00000000001010101110;
logic signed [WIDTH-1:0] w_iz_5_2 = 'b11111111101001110010;
logic signed [WIDTH-1:0] w_iz_5_3 = 'b00000000100000011111;
logic signed [WIDTH-1:0] w_iz_5_4 = 'b11111111110011000001;
logic signed [WIDTH-1:0] w_iz_5_5 = 'b00000000001100110101;
logic signed [WIDTH-1:0] w_iz_5_6 = 'b00000000010101000111;
logic signed [WIDTH-1:0] w_iz_5_7 = 'b00000000001101101000;
logic signed [WIDTH-1:0] w_iz_5_8 = 'b00000000110101000101;
logic signed [WIDTH-1:0] w_iz_5_9 = 'b00000000001011101001;
logic signed [WIDTH-1:0] w_iz_5_10 = 'b11111111111000100001;
logic signed [WIDTH-1:0] w_iz_5_11 = 'b11111111101100101011;
logic signed [WIDTH-1:0] w_iz_5_12 = 'b00000000001011010100;
logic signed [WIDTH-1:0] w_iz_5_13 = 'b00000000001001100010;
logic signed [WIDTH-1:0] w_iz_5_14 = 'b11111111011110000001;
logic signed [WIDTH-1:0] w_iz_5_15 = 'b00000001000010001111;
logic signed [WIDTH-1:0] w_iz_6_0 = 'b00000000100001111100;
logic signed [WIDTH-1:0] w_iz_6_1 = 'b11111111011000100111;
logic signed [WIDTH-1:0] w_iz_6_2 = 'b00000000010000000011;
logic signed [WIDTH-1:0] w_iz_6_3 = 'b00000000001001001101;
logic signed [WIDTH-1:0] w_iz_6_4 = 'b00000000001011110000;
logic signed [WIDTH-1:0] w_iz_6_5 = 'b11111111000111111010;
logic signed [WIDTH-1:0] w_iz_6_6 = 'b00000000011000100100;
logic signed [WIDTH-1:0] w_iz_6_7 = 'b00000000000011100111;
logic signed [WIDTH-1:0] w_iz_6_8 = 'b11111111111110110100;
logic signed [WIDTH-1:0] w_iz_6_9 = 'b00000000100101010101;
logic signed [WIDTH-1:0] w_iz_6_10 = 'b11111111010110001101;
logic signed [WIDTH-1:0] w_iz_6_11 = 'b00000000000110000100;
logic signed [WIDTH-1:0] w_iz_6_12 = 'b11111111101001111111;
logic signed [WIDTH-1:0] w_iz_6_13 = 'b11111111101110001001;
logic signed [WIDTH-1:0] w_iz_6_14 = 'b00000000110001011110;
logic signed [WIDTH-1:0] w_iz_6_15 = 'b11111111101000111000;
logic signed [WIDTH-1:0] w_iz_7_0 = 'b11111111110010100010;
logic signed [WIDTH-1:0] w_iz_7_1 = 'b11111111110110011000;
logic signed [WIDTH-1:0] w_iz_7_2 = 'b11111111100011111111;
logic signed [WIDTH-1:0] w_iz_7_3 = 'b11111111101000000101;
logic signed [WIDTH-1:0] w_iz_7_4 = 'b11111111100101111010;
logic signed [WIDTH-1:0] w_iz_7_5 = 'b11111111100010110101;
logic signed [WIDTH-1:0] w_iz_7_6 = 'b11111111101111011000;
logic signed [WIDTH-1:0] w_iz_7_7 = 'b11111111000110000010;
logic signed [WIDTH-1:0] w_iz_7_8 = 'b11111111100100110010;
logic signed [WIDTH-1:0] w_iz_7_9 = 'b00000000011111001110;
logic signed [WIDTH-1:0] w_iz_7_10 = 'b11111111011100111000;
logic signed [WIDTH-1:0] w_iz_7_11 = 'b11111111100111000111;
logic signed [WIDTH-1:0] w_iz_7_12 = 'b11111111100111111111;
logic signed [WIDTH-1:0] w_iz_7_13 = 'b11111111101011010101;
logic signed [WIDTH-1:0] w_iz_7_14 = 'b11111111010000010010;
logic signed [WIDTH-1:0] w_iz_7_15 = 'b11111111101100000011;

logic signed [WIDTH-1:0] w_in_0_0 = 'b11111111111100100000;
logic signed [WIDTH-1:0] w_in_0_1 = 'b11111111110011011010;
logic signed [WIDTH-1:0] w_in_0_2 = 'b11111111110110101110;
logic signed [WIDTH-1:0] w_in_0_3 = 'b11111111100111001111;
logic signed [WIDTH-1:0] w_in_0_4 = 'b00000000000001010001;
logic signed [WIDTH-1:0] w_in_0_5 = 'b00000000010111000110;
logic signed [WIDTH-1:0] w_in_0_6 = 'b11111111100011010111;
logic signed [WIDTH-1:0] w_in_0_7 = 'b11111111010111010010;
logic signed [WIDTH-1:0] w_in_0_8 = 'b11111111000101000000;
logic signed [WIDTH-1:0] w_in_0_9 = 'b11111111101001011001;
logic signed [WIDTH-1:0] w_in_0_10 = 'b11111111001011100001;
logic signed [WIDTH-1:0] w_in_0_11 = 'b11111111101111000010;
logic signed [WIDTH-1:0] w_in_0_12 = 'b11111111110110100110;
logic signed [WIDTH-1:0] w_in_0_13 = 'b00000000010111000011;
logic signed [WIDTH-1:0] w_in_0_14 = 'b00000000000110010010;
logic signed [WIDTH-1:0] w_in_0_15 = 'b11111111110110100101;
logic signed [WIDTH-1:0] w_in_1_0 = 'b11111111100000110100;
logic signed [WIDTH-1:0] w_in_1_1 = 'b11111111101000100110;
logic signed [WIDTH-1:0] w_in_1_2 = 'b11111111100001100110;
logic signed [WIDTH-1:0] w_in_1_3 = 'b11111111011010100111;
logic signed [WIDTH-1:0] w_in_1_4 = 'b11111111110111001000;
logic signed [WIDTH-1:0] w_in_1_5 = 'b00000000011010110011;
logic signed [WIDTH-1:0] w_in_1_6 = 'b00000001000011101101;
logic signed [WIDTH-1:0] w_in_1_7 = 'b00000000100101011111;
logic signed [WIDTH-1:0] w_in_1_8 = 'b11111111001000001001;
logic signed [WIDTH-1:0] w_in_1_9 = 'b11111111010010110101;
logic signed [WIDTH-1:0] w_in_1_10 = 'b00000000000011101001;
logic signed [WIDTH-1:0] w_in_1_11 = 'b11111111001000000110;
logic signed [WIDTH-1:0] w_in_1_12 = 'b00000000101111100100;
logic signed [WIDTH-1:0] w_in_1_13 = 'b11111111111101101100;
logic signed [WIDTH-1:0] w_in_1_14 = 'b00000000101101011110;
logic signed [WIDTH-1:0] w_in_1_15 = 'b11111111100001001001;
logic signed [WIDTH-1:0] w_in_2_0 = 'b11111111001100000000;
logic signed [WIDTH-1:0] w_in_2_1 = 'b11111111010010101011;
logic signed [WIDTH-1:0] w_in_2_2 = 'b11111111100001100100;
logic signed [WIDTH-1:0] w_in_2_3 = 'b11111111011110111001;
logic signed [WIDTH-1:0] w_in_2_4 = 'b11111111001101100111;
logic signed [WIDTH-1:0] w_in_2_5 = 'b11111111010101010111;
logic signed [WIDTH-1:0] w_in_2_6 = 'b11111111100100100001;
logic signed [WIDTH-1:0] w_in_2_7 = 'b00000000010001001110;
logic signed [WIDTH-1:0] w_in_2_8 = 'b00000000001011111111;
logic signed [WIDTH-1:0] w_in_2_9 = 'b11111111100011000111;
logic signed [WIDTH-1:0] w_in_2_10 = 'b11111111111011111010;
logic signed [WIDTH-1:0] w_in_2_11 = 'b11111111101001111010;
logic signed [WIDTH-1:0] w_in_2_12 = 'b11111111000010001110;
logic signed [WIDTH-1:0] w_in_2_13 = 'b11111111110101011111;
logic signed [WIDTH-1:0] w_in_2_14 = 'b11111111110101010010;
logic signed [WIDTH-1:0] w_in_2_15 = 'b11111111111000010110;
logic signed [WIDTH-1:0] w_in_3_0 = 'b00000000000000001001;
logic signed [WIDTH-1:0] w_in_3_1 = 'b11111111110010011110;
logic signed [WIDTH-1:0] w_in_3_2 = 'b00000000101001110011;
logic signed [WIDTH-1:0] w_in_3_3 = 'b11111111100110111110;
logic signed [WIDTH-1:0] w_in_3_4 = 'b00000000111010100011;
logic signed [WIDTH-1:0] w_in_3_5 = 'b00000000011100010100;
logic signed [WIDTH-1:0] w_in_3_6 = 'b00000000111101100010;
logic signed [WIDTH-1:0] w_in_3_7 = 'b00000000110011010110;
logic signed [WIDTH-1:0] w_in_3_8 = 'b00000000010100000100;
logic signed [WIDTH-1:0] w_in_3_9 = 'b11111111001000011110;
logic signed [WIDTH-1:0] w_in_3_10 = 'b00000000100000110101;
logic signed [WIDTH-1:0] w_in_3_11 = 'b00000001101110110100;
logic signed [WIDTH-1:0] w_in_3_12 = 'b00000001010010110011;
logic signed [WIDTH-1:0] w_in_3_13 = 'b00000001010111010110;
logic signed [WIDTH-1:0] w_in_3_14 = 'b00000001100111001001;
logic signed [WIDTH-1:0] w_in_3_15 = 'b00000001011100000010;
logic signed [WIDTH-1:0] w_in_4_0 = 'b00000000001010100010;
logic signed [WIDTH-1:0] w_in_4_1 = 'b00000000001011010101;
logic signed [WIDTH-1:0] w_in_4_2 = 'b00000000001101011000;
logic signed [WIDTH-1:0] w_in_4_3 = 'b11111111111000001110;
logic signed [WIDTH-1:0] w_in_4_4 = 'b11111111110111011000;
logic signed [WIDTH-1:0] w_in_4_5 = 'b11111111011011000010;
logic signed [WIDTH-1:0] w_in_4_6 = 'b00000000110001110101;
logic signed [WIDTH-1:0] w_in_4_7 = 'b11111111000101010100;
logic signed [WIDTH-1:0] w_in_4_8 = 'b11111111010010011101;
logic signed [WIDTH-1:0] w_in_4_9 = 'b11111111101111011001;
logic signed [WIDTH-1:0] w_in_4_10 = 'b11111111111110101001;
logic signed [WIDTH-1:0] w_in_4_11 = 'b11111111110110100111;
logic signed [WIDTH-1:0] w_in_4_12 = 'b11111111011100001011;
logic signed [WIDTH-1:0] w_in_4_13 = 'b11111111110101100001;
logic signed [WIDTH-1:0] w_in_4_14 = 'b11111111100000111100;
logic signed [WIDTH-1:0] w_in_4_15 = 'b11111111011111110110;
logic signed [WIDTH-1:0] w_in_5_0 = 'b00000000100100111110;
logic signed [WIDTH-1:0] w_in_5_1 = 'b11111111010111110001;
logic signed [WIDTH-1:0] w_in_5_2 = 'b00000000000111101111;
logic signed [WIDTH-1:0] w_in_5_3 = 'b11111111001101111011;
logic signed [WIDTH-1:0] w_in_5_4 = 'b11111111110110000001;
logic signed [WIDTH-1:0] w_in_5_5 = 'b00000000000001010111;
logic signed [WIDTH-1:0] w_in_5_6 = 'b00000000010100100111;
logic signed [WIDTH-1:0] w_in_5_7 = 'b00000000001100110111;
logic signed [WIDTH-1:0] w_in_5_8 = 'b11111111111010111111;
logic signed [WIDTH-1:0] w_in_5_9 = 'b11111111100111100111;
logic signed [WIDTH-1:0] w_in_5_10 = 'b11111111111011001111;
logic signed [WIDTH-1:0] w_in_5_11 = 'b00000000010111001101;
logic signed [WIDTH-1:0] w_in_5_12 = 'b00000000000101000000;
logic signed [WIDTH-1:0] w_in_5_13 = 'b11111111100010100001;
logic signed [WIDTH-1:0] w_in_5_14 = 'b11111111110001000100;
logic signed [WIDTH-1:0] w_in_5_15 = 'b11111111001000100001;
logic signed [WIDTH-1:0] w_in_6_0 = 'b11111111111100010110;
logic signed [WIDTH-1:0] w_in_6_1 = 'b11111111000000000100;
logic signed [WIDTH-1:0] w_in_6_2 = 'b11111111101111110110;
logic signed [WIDTH-1:0] w_in_6_3 = 'b00000000011111001001;
logic signed [WIDTH-1:0] w_in_6_4 = 'b11111111100000100000;
logic signed [WIDTH-1:0] w_in_6_5 = 'b11111111010001000111;
logic signed [WIDTH-1:0] w_in_6_6 = 'b11111110111010010101;
logic signed [WIDTH-1:0] w_in_6_7 = 'b00000000101000111000;
logic signed [WIDTH-1:0] w_in_6_8 = 'b11111111101011101010;
logic signed [WIDTH-1:0] w_in_6_9 = 'b11111111110111111111;
logic signed [WIDTH-1:0] w_in_6_10 = 'b00000000000011011011;
logic signed [WIDTH-1:0] w_in_6_11 = 'b11111111101001100011;
logic signed [WIDTH-1:0] w_in_6_12 = 'b00000000001000010010;
logic signed [WIDTH-1:0] w_in_6_13 = 'b11111111101010100000;
logic signed [WIDTH-1:0] w_in_6_14 = 'b11111111110110110011;
logic signed [WIDTH-1:0] w_in_6_15 = 'b00000000011110100010;
logic signed [WIDTH-1:0] w_in_7_0 = 'b00000000001111001110;
logic signed [WIDTH-1:0] w_in_7_1 = 'b00000000001100100001;
logic signed [WIDTH-1:0] w_in_7_2 = 'b00000000001010101010;
logic signed [WIDTH-1:0] w_in_7_3 = 'b00000000001011000111;
logic signed [WIDTH-1:0] w_in_7_4 = 'b11111111101110110010;
logic signed [WIDTH-1:0] w_in_7_5 = 'b11111111101011011110;
logic signed [WIDTH-1:0] w_in_7_6 = 'b00000000001110101001;
logic signed [WIDTH-1:0] w_in_7_7 = 'b00000000000000001011;
logic signed [WIDTH-1:0] w_in_7_8 = 'b00000000001011000011;
logic signed [WIDTH-1:0] w_in_7_9 = 'b11111111011011111000;
logic signed [WIDTH-1:0] w_in_7_10 = 'b11111111011110011010;
logic signed [WIDTH-1:0] w_in_7_11 = 'b11111111101101100010;
logic signed [WIDTH-1:0] w_in_7_12 = 'b00000000111011101010;
logic signed [WIDTH-1:0] w_in_7_13 = 'b00000000101000011101;
logic signed [WIDTH-1:0] w_in_7_14 = 'b11111111101100000011;
logic signed [WIDTH-1:0] w_in_7_15 = 'b00000000100100001110;

// Recurrent weights (h×h for each gate)
logic signed [WIDTH-1:0] w_hr_0_0 = 'b00000000000011100100;
logic signed [WIDTH-1:0] w_hr_0_1 = 'b00000000001001101010;
logic signed [WIDTH-1:0] w_hr_0_2 = 'b00000000001111100111;
logic signed [WIDTH-1:0] w_hr_0_3 = 'b11111111010111000111;
logic signed [WIDTH-1:0] w_hr_0_4 = 'b00000001000110000100;
logic signed [WIDTH-1:0] w_hr_0_5 = 'b00000001001011010111;
logic signed [WIDTH-1:0] w_hr_0_6 = 'b00000001001010101110;
logic signed [WIDTH-1:0] w_hr_0_7 = 'b11111110110110001000;
logic signed [WIDTH-1:0] w_hr_1_0 = 'b00000000111111100001;
logic signed [WIDTH-1:0] w_hr_1_1 = 'b00000001000111111010;
logic signed [WIDTH-1:0] w_hr_1_2 = 'b11111111011111011100;
logic signed [WIDTH-1:0] w_hr_1_3 = 'b11111111011000110111;
logic signed [WIDTH-1:0] w_hr_1_4 = 'b00000000011111010000;
logic signed [WIDTH-1:0] w_hr_1_5 = 'b00000000100111111110;
logic signed [WIDTH-1:0] w_hr_1_6 = 'b00000001011010000100;
logic signed [WIDTH-1:0] w_hr_1_7 = 'b11111111000011010010;
logic signed [WIDTH-1:0] w_hr_2_0 = 'b00000000110110111110;
logic signed [WIDTH-1:0] w_hr_2_1 = 'b00000000011100101000;
logic signed [WIDTH-1:0] w_hr_2_2 = 'b11111111101011000100;
logic signed [WIDTH-1:0] w_hr_2_3 = 'b00000000100000100111;
logic signed [WIDTH-1:0] w_hr_2_4 = 'b00000001101000010011;
logic signed [WIDTH-1:0] w_hr_2_5 = 'b11111110011110010001;
logic signed [WIDTH-1:0] w_hr_2_6 = 'b00000000000001101010;
logic signed [WIDTH-1:0] w_hr_2_7 = 'b00000001000111101101;
logic signed [WIDTH-1:0] w_hr_3_0 = 'b00000000110110010110;
logic signed [WIDTH-1:0] w_hr_3_1 = 'b00000000000001010101;
logic signed [WIDTH-1:0] w_hr_3_2 = 'b11111110000010100100;
logic signed [WIDTH-1:0] w_hr_3_3 = 'b00000001110001110110;
logic signed [WIDTH-1:0] w_hr_3_4 = 'b00000001011111101110;
logic signed [WIDTH-1:0] w_hr_3_5 = 'b00000000100010111000;
logic signed [WIDTH-1:0] w_hr_3_6 = 'b11111110110100110001;
logic signed [WIDTH-1:0] w_hr_3_7 = 'b00000010100101110110;
logic signed [WIDTH-1:0] w_hr_4_0 = 'b11111111110101110100;
logic signed [WIDTH-1:0] w_hr_4_1 = 'b11111111101100110010;
logic signed [WIDTH-1:0] w_hr_4_2 = 'b00000000100100011000;
logic signed [WIDTH-1:0] w_hr_4_3 = 'b11111111001100010110;
logic signed [WIDTH-1:0] w_hr_4_4 = 'b11111111010010110100;
logic signed [WIDTH-1:0] w_hr_4_5 = 'b11111111111001110101;
logic signed [WIDTH-1:0] w_hr_4_6 = 'b00000010111011100001;
logic signed [WIDTH-1:0] w_hr_4_7 = 'b11111110100010000101;
logic signed [WIDTH-1:0] w_hr_5_0 = 'b11111111110101110010;
logic signed [WIDTH-1:0] w_hr_5_1 = 'b00000001101100111000;
logic signed [WIDTH-1:0] w_hr_5_2 = 'b00000010011111000111;
logic signed [WIDTH-1:0] w_hr_5_3 = 'b11111110010000010100;
logic signed [WIDTH-1:0] w_hr_5_4 = 'b11111111010110010110;
logic signed [WIDTH-1:0] w_hr_5_5 = 'b11111110110011000110;
logic signed [WIDTH-1:0] w_hr_5_6 = 'b11111111001011100001;
logic signed [WIDTH-1:0] w_hr_5_7 = 'b00000001001110101011;
logic signed [WIDTH-1:0] w_hr_6_0 = 'b00000000000011100100;
logic signed [WIDTH-1:0] w_hr_6_1 = 'b00000000001001101010;
logic signed [WIDTH-1:0] w_hr_6_2 = 'b00000000001111100111;
logic signed [WIDTH-1:0] w_hr_6_3 = 'b11111111010111000111;
logic signed [WIDTH-1:0] w_hr_6_4 = 'b00000001000110000100;
logic signed [WIDTH-1:0] w_hr_6_5 = 'b00000001001011010111;
logic signed [WIDTH-1:0] w_hr_6_6 = 'b00000001001010101110;
logic signed [WIDTH-1:0] w_hr_6_7 = 'b11111110110110001000;
logic signed [WIDTH-1:0] w_hr_7_0 = 'b00000000111111100001;
logic signed [WIDTH-1:0] w_hr_7_1 = 'b00000001000111111010;
logic signed [WIDTH-1:0] w_hr_7_2 = 'b11111111011111011100;
logic signed [WIDTH-1:0] w_hr_7_3 = 'b11111111011000110111;
logic signed [WIDTH-1:0] w_hr_7_4 = 'b00000000011111010000;
logic signed [WIDTH-1:0] w_hr_7_5 = 'b00000000100111111110;
logic signed [WIDTH-1:0] w_hr_7_6 = 'b00000001011010000100;
logic signed [WIDTH-1:0] w_hr_7_7 = 'b11111111000011010010;

logic signed [WIDTH-1:0] w_hz_0_0 = 'b00000000110110111110;
logic signed [WIDTH-1:0] w_hz_0_1 = 'b00000000011100101000;
logic signed [WIDTH-1:0] w_hz_0_2 = 'b11111111101011000100;
logic signed [WIDTH-1:0] w_hz_0_3 = 'b00000000100000100111;
logic signed [WIDTH-1:0] w_hz_0_4 = 'b00000001101000010011;
logic signed [WIDTH-1:0] w_hz_0_5 = 'b11111110011110010001;
logic signed [WIDTH-1:0] w_hz_0_6 = 'b00000000000001101010;
logic signed [WIDTH-1:0] w_hz_0_7 = 'b00000001000111101101;
logic signed [WIDTH-1:0] w_hz_1_0 = 'b00000000110110010110;
logic signed [WIDTH-1:0] w_hz_1_1 = 'b00000000000001010101;
logic signed [WIDTH-1:0] w_hz_1_2 = 'b11111110000010100100;
logic signed [WIDTH-1:0] w_hz_1_3 = 'b00000001110001110110;
logic signed [WIDTH-1:0] w_hz_1_4 = 'b00000001011111101110;
logic signed [WIDTH-1:0] w_hz_1_5 = 'b00000000100010111000;
logic signed [WIDTH-1:0] w_hz_1_6 = 'b11111110110100110001;
logic signed [WIDTH-1:0] w_hz_1_7 = 'b00000010100101110110;
logic signed [WIDTH-1:0] w_hz_2_0 = 'b11111111110101110100;
logic signed [WIDTH-1:0] w_hz_2_1 = 'b11111111101100110010;
logic signed [WIDTH-1:0] w_hz_2_2 = 'b00000000100100011000;
logic signed [WIDTH-1:0] w_hz_2_3 = 'b11111111001100010110;
logic signed [WIDTH-1:0] w_hz_2_4 = 'b11111111010010110100;
logic signed [WIDTH-1:0] w_hz_2_5 = 'b11111111111001110101;
logic signed [WIDTH-1:0] w_hz_2_6 = 'b00000010111011100001;
logic signed [WIDTH-1:0] w_hz_2_7 = 'b11111110100010000101;
logic signed [WIDTH-1:0] w_hz_3_0 = 'b11111111110101110010;
logic signed [WIDTH-1:0] w_hz_3_1 = 'b00000001101100111000;
logic signed [WIDTH-1:0] w_hz_3_2 = 'b00000010011111000111;
logic signed [WIDTH-1:0] w_hz_3_3 = 'b11111110010000010100;
logic signed [WIDTH-1:0] w_hz_3_4 = 'b11111111010110010110;
logic signed [WIDTH-1:0] w_hz_3_5 = 'b11111110110011000110;
logic signed [WIDTH-1:0] w_hz_3_6 = 'b11111111001011100001;
logic signed [WIDTH-1:0] w_hz_3_7 = 'b00000001001110101011;
logic signed [WIDTH-1:0] w_hz_4_0 = 'b00000000000011100100;
logic signed [WIDTH-1:0] w_hz_4_1 = 'b00000000001001101010;
logic signed [WIDTH-1:0] w_hz_4_2 = 'b00000000001111100111;
logic signed [WIDTH-1:0] w_hz_4_3 = 'b11111111010111000111;
logic signed [WIDTH-1:0] w_hz_4_4 = 'b00000001000110000100;
logic signed [WIDTH-1:0] w_hz_4_5 = 'b00000001001011010111;
logic signed [WIDTH-1:0] w_hz_4_6 = 'b00000001001010101110;
logic signed [WIDTH-1:0] w_hz_4_7 = 'b11111110110110001000;
logic signed [WIDTH-1:0] w_hz_5_0 = 'b00000000111111100001;
logic signed [WIDTH-1:0] w_hz_5_1 = 'b00000001000111111010;
logic signed [WIDTH-1:0] w_hz_5_2 = 'b11111111011111011100;
logic signed [WIDTH-1:0] w_hz_5_3 = 'b11111111011000110111;
logic signed [WIDTH-1:0] w_hz_5_4 = 'b00000000011111010000;
logic signed [WIDTH-1:0] w_hz_5_5 = 'b00000000100111111110;
logic signed [WIDTH-1:0] w_hz_5_6 = 'b00000001011010000100;
logic signed [WIDTH-1:0] w_hz_5_7 = 'b11111111000011010010;
logic signed [WIDTH-1:0] w_hz_6_0 = 'b00000000110110111110;
logic signed [WIDTH-1:0] w_hz_6_1 = 'b00000000011100101000;
logic signed [WIDTH-1:0] w_hz_6_2 = 'b11111111101011000100;
logic signed [WIDTH-1:0] w_hz_6_3 = 'b00000000100000100111;
logic signed [WIDTH-1:0] w_hz_6_4 = 'b00000001101000010011;
logic signed [WIDTH-1:0] w_hz_6_5 = 'b11111110011110010001;
logic signed [WIDTH-1:0] w_hz_6_6 = 'b00000000000001101010;
logic signed [WIDTH-1:0] w_hz_6_7 = 'b00000001000111101101;
logic signed [WIDTH-1:0] w_hz_7_0 = 'b00000000110110010110;
logic signed [WIDTH-1:0] w_hz_7_1 = 'b00000000000001010101;
logic signed [WIDTH-1:0] w_hz_7_2 = 'b11111110000010100100;
logic signed [WIDTH-1:0] w_hz_7_3 = 'b00000001110001110110;
logic signed [WIDTH-1:0] w_hz_7_4 = 'b00000001011111101110;
logic signed [WIDTH-1:0] w_hz_7_5 = 'b00000000100010111000;
logic signed [WIDTH-1:0] w_hz_7_6 = 'b11111110110100110001;
logic signed [WIDTH-1:0] w_hz_7_7 = 'b00000010100101110110;

logic signed [WIDTH-1:0] w_hn_0_0 = 'b11111111110101110100;
logic signed [WIDTH-1:0] w_hn_0_1 = 'b11111111101100110010;
logic signed [WIDTH-1:0] w_hn_0_2 = 'b00000000100100011000;
logic signed [WIDTH-1:0] w_hn_0_3 = 'b11111111001100010110;
logic signed [WIDTH-1:0] w_hn_0_4 = 'b11111111010010110100;
logic signed [WIDTH-1:0] w_hn_0_5 = 'b11111111111001110101;
logic signed [WIDTH-1:0] w_hn_0_6 = 'b00000010111011100001;
logic signed [WIDTH-1:0] w_hn_0_7 = 'b11111110100010000101;
logic signed [WIDTH-1:0] w_hn_1_0 = 'b11111111110101110010;
logic signed [WIDTH-1:0] w_hn_1_1 = 'b00000001101100111000;
logic signed [WIDTH-1:0] w_hn_1_2 = 'b00000010011111000111;
logic signed [WIDTH-1:0] w_hn_1_3 = 'b11111110010000010100;
logic signed [WIDTH-1:0] w_hn_1_4 = 'b11111111010110010110;
logic signed [WIDTH-1:0] w_hn_1_5 = 'b11111110110011000110;
logic signed [WIDTH-1:0] w_hn_1_6 = 'b11111111001011100001;
logic signed [WIDTH-1:0] w_hn_1_7 = 'b00000001001110101011;
logic signed [WIDTH-1:0] w_hn_2_0 = 'b00000000000011100100;
logic signed [WIDTH-1:0] w_hn_2_1 = 'b00000000001001101010;
logic signed [WIDTH-1:0] w_hn_2_2 = 'b00000000001111100111;
logic signed [WIDTH-1:0] w_hn_2_3 = 'b11111111010111000111;
logic signed [WIDTH-1:0] w_hn_2_4 = 'b00000001000110000100;
logic signed [WIDTH-1:0] w_hn_2_5 = 'b00000001001011010111;
logic signed [WIDTH-1:0] w_hn_2_6 = 'b00000001001010101110;
logic signed [WIDTH-1:0] w_hn_2_7 = 'b11111110110110001000;
logic signed [WIDTH-1:0] w_hn_3_0 = 'b00000000111111100001;
logic signed [WIDTH-1:0] w_hn_3_1 = 'b00000001000111111010;
logic signed [WIDTH-1:0] w_hn_3_2 = 'b11111111011111011100;
logic signed [WIDTH-1:0] w_hn_3_3 = 'b11111111011000110111;
logic signed [WIDTH-1:0] w_hn_3_4 = 'b00000000011111010000;
logic signed [WIDTH-1:0] w_hn_3_5 = 'b00000000100111111110;
logic signed [WIDTH-1:0] w_hn_3_6 = 'b00000001011010000100;
logic signed [WIDTH-1:0] w_hn_3_7 = 'b11111111000011010010;
logic signed [WIDTH-1:0] w_hn_4_0 = 'b00000000110110111110;
logic signed [WIDTH-1:0] w_hn_4_1 = 'b00000000011100101000;
logic signed [WIDTH-1:0] w_hn_4_2 = 'b11111111101011000100;
logic signed [WIDTH-1:0] w_hn_4_3 = 'b00000000100000100111;
logic signed [WIDTH-1:0] w_hn_4_4 = 'b00000001101000010011;
logic signed [WIDTH-1:0] w_hn_4_5 = 'b11111110011110010001;
logic signed [WIDTH-1:0] w_hn_4_6 = 'b00000000000001101010;
logic signed [WIDTH-1:0] w_hn_4_7 = 'b00000001000111101101;
logic signed [WIDTH-1:0] w_hn_5_0 = 'b00000000110110010110;
logic signed [WIDTH-1:0] w_hn_5_1 = 'b00000000000001010101;
logic signed [WIDTH-1:0] w_hn_5_2 = 'b11111110000010100100;
logic signed [WIDTH-1:0] w_hn_5_3 = 'b00000001110001110110;
logic signed [WIDTH-1:0] w_hn_5_4 = 'b00000001011111101110;
logic signed [WIDTH-1:0] w_hn_5_5 = 'b00000000100010111000;
logic signed [WIDTH-1:0] w_hn_5_6 = 'b11111110110100110001;
logic signed [WIDTH-1:0] w_hn_5_7 = 'b00000010100101110110;
logic signed [WIDTH-1:0] w_hn_6_0 = 'b11111111110101110100;
logic signed [WIDTH-1:0] w_hn_6_1 = 'b11111111101100110010;
logic signed [WIDTH-1:0] w_hn_6_2 = 'b00000000100100011000;
logic signed [WIDTH-1:0] w_hn_6_3 = 'b11111111001100010110;
logic signed [WIDTH-1:0] w_hn_6_4 = 'b11111111010010110100;
logic signed [WIDTH-1:0] w_hn_6_5 = 'b11111111111001110101;
logic signed [WIDTH-1:0] w_hn_6_6 = 'b00000010111011100001;
logic signed [WIDTH-1:0] w_hn_6_7 = 'b11111110100010000101;
logic signed [WIDTH-1:0] w_hn_7_0 = 'b11111111110101110010;
logic signed [WIDTH-1:0] w_hn_7_1 = 'b00000001101100111000;
logic signed [WIDTH-1:0] w_hn_7_2 = 'b00000010011111000111;
logic signed [WIDTH-1:0] w_hn_7_3 = 'b11111110010000010100;
logic signed [WIDTH-1:0] w_hn_7_4 = 'b11111111010110010110;
logic signed [WIDTH-1:0] w_hn_7_5 = 'b11111110110011000110;
logic signed [WIDTH-1:0] w_hn_7_6 = 'b11111111001011100001;
logic signed [WIDTH-1:0] w_hn_7_7 = 'b00000001001110101011;

// Biases (h for each gate type)
logic signed [WIDTH-1:0] b_ir_0 = 'b00000000000101110001;
logic signed [WIDTH-1:0] b_ir_1 = 'b00000001000010101100;
logic signed [WIDTH-1:0] b_ir_2 = 'b00000001110110110001;
logic signed [WIDTH-1:0] b_ir_3 = 'b00000000101000110101;
logic signed [WIDTH-1:0] b_ir_4 = 'b00000000110000100110;
logic signed [WIDTH-1:0] b_ir_5 = 'b00000000100010010111;
logic signed [WIDTH-1:0] b_ir_6 = 'b00000001111110001000;
logic signed [WIDTH-1:0] b_ir_7 = 'b11111111111101000000;

logic signed [WIDTH-1:0] b_iz_0 = 'b00000001010101000011;
logic signed [WIDTH-1:0] b_iz_1 = 'b00000000001110100001;
logic signed [WIDTH-1:0] b_iz_2 = 'b00000001110000100001;
logic signed [WIDTH-1:0] b_iz_3 = 'b00000000010011000011;
logic signed [WIDTH-1:0] b_iz_4 = 'b00000000010010010011;
logic signed [WIDTH-1:0] b_iz_5 = 'b00000001001110001101;
logic signed [WIDTH-1:0] b_iz_6 = 'b00000000110111000001;
logic signed [WIDTH-1:0] b_iz_7 = 'b00000001101000110100;

logic signed [WIDTH-1:0] b_in_0 = 'b00000000110100010010;
logic signed [WIDTH-1:0] b_in_1 = 'b00000001001001001100;
logic signed [WIDTH-1:0] b_in_2 = 'b00000000100111111010;
logic signed [WIDTH-1:0] b_in_3 = 'b00000011001110110011;
logic signed [WIDTH-1:0] b_in_4 = 'b00000000011000010011;
logic signed [WIDTH-1:0] b_in_5 = 'b00000010010111111001;
logic signed [WIDTH-1:0] b_in_6 = 'b00000000111010100000;
logic signed [WIDTH-1:0] b_in_7 = 'b11111110000100001001;

logic signed [WIDTH-1:0] b_hr_0 = 'b00000000000101110001;
logic signed [WIDTH-1:0] b_hr_1 = 'b00000001000010101100;
logic signed [WIDTH-1:0] b_hr_2 = 'b00000001110110110001;
logic signed [WIDTH-1:0] b_hr_3 = 'b00000000101000110101;
logic signed [WIDTH-1:0] b_hr_4 = 'b00000000110000100110;
logic signed [WIDTH-1:0] b_hr_5 = 'b00000000100010010111;
logic signed [WIDTH-1:0] b_hr_6 = 'b00000001111110001000;
logic signed [WIDTH-1:0] b_hr_7 = 'b11111111111101000000;

logic signed [WIDTH-1:0] b_hz_0 = 'b00000001010101000011;
logic signed [WIDTH-1:0] b_hz_1 = 'b00000000001110100001;
logic signed [WIDTH-1:0] b_hz_2 = 'b00000001110000100001;
logic signed [WIDTH-1:0] b_hz_3 = 'b00000000010011000011;
logic signed [WIDTH-1:0] b_hz_4 = 'b00000000010010010011;
logic signed [WIDTH-1:0] b_hz_5 = 'b00000001001110001101;
logic signed [WIDTH-1:0] b_hz_6 = 'b00000000110111000001;
logic signed [WIDTH-1:0] b_hz_7 = 'b00000001101000110100;

logic signed [WIDTH-1:0] b_hn_0 = 'b00000000110100010010;
logic signed [WIDTH-1:0] b_hn_1 = 'b00000001001001001100;
logic signed [WIDTH-1:0] b_hn_2 = 'b00000000100111111010;
logic signed [WIDTH-1:0] b_hn_3 = 'b00000011001110110011;
logic signed [WIDTH-1:0] b_hn_4 = 'b00000000011000010011;
logic signed [WIDTH-1:0] b_hn_5 = 'b00000010010111111001;
logic signed [WIDTH-1:0] b_hn_6 = 'b00000000111010100000;
logic signed [WIDTH-1:0] b_hn_7 = 'b11111110000100001001;

// Outputs (h=8)
logic signed [WIDTH-1:0]  y_0 = 0;
logic signed [WIDTH-1:0]  y_1 = 0;
logic signed [WIDTH-1:0]  y_2 = 0;
logic signed [WIDTH-1:0]  y_3 = 0;
logic signed [WIDTH-1:0]  y_4 = 0;
logic signed [WIDTH-1:0]  y_5 = 0;
logic signed [WIDTH-1:0]  y_6 = 0;
logic signed [WIDTH-1:0]  y_7 = 0;

gru #(
        .INT_WIDTH(INT_WIDTH),
        .FRAC_WIDTH(FRAC_WIDTH)
    ) gru_inst (
        .clk(clk),
        .reset(reset),
        // Input features (d=64)
        	
.x_0(x_0), .x_1(x_1), .x_2(x_2), .x_3(x_3), .x_4(x_4), .x_5(x_5), .x_6(x_6), .x_7(x_7), .x_8(x_8), .x_9(x_9), .x_10(x_10), .x_11(x_11), .x_12(x_12), .x_13(x_13), .x_14(x_14), .x_15(x_15), 	
.h_0(h_0), .h_1(h_1), .h_2(h_2), .h_3(h_3), .h_4(h_4), .h_5(h_5), .h_6(h_6), .h_7(h_7), 	
.w_ir_0_0(w_ir_0_0), .w_ir_0_1(w_ir_0_1), .w_ir_0_2(w_ir_0_2), .w_ir_0_3(w_ir_0_3), .w_ir_0_4(w_ir_0_4), .w_ir_0_5(w_ir_0_5), .w_ir_0_6(w_ir_0_6), .w_ir_0_7(w_ir_0_7), .w_ir_0_8(w_ir_0_8), .w_ir_0_9(w_ir_0_9), .w_ir_0_10(w_ir_0_10), .w_ir_0_11(w_ir_0_11), .w_ir_0_12(w_ir_0_12), .w_ir_0_13(w_ir_0_13), .w_ir_0_14(w_ir_0_14), .w_ir_0_15(w_ir_0_15), .w_ir_1_0(w_ir_1_0), .w_ir_1_1(w_ir_1_1), .w_ir_1_2(w_ir_1_2), .w_ir_1_3(w_ir_1_3), .w_ir_1_4(w_ir_1_4), .w_ir_1_5(w_ir_1_5), .w_ir_1_6(w_ir_1_6), .w_ir_1_7(w_ir_1_7), .w_ir_1_8(w_ir_1_8), .w_ir_1_9(w_ir_1_9), .w_ir_1_10(w_ir_1_10), .w_ir_1_11(w_ir_1_11), .w_ir_1_12(w_ir_1_12), .w_ir_1_13(w_ir_1_13), .w_ir_1_14(w_ir_1_14), .w_ir_1_15(w_ir_1_15), .w_ir_2_0(w_ir_2_0), .w_ir_2_1(w_ir_2_1), .w_ir_2_2(w_ir_2_2), .w_ir_2_3(w_ir_2_3), .w_ir_2_4(w_ir_2_4), .w_ir_2_5(w_ir_2_5), .w_ir_2_6(w_ir_2_6), .w_ir_2_7(w_ir_2_7), .w_ir_2_8(w_ir_2_8), .w_ir_2_9(w_ir_2_9), .w_ir_2_10(w_ir_2_10), .w_ir_2_11(w_ir_2_11), .w_ir_2_12(w_ir_2_12), .w_ir_2_13(w_ir_2_13), .w_ir_2_14(w_ir_2_14), .w_ir_2_15(w_ir_2_15), .w_ir_3_0(w_ir_3_0), .w_ir_3_1(w_ir_3_1), .w_ir_3_2(w_ir_3_2), .w_ir_3_3(w_ir_3_3), .w_ir_3_4(w_ir_3_4), .w_ir_3_5(w_ir_3_5), .w_ir_3_6(w_ir_3_6), .w_ir_3_7(w_ir_3_7), .w_ir_3_8(w_ir_3_8), .w_ir_3_9(w_ir_3_9), .w_ir_3_10(w_ir_3_10), .w_ir_3_11(w_ir_3_11), .w_ir_3_12(w_ir_3_12), .w_ir_3_13(w_ir_3_13), .w_ir_3_14(w_ir_3_14), .w_ir_3_15(w_ir_3_15), .w_ir_4_0(w_ir_4_0), .w_ir_4_1(w_ir_4_1), .w_ir_4_2(w_ir_4_2), .w_ir_4_3(w_ir_4_3), .w_ir_4_4(w_ir_4_4), .w_ir_4_5(w_ir_4_5), .w_ir_4_6(w_ir_4_6), .w_ir_4_7(w_ir_4_7), .w_ir_4_8(w_ir_4_8), .w_ir_4_9(w_ir_4_9), .w_ir_4_10(w_ir_4_10), .w_ir_4_11(w_ir_4_11), .w_ir_4_12(w_ir_4_12), .w_ir_4_13(w_ir_4_13), .w_ir_4_14(w_ir_4_14), .w_ir_4_15(w_ir_4_15), .w_ir_5_0(w_ir_5_0), .w_ir_5_1(w_ir_5_1), .w_ir_5_2(w_ir_5_2), .w_ir_5_3(w_ir_5_3), .w_ir_5_4(w_ir_5_4), .w_ir_5_5(w_ir_5_5), .w_ir_5_6(w_ir_5_6), .w_ir_5_7(w_ir_5_7), .w_ir_5_8(w_ir_5_8), .w_ir_5_9(w_ir_5_9), .w_ir_5_10(w_ir_5_10), .w_ir_5_11(w_ir_5_11), .w_ir_5_12(w_ir_5_12), .w_ir_5_13(w_ir_5_13), .w_ir_5_14(w_ir_5_14), .w_ir_5_15(w_ir_5_15), .w_ir_6_0(w_ir_6_0), .w_ir_6_1(w_ir_6_1), .w_ir_6_2(w_ir_6_2), .w_ir_6_3(w_ir_6_3), .w_ir_6_4(w_ir_6_4), .w_ir_6_5(w_ir_6_5), .w_ir_6_6(w_ir_6_6), .w_ir_6_7(w_ir_6_7), .w_ir_6_8(w_ir_6_8), .w_ir_6_9(w_ir_6_9), .w_ir_6_10(w_ir_6_10), .w_ir_6_11(w_ir_6_11), .w_ir_6_12(w_ir_6_12), .w_ir_6_13(w_ir_6_13), .w_ir_6_14(w_ir_6_14), .w_ir_6_15(w_ir_6_15), .w_ir_7_0(w_ir_7_0), .w_ir_7_1(w_ir_7_1), .w_ir_7_2(w_ir_7_2), .w_ir_7_3(w_ir_7_3), .w_ir_7_4(w_ir_7_4), .w_ir_7_5(w_ir_7_5), .w_ir_7_6(w_ir_7_6), .w_ir_7_7(w_ir_7_7), .w_ir_7_8(w_ir_7_8), .w_ir_7_9(w_ir_7_9), .w_ir_7_10(w_ir_7_10), .w_ir_7_11(w_ir_7_11), .w_ir_7_12(w_ir_7_12), .w_ir_7_13(w_ir_7_13), .w_ir_7_14(w_ir_7_14), .w_ir_7_15(w_ir_7_15), 	
.w_iz_0_0(w_iz_0_0), .w_iz_0_1(w_iz_0_1), .w_iz_0_2(w_iz_0_2), .w_iz_0_3(w_iz_0_3), .w_iz_0_4(w_iz_0_4), .w_iz_0_5(w_iz_0_5), .w_iz_0_6(w_iz_0_6), .w_iz_0_7(w_iz_0_7), .w_iz_0_8(w_iz_0_8), .w_iz_0_9(w_iz_0_9), .w_iz_0_10(w_iz_0_10), .w_iz_0_11(w_iz_0_11), .w_iz_0_12(w_iz_0_12), .w_iz_0_13(w_iz_0_13), .w_iz_0_14(w_iz_0_14), .w_iz_0_15(w_iz_0_15), .w_iz_1_0(w_iz_1_0), .w_iz_1_1(w_iz_1_1), .w_iz_1_2(w_iz_1_2), .w_iz_1_3(w_iz_1_3), .w_iz_1_4(w_iz_1_4), .w_iz_1_5(w_iz_1_5), .w_iz_1_6(w_iz_1_6), .w_iz_1_7(w_iz_1_7), .w_iz_1_8(w_iz_1_8), .w_iz_1_9(w_iz_1_9), .w_iz_1_10(w_iz_1_10), .w_iz_1_11(w_iz_1_11), .w_iz_1_12(w_iz_1_12), .w_iz_1_13(w_iz_1_13), .w_iz_1_14(w_iz_1_14), .w_iz_1_15(w_iz_1_15), .w_iz_2_0(w_iz_2_0), .w_iz_2_1(w_iz_2_1), .w_iz_2_2(w_iz_2_2), .w_iz_2_3(w_iz_2_3), .w_iz_2_4(w_iz_2_4), .w_iz_2_5(w_iz_2_5), .w_iz_2_6(w_iz_2_6), .w_iz_2_7(w_iz_2_7), .w_iz_2_8(w_iz_2_8), .w_iz_2_9(w_iz_2_9), .w_iz_2_10(w_iz_2_10), .w_iz_2_11(w_iz_2_11), .w_iz_2_12(w_iz_2_12), .w_iz_2_13(w_iz_2_13), .w_iz_2_14(w_iz_2_14), .w_iz_2_15(w_iz_2_15), .w_iz_3_0(w_iz_3_0), .w_iz_3_1(w_iz_3_1), .w_iz_3_2(w_iz_3_2), .w_iz_3_3(w_iz_3_3), .w_iz_3_4(w_iz_3_4), .w_iz_3_5(w_iz_3_5), .w_iz_3_6(w_iz_3_6), .w_iz_3_7(w_iz_3_7), .w_iz_3_8(w_iz_3_8), .w_iz_3_9(w_iz_3_9), .w_iz_3_10(w_iz_3_10), .w_iz_3_11(w_iz_3_11), .w_iz_3_12(w_iz_3_12), .w_iz_3_13(w_iz_3_13), .w_iz_3_14(w_iz_3_14), .w_iz_3_15(w_iz_3_15), .w_iz_4_0(w_iz_4_0), .w_iz_4_1(w_iz_4_1), .w_iz_4_2(w_iz_4_2), .w_iz_4_3(w_iz_4_3), .w_iz_4_4(w_iz_4_4), .w_iz_4_5(w_iz_4_5), .w_iz_4_6(w_iz_4_6), .w_iz_4_7(w_iz_4_7), .w_iz_4_8(w_iz_4_8), .w_iz_4_9(w_iz_4_9), .w_iz_4_10(w_iz_4_10), .w_iz_4_11(w_iz_4_11), .w_iz_4_12(w_iz_4_12), .w_iz_4_13(w_iz_4_13), .w_iz_4_14(w_iz_4_14), .w_iz_4_15(w_iz_4_15), .w_iz_5_0(w_iz_5_0), .w_iz_5_1(w_iz_5_1), .w_iz_5_2(w_iz_5_2), .w_iz_5_3(w_iz_5_3), .w_iz_5_4(w_iz_5_4), .w_iz_5_5(w_iz_5_5), .w_iz_5_6(w_iz_5_6), .w_iz_5_7(w_iz_5_7), .w_iz_5_8(w_iz_5_8), .w_iz_5_9(w_iz_5_9), .w_iz_5_10(w_iz_5_10), .w_iz_5_11(w_iz_5_11), .w_iz_5_12(w_iz_5_12), .w_iz_5_13(w_iz_5_13), .w_iz_5_14(w_iz_5_14), .w_iz_5_15(w_iz_5_15), .w_iz_6_0(w_iz_6_0), .w_iz_6_1(w_iz_6_1), .w_iz_6_2(w_iz_6_2), .w_iz_6_3(w_iz_6_3), .w_iz_6_4(w_iz_6_4), .w_iz_6_5(w_iz_6_5), .w_iz_6_6(w_iz_6_6), .w_iz_6_7(w_iz_6_7), .w_iz_6_8(w_iz_6_8), .w_iz_6_9(w_iz_6_9), .w_iz_6_10(w_iz_6_10), .w_iz_6_11(w_iz_6_11), .w_iz_6_12(w_iz_6_12), .w_iz_6_13(w_iz_6_13), .w_iz_6_14(w_iz_6_14), .w_iz_6_15(w_iz_6_15), .w_iz_7_0(w_iz_7_0), .w_iz_7_1(w_iz_7_1), .w_iz_7_2(w_iz_7_2), .w_iz_7_3(w_iz_7_3), .w_iz_7_4(w_iz_7_4), .w_iz_7_5(w_iz_7_5), .w_iz_7_6(w_iz_7_6), .w_iz_7_7(w_iz_7_7), .w_iz_7_8(w_iz_7_8), .w_iz_7_9(w_iz_7_9), .w_iz_7_10(w_iz_7_10), .w_iz_7_11(w_iz_7_11), .w_iz_7_12(w_iz_7_12), .w_iz_7_13(w_iz_7_13), .w_iz_7_14(w_iz_7_14), .w_iz_7_15(w_iz_7_15), 
.w_in_0_0(w_in_0_0), .w_in_0_1(w_in_0_1), .w_in_0_2(w_in_0_2), .w_in_0_3(w_in_0_3), .w_in_0_4(w_in_0_4), .w_in_0_5(w_in_0_5), .w_in_0_6(w_in_0_6), .w_in_0_7(w_in_0_7), .w_in_0_8(w_in_0_8), .w_in_0_9(w_in_0_9), .w_in_0_10(w_in_0_10), .w_in_0_11(w_in_0_11), .w_in_0_12(w_in_0_12), .w_in_0_13(w_in_0_13), .w_in_0_14(w_in_0_14), .w_in_0_15(w_in_0_15), .w_in_1_0(w_in_1_0), .w_in_1_1(w_in_1_1), .w_in_1_2(w_in_1_2), .w_in_1_3(w_in_1_3), .w_in_1_4(w_in_1_4), .w_in_1_5(w_in_1_5), .w_in_1_6(w_in_1_6), .w_in_1_7(w_in_1_7), .w_in_1_8(w_in_1_8), .w_in_1_9(w_in_1_9), .w_in_1_10(w_in_1_10), .w_in_1_11(w_in_1_11), .w_in_1_12(w_in_1_12), .w_in_1_13(w_in_1_13), .w_in_1_14(w_in_1_14), .w_in_1_15(w_in_1_15), .w_in_2_0(w_in_2_0), .w_in_2_1(w_in_2_1), .w_in_2_2(w_in_2_2), .w_in_2_3(w_in_2_3), .w_in_2_4(w_in_2_4), .w_in_2_5(w_in_2_5), .w_in_2_6(w_in_2_6), .w_in_2_7(w_in_2_7), .w_in_2_8(w_in_2_8), .w_in_2_9(w_in_2_9), .w_in_2_10(w_in_2_10), .w_in_2_11(w_in_2_11), .w_in_2_12(w_in_2_12), .w_in_2_13(w_in_2_13), .w_in_2_14(w_in_2_14), .w_in_2_15(w_in_2_15), .w_in_3_0(w_in_3_0), .w_in_3_1(w_in_3_1), .w_in_3_2(w_in_3_2), .w_in_3_3(w_in_3_3), .w_in_3_4(w_in_3_4), .w_in_3_5(w_in_3_5), .w_in_3_6(w_in_3_6), .w_in_3_7(w_in_3_7), .w_in_3_8(w_in_3_8), .w_in_3_9(w_in_3_9), .w_in_3_10(w_in_3_10), .w_in_3_11(w_in_3_11), .w_in_3_12(w_in_3_12), .w_in_3_13(w_in_3_13), .w_in_3_14(w_in_3_14), .w_in_3_15(w_in_3_15), .w_in_4_0(w_in_4_0), .w_in_4_1(w_in_4_1), .w_in_4_2(w_in_4_2), .w_in_4_3(w_in_4_3), .w_in_4_4(w_in_4_4), .w_in_4_5(w_in_4_5), .w_in_4_6(w_in_4_6), .w_in_4_7(w_in_4_7), .w_in_4_8(w_in_4_8), .w_in_4_9(w_in_4_9), .w_in_4_10(w_in_4_10), .w_in_4_11(w_in_4_11), .w_in_4_12(w_in_4_12), .w_in_4_13(w_in_4_13), .w_in_4_14(w_in_4_14), .w_in_4_15(w_in_4_15), .w_in_5_0(w_in_5_0), .w_in_5_1(w_in_5_1), .w_in_5_2(w_in_5_2), .w_in_5_3(w_in_5_3), .w_in_5_4(w_in_5_4), .w_in_5_5(w_in_5_5), .w_in_5_6(w_in_5_6), .w_in_5_7(w_in_5_7), .w_in_5_8(w_in_5_8), .w_in_5_9(w_in_5_9), .w_in_5_10(w_in_5_10), .w_in_5_11(w_in_5_11), .w_in_5_12(w_in_5_12), .w_in_5_13(w_in_5_13), .w_in_5_14(w_in_5_14), .w_in_5_15(w_in_5_15), .w_in_6_0(w_in_6_0), .w_in_6_1(w_in_6_1), .w_in_6_2(w_in_6_2), .w_in_6_3(w_in_6_3), .w_in_6_4(w_in_6_4), .w_in_6_5(w_in_6_5), .w_in_6_6(w_in_6_6), .w_in_6_7(w_in_6_7), .w_in_6_8(w_in_6_8), .w_in_6_9(w_in_6_9), .w_in_6_10(w_in_6_10), .w_in_6_11(w_in_6_11), .w_in_6_12(w_in_6_12), .w_in_6_13(w_in_6_13), .w_in_6_14(w_in_6_14), .w_in_6_15(w_in_6_15), .w_in_7_0(w_in_7_0), .w_in_7_1(w_in_7_1), .w_in_7_2(w_in_7_2), .w_in_7_3(w_in_7_3), .w_in_7_4(w_in_7_4), .w_in_7_5(w_in_7_5), .w_in_7_6(w_in_7_6), .w_in_7_7(w_in_7_7), .w_in_7_8(w_in_7_8), .w_in_7_9(w_in_7_9), .w_in_7_10(w_in_7_10), .w_in_7_11(w_in_7_11), .w_in_7_12(w_in_7_12), .w_in_7_13(w_in_7_13), .w_in_7_14(w_in_7_14), .w_in_7_15(w_in_7_15), 
.w_hr_0_0(w_hr_0_0), .w_hr_0_1(w_hr_0_1), .w_hr_0_2(w_hr_0_2), .w_hr_0_3(w_hr_0_3), .w_hr_0_4(w_hr_0_4), .w_hr_0_5(w_hr_0_5), .w_hr_0_6(w_hr_0_6), .w_hr_0_7(w_hr_0_7), .w_hr_1_0(w_hr_1_0), .w_hr_1_1(w_hr_1_1), .w_hr_1_2(w_hr_1_2), .w_hr_1_3(w_hr_1_3), .w_hr_1_4(w_hr_1_4), .w_hr_1_5(w_hr_1_5), .w_hr_1_6(w_hr_1_6), .w_hr_1_7(w_hr_1_7), .w_hr_2_0(w_hr_2_0), .w_hr_2_1(w_hr_2_1), .w_hr_2_2(w_hr_2_2), .w_hr_2_3(w_hr_2_3), .w_hr_2_4(w_hr_2_4), .w_hr_2_5(w_hr_2_5), .w_hr_2_6(w_hr_2_6), .w_hr_2_7(w_hr_2_7), .w_hr_3_0(w_hr_3_0), .w_hr_3_1(w_hr_3_1), .w_hr_3_2(w_hr_3_2), .w_hr_3_3(w_hr_3_3), .w_hr_3_4(w_hr_3_4), .w_hr_3_5(w_hr_3_5), .w_hr_3_6(w_hr_3_6), .w_hr_3_7(w_hr_3_7), .w_hr_4_0(w_hr_4_0), .w_hr_4_1(w_hr_4_1), .w_hr_4_2(w_hr_4_2), .w_hr_4_3(w_hr_4_3), .w_hr_4_4(w_hr_4_4), .w_hr_4_5(w_hr_4_5), .w_hr_4_6(w_hr_4_6), .w_hr_4_7(w_hr_4_7), .w_hr_5_0(w_hr_5_0), .w_hr_5_1(w_hr_5_1), .w_hr_5_2(w_hr_5_2), .w_hr_5_3(w_hr_5_3), .w_hr_5_4(w_hr_5_4), .w_hr_5_5(w_hr_5_5), .w_hr_5_6(w_hr_5_6), .w_hr_5_7(w_hr_5_7), .w_hr_6_0(w_hr_6_0), .w_hr_6_1(w_hr_6_1), .w_hr_6_2(w_hr_6_2), .w_hr_6_3(w_hr_6_3), .w_hr_6_4(w_hr_6_4), .w_hr_6_5(w_hr_6_5), .w_hr_6_6(w_hr_6_6), .w_hr_6_7(w_hr_6_7), .w_hr_7_0(w_hr_7_0), .w_hr_7_1(w_hr_7_1), .w_hr_7_2(w_hr_7_2), .w_hr_7_3(w_hr_7_3), .w_hr_7_4(w_hr_7_4), .w_hr_7_5(w_hr_7_5), .w_hr_7_6(w_hr_7_6), .w_hr_7_7(w_hr_7_7), 
.w_hz_0_0(w_hz_0_0), .w_hz_0_1(w_hz_0_1), .w_hz_0_2(w_hz_0_2), .w_hz_0_3(w_hz_0_3), .w_hz_0_4(w_hz_0_4), .w_hz_0_5(w_hz_0_5), .w_hz_0_6(w_hz_0_6), .w_hz_0_7(w_hz_0_7), .w_hz_1_0(w_hz_1_0), .w_hz_1_1(w_hz_1_1), .w_hz_1_2(w_hz_1_2), .w_hz_1_3(w_hz_1_3), .w_hz_1_4(w_hz_1_4), .w_hz_1_5(w_hz_1_5), .w_hz_1_6(w_hz_1_6), .w_hz_1_7(w_hz_1_7), .w_hz_2_0(w_hz_2_0), .w_hz_2_1(w_hz_2_1), .w_hz_2_2(w_hz_2_2), .w_hz_2_3(w_hz_2_3), .w_hz_2_4(w_hz_2_4), .w_hz_2_5(w_hz_2_5), .w_hz_2_6(w_hz_2_6), .w_hz_2_7(w_hz_2_7), .w_hz_3_0(w_hz_3_0), .w_hz_3_1(w_hz_3_1), .w_hz_3_2(w_hz_3_2), .w_hz_3_3(w_hz_3_3), .w_hz_3_4(w_hz_3_4), .w_hz_3_5(w_hz_3_5), .w_hz_3_6(w_hz_3_6), .w_hz_3_7(w_hz_3_7), .w_hz_4_0(w_hz_4_0), .w_hz_4_1(w_hz_4_1), .w_hz_4_2(w_hz_4_2), .w_hz_4_3(w_hz_4_3), .w_hz_4_4(w_hz_4_4), .w_hz_4_5(w_hz_4_5), .w_hz_4_6(w_hz_4_6), .w_hz_4_7(w_hz_4_7), .w_hz_5_0(w_hz_5_0), .w_hz_5_1(w_hz_5_1), .w_hz_5_2(w_hz_5_2), .w_hz_5_3(w_hz_5_3), .w_hz_5_4(w_hz_5_4), .w_hz_5_5(w_hz_5_5), .w_hz_5_6(w_hz_5_6), .w_hz_5_7(w_hz_5_7), .w_hz_6_0(w_hz_6_0), .w_hz_6_1(w_hz_6_1), .w_hz_6_2(w_hz_6_2), .w_hz_6_3(w_hz_6_3), .w_hz_6_4(w_hz_6_4), .w_hz_6_5(w_hz_6_5), .w_hz_6_6(w_hz_6_6), .w_hz_6_7(w_hz_6_7), .w_hz_7_0(w_hz_7_0), .w_hz_7_1(w_hz_7_1), .w_hz_7_2(w_hz_7_2), .w_hz_7_3(w_hz_7_3), .w_hz_7_4(w_hz_7_4), .w_hz_7_5(w_hz_7_5), .w_hz_7_6(w_hz_7_6), .w_hz_7_7(w_hz_7_7), 
.w_hn_0_0(w_hn_0_0), .w_hn_0_1(w_hn_0_1), .w_hn_0_2(w_hn_0_2), .w_hn_0_3(w_hn_0_3), .w_hn_0_4(w_hn_0_4), .w_hn_0_5(w_hn_0_5), .w_hn_0_6(w_hn_0_6), .w_hn_0_7(w_hn_0_7), .w_hn_1_0(w_hn_1_0), .w_hn_1_1(w_hn_1_1), .w_hn_1_2(w_hn_1_2), .w_hn_1_3(w_hn_1_3), .w_hn_1_4(w_hn_1_4), .w_hn_1_5(w_hn_1_5), .w_hn_1_6(w_hn_1_6), .w_hn_1_7(w_hn_1_7), .w_hn_2_0(w_hn_2_0), .w_hn_2_1(w_hn_2_1), .w_hn_2_2(w_hn_2_2), .w_hn_2_3(w_hn_2_3), .w_hn_2_4(w_hn_2_4), .w_hn_2_5(w_hn_2_5), .w_hn_2_6(w_hn_2_6), .w_hn_2_7(w_hn_2_7), .w_hn_3_0(w_hn_3_0), .w_hn_3_1(w_hn_3_1), .w_hn_3_2(w_hn_3_2), .w_hn_3_3(w_hn_3_3), .w_hn_3_4(w_hn_3_4), .w_hn_3_5(w_hn_3_5), .w_hn_3_6(w_hn_3_6), .w_hn_3_7(w_hn_3_7), .w_hn_4_0(w_hn_4_0), .w_hn_4_1(w_hn_4_1), .w_hn_4_2(w_hn_4_2), .w_hn_4_3(w_hn_4_3), .w_hn_4_4(w_hn_4_4), .w_hn_4_5(w_hn_4_5), .w_hn_4_6(w_hn_4_6), .w_hn_4_7(w_hn_4_7), .w_hn_5_0(w_hn_5_0), .w_hn_5_1(w_hn_5_1), .w_hn_5_2(w_hn_5_2), .w_hn_5_3(w_hn_5_3), .w_hn_5_4(w_hn_5_4), .w_hn_5_5(w_hn_5_5), .w_hn_5_6(w_hn_5_6), .w_hn_5_7(w_hn_5_7), .w_hn_6_0(w_hn_6_0), .w_hn_6_1(w_hn_6_1), .w_hn_6_2(w_hn_6_2), .w_hn_6_3(w_hn_6_3), .w_hn_6_4(w_hn_6_4), .w_hn_6_5(w_hn_6_5), .w_hn_6_6(w_hn_6_6), .w_hn_6_7(w_hn_6_7), .w_hn_7_0(w_hn_7_0), .w_hn_7_1(w_hn_7_1), .w_hn_7_2(w_hn_7_2), .w_hn_7_3(w_hn_7_3), .w_hn_7_4(w_hn_7_4), .w_hn_7_5(w_hn_7_5), .w_hn_7_6(w_hn_7_6), .w_hn_7_7(w_hn_7_7), 
.b_ir_0(b_ir_0), .b_ir_1(b_ir_1), .b_ir_2(b_ir_2), .b_ir_3(b_ir_3), .b_ir_4(b_ir_4), .b_ir_5(b_ir_5), .b_ir_6(b_ir_6), .b_ir_7(b_ir_7), 
.b_iz_0(b_iz_0), .b_iz_1(b_iz_1), .b_iz_2(b_iz_2), .b_iz_3(b_iz_3), .b_iz_4(b_iz_4), .b_iz_5(b_iz_5), .b_iz_6(b_iz_6), .b_iz_7(b_iz_7), 
.b_in_0(b_in_0), .b_in_1(b_in_1), .b_in_2(b_in_2), .b_in_3(b_in_3), .b_in_4(b_in_4), .b_in_5(b_in_5), .b_in_6(b_in_6), .b_in_7(b_in_7), 
.b_hr_0(b_hr_0), .b_hr_1(b_hr_1), .b_hr_2(b_hr_2), .b_hr_3(b_hr_3), .b_hr_4(b_hr_4), .b_hr_5(b_hr_5), .b_hr_6(b_hr_6), .b_hr_7(b_hr_7), 
.b_hz_0(b_hz_0), .b_hz_1(b_hz_1), .b_hz_2(b_hz_2), .b_hz_3(b_hz_3), .b_hz_4(b_hz_4), .b_hz_5(b_hz_5), .b_hz_6(b_hz_6), .b_hz_7(b_hz_7), 
.b_hn_0(b_hn_0), .b_hn_1(b_hn_1), .b_hn_2(b_hn_2), .b_hn_3(b_hn_3), .b_hn_4(b_hn_4), .b_hn_5(b_hn_5), .b_hn_6(b_hn_6), .b_hn_7(b_hn_7), 
.y_0(y_0), .y_1(y_1), .y_2(y_2), .y_3(y_3), .y_4(y_4), .y_5(y_5), .y_6(y_6), .y_7(y_7)
);

    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end
    
    initial begin
        // Open file for writing (overwrite existing)
        integer fd;
        fd = $fopen("../../../../../output_d16_h8_int6_frac14.txt", "w+");
        if (fd == 0) begin
            $display("ERROR: Failed to open file!");
            $finish;
        end
        x_0 = 'b00000100100010010100;
    x_1 = 'b00000110110110001001;
    x_2 = 'b00001000001001001101;
    x_3 = 'b00001001000110011110;
    x_4 = 'b00000111010100111000;
    x_5 = 'b00000110101110000100;
    x_6 = 'b00000100111010001100;
    x_7 = 'b00000100100111110001;
    x_8 = 'b00000111100001010001;
    x_9 = 'b00001001000010001000;
    x_10 = 'b00001001011010010111;
    x_11 = 'b00001001001001001011;
    x_12 = 'b00001000111011000001;
    x_13 = 'b00000101100100011010;
    x_14 = 'b00000111010101110111;
    x_15 = 'b00001000110010000011;

    h_0 = 'b00000100100010010100;
    h_1 = 'b00000110110110001001;
    h_2 = 'b00001000001001001101;
    h_3 = 'b00001001000110011110;
    h_4 = 'b00000111010100111000;
    h_5 = 'b00000110101110000100;
    h_6 = 'b00000100111010001100;
    h_7 = 'b00000100100111110001;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000101110001001111;
    x_1 = 'b00001001001000111110;
    x_2 = 'b00001010001100010100;
    x_3 = 'b00001010101011111111;
    x_4 = 'b00001001111011100110;
    x_5 = 'b00001001011111100101;
    x_6 = 'b00000111111011000111;
    x_7 = 'b00000110110110010001;
    x_8 = 'b00001010001011011101;
    x_9 = 'b00001011001110011100;
    x_10 = 'b00001011010100101010;
    x_11 = 'b00001011110110011100;
    x_12 = 'b00001011010011001100;
    x_13 = 'b00001000000001001001;
    x_14 = 'b00001001101001100001;
    x_15 = 'b00001010110110010001;

    h_0 = 'b00000101110001001111;
    h_1 = 'b00001001001000111110;
    h_2 = 'b00001010001100010100;
    h_3 = 'b00001010101011111111;
    h_4 = 'b00001001111011100110;
    h_5 = 'b00001001011111100101;
    h_6 = 'b00000111111011000111;
    h_7 = 'b00000110110110010001;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000111111011010110;
    x_1 = 'b00001000011000000010;
    x_2 = 'b00001000000100010111;
    x_3 = 'b00000111111101111101;
    x_4 = 'b00000110110110100100;
    x_5 = 'b00000101100101111101;
    x_6 = 'b00000011101111100000;
    x_7 = 'b00000110001101100011;
    x_8 = 'b00001000001111101011;
    x_9 = 'b00001000001011000000;
    x_10 = 'b00001000000010010010;
    x_11 = 'b00001000011011010100;
    x_12 = 'b00000110100010110101;
    x_13 = 'b00000001101111000110;
    x_14 = 'b00001000000101010101;
    x_15 = 'b00001000010011100010;

    h_0 = 'b00000111111011010110;
    h_1 = 'b00001000011000000010;
    h_2 = 'b00001000000100010111;
    h_3 = 'b00000111111101111101;
    h_4 = 'b00000110110110100100;
    h_5 = 'b00000101100101111101;
    h_6 = 'b00000011101111100000;
    h_7 = 'b00000110001101100011;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000101100111010111;
    x_1 = 'b00000101111011011010;
    x_2 = 'b00000110100011001111;
    x_3 = 'b00000111001101100111;
    x_4 = 'b00000110000100000011;
    x_5 = 'b00000100100011011001;
    x_6 = 'b00000011011100110101;
    x_7 = 'b00000011110100110111;
    x_8 = 'b00000110000100011011;
    x_9 = 'b00000110101011110010;
    x_10 = 'b00000110111101110011;
    x_11 = 'b00000111011110001010;
    x_12 = 'b00000101010110101111;
    x_13 = 'b00000010001010010110;
    x_14 = 'b00000101110001101011;
    x_15 = 'b00000110101101110100;

    h_0 = 'b00000101100111010111;
    h_1 = 'b00000101111011011010;
    h_2 = 'b00000110100011001111;
    h_3 = 'b00000111001101100111;
    h_4 = 'b00000110000100000011;
    h_5 = 'b00000100100011011001;
    h_6 = 'b00000011011100110101;
    h_7 = 'b00000011110100110111;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000011100010001100;
    x_1 = 'b00000100101101000110;
    x_2 = 'b00000101001011110101;
    x_3 = 'b00000110001001111100;
    x_4 = 'b00000101100000101011;
    x_5 = 'b00000100000010000111;
    x_6 = 'b00000011101001010010;
    x_7 = 'b00000010100011011011;
    x_8 = 'b00000100001000101010;
    x_9 = 'b00000100111000100010;
    x_10 = 'b00000101010010001010;
    x_11 = 'b00000110000010011100;
    x_12 = 'b00000100000100110011;
    x_13 = 'b00000001111100101110;
    x_14 = 'b00000100010010110000;
    x_15 = 'b00000101000011000010;

    h_0 = 'b00000011100010001100;
    h_1 = 'b00000100101101000110;
    h_2 = 'b00000101001011110101;
    h_3 = 'b00000110001001111100;
    h_4 = 'b00000101100000101011;
    h_5 = 'b00000100000010000111;
    h_6 = 'b00000011101001010010;
    h_7 = 'b00000010100011011011;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000010011000001100;
    x_1 = 'b00000011110111010001;
    x_2 = 'b00000100100000001001;
    x_3 = 'b00000101011110011011;
    x_4 = 'b00000100101001000111;
    x_5 = 'b00000010110100011101;
    x_6 = 'b00000010100100110100;
    x_7 = 'b00000001010111000101;
    x_8 = 'b00000011100100100011;
    x_9 = 'b00000100101001100000;
    x_10 = 'b00000101000011011111;
    x_11 = 'b00000101111000010000;
    x_12 = 'b00000011110011001111;
    x_13 = 'b00000001101000010010;
    x_14 = 'b00000011111101101010;
    x_15 = 'b00000100111000110111;

    h_0 = 'b00000010011000001100;
    h_1 = 'b00000011110111010001;
    h_2 = 'b00000100100000001001;
    h_3 = 'b00000101011110011011;
    h_4 = 'b00000100101001000111;
    h_5 = 'b00000010110100011101;
    h_6 = 'b00000010100100110100;
    h_7 = 'b00000001010111000101;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000011000100100101;
    x_1 = 'b00000100101000001101;
    x_2 = 'b00000101011111010001;
    x_3 = 'b00000110100110111100;
    x_4 = 'b00000101110100111001;
    x_5 = 'b00000100010010110000;
    x_6 = 'b00000011100011000100;
    x_7 = 'b00000000110011011101;
    x_8 = 'b00000100000011100000;
    x_9 = 'b00000101010110100110;
    x_10 = 'b00000110000111111111;
    x_11 = 'b00000111010011111110;
    x_12 = 'b00000101110100000000;
    x_13 = 'b00000011100010111100;
    x_14 = 'b00000010011001011101;
    x_15 = 'b00000100100100100001;

    h_0 = 'b00000011000100100101;
    h_1 = 'b00000100101000001101;
    h_2 = 'b00000101011111010001;
    h_3 = 'b00000110100110111100;
    h_4 = 'b00000101110100111001;
    h_5 = 'b00000100010010110000;
    h_6 = 'b00000011100011000100;
    h_7 = 'b00000000110011011101;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000011000100100101;
    x_1 = 'b00000100010100101000;
    x_2 = 'b00000101001011110101;
    x_3 = 'b00000110101011110001;
    x_4 = 'b00000110001001000110;
    x_5 = 'b00000100111001100101;
    x_6 = 'b00000100101101101111;
    x_7 = 'b00000001000111110100;
    x_8 = 'b00000011011111011001;
    x_9 = 'b00000100100100011111;
    x_10 = 'b00000101101111100001;
    x_11 = 'b00000111010011111110;
    x_12 = 'b00000110010111001000;
    x_13 = 'b00000100110100101101;
    x_14 = 'b00000010010100001100;
    x_15 = 'b00000100000000111011;

    h_0 = 'b00000011000100100101;
    h_1 = 'b00000100010100101000;
    h_2 = 'b00000101001011110101;
    h_3 = 'b00000110101011110001;
    h_4 = 'b00000110001001000110;
    h_5 = 'b00000100111001100101;
    h_6 = 'b00000100101101101111;
    h_7 = 'b00000001000111110100;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000010111010101110;
    x_1 = 'b00000011101101011110;
    x_2 = 'b00000100101110101101;
    x_3 = 'b00000101111011011100;
    x_4 = 'b00000101011011101000;
    x_5 = 'b00000100011101110110;
    x_6 = 'b00000100101101101111;
    x_7 = 'b00000000101110010111;
    x_8 = 'b00000010100110101011;
    x_9 = 'b00000011101000010111;
    x_10 = 'b00000100101011000001;
    x_11 = 'b00000110100001000001;
    x_12 = 'b00000101100010011100;
    x_13 = 'b00000101001001001010;
    x_14 = 'b00000001101111010001;
    x_15 = 'b00000011000011111001;

    h_0 = 'b00000010111010101110;
    h_1 = 'b00000011101101011110;
    h_2 = 'b00000100101110101101;
    h_3 = 'b00000101111011011100;
    h_4 = 'b00000101011011101000;
    h_5 = 'b00000100011101110110;
    h_6 = 'b00000100101101101111;
    h_7 = 'b00000000101110010111;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000010001001011001;
    x_1 = 'b00000010011010010001;
    x_2 = 'b00000011001101100101;
    x_3 = 'b00000100010001000101;
    x_4 = 'b00000011110110100101;
    x_5 = 'b00000010011000101110;
    x_6 = 'b00000001110011000010;
    x_7 = 'b00000001000010101110;
    x_8 = 'b00000001111101011010;
    x_9 = 'b00000010100010001101;
    x_10 = 'b00000011010010111101;
    x_11 = 'b00000100100110101110;
    x_12 = 'b00000011010000000111;
    x_13 = 'b00000001000110001101;
    x_14 = 'b00000010010100001100;
    x_15 = 'b00000011001110000100;

    h_0 = 'b00000010001001011001;
    h_1 = 'b00000010011010010001;
    h_2 = 'b00000011001101100101;
    h_3 = 'b00000100010001000101;
    h_4 = 'b00000011110110100101;
    h_5 = 'b00000010011000101110;
    h_6 = 'b00000001110011000010;
    h_7 = 'b00000001000010101110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000000110000100110;
    x_1 = 'b00000000111000011001;
    x_2 = 'b00000001010100001100;
    x_3 = 'b00000010000100111001;
    x_4 = 'b00000001101001001000;
    x_5 = 'b11111111111101011001;
    x_6 = 'b11111111011101101011;
    x_7 = 'b11111111111011011110;
    x_8 = 'b00000001100011101000;
    x_9 = 'b00000001110101000110;
    x_10 = 'b00000010001001100101;
    x_11 = 'b00000010001101110101;
    x_12 = 'b00000001011011000011;
    x_13 = 'b11111111011111111111;
    x_14 = 'b00000011000011101001;
    x_15 = 'b00000011100010011010;

    h_0 = 'b00000000110000100110;
    h_1 = 'b00000000111000011001;
    h_2 = 'b00000001010100001100;
    h_3 = 'b00000010000100111001;
    h_4 = 'b00000001101001001000;
    h_5 = 'b11111111111101011001;
    h_6 = 'b11111111011101101011;
    h_7 = 'b11111111111011011110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000010100110111111;
    x_1 = 'b00000010000001110011;
    x_2 = 'b00000001111111111001;
    x_3 = 'b00000010000100111001;
    x_4 = 'b00000001100100000101;
    x_5 = 'b11111111100111001101;
    x_6 = 'b11111111010111011100;
    x_7 = 'b00000001101011011100;
    x_8 = 'b00000010011100010110;
    x_9 = 'b00000010001001001001;
    x_10 = 'b00000001110001000111;
    x_11 = 'b00000001111001011101;
    x_12 = 'b00000000110010000101;
    x_13 = 'b11111111011001001011;
    x_14 = 'b00000100000010111011;
    x_15 = 'b00000011111011110101;

    h_0 = 'b00000010100110111111;
    h_1 = 'b00000010000001110011;
    h_2 = 'b00000001111111111001;
    h_3 = 'b00000010000100111001;
    h_4 = 'b00000001100100000101;
    h_5 = 'b11111111100111001101;
    h_6 = 'b11111111010111011100;
    h_7 = 'b00000001101011011100;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000010101011111011;
    x_1 = 'b00000010010000011111;
    x_2 = 'b00000010001001100111;
    x_3 = 'b00000010001110100100;
    x_4 = 'b00000001001111111000;
    x_5 = 'b11111111000101111011;
    x_6 = 'b11111110111110100011;
    x_7 = 'b00000001111111110011;
    x_8 = 'b00000010010010000010;
    x_9 = 'b00000001110000000110;
    x_10 = 'b00000001100111010101;
    x_11 = 'b00000001100101000100;
    x_12 = 'b11111111111101011010;
    x_13 = 'b11111110001110001110;
    x_14 = 'b00000011111101101010;
    x_15 = 'b00000011011101010100;

    h_0 = 'b00000010101011111011;
    h_1 = 'b00000010010000011111;
    h_2 = 'b00000010001001100111;
    h_3 = 'b00000010001110100100;
    h_4 = 'b00000001001111111000;
    h_5 = 'b11111111000101111011;
    h_6 = 'b11111110111110100011;
    h_7 = 'b00000001111111110011;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000001111010100110;
    x_1 = 'b00000000101110100110;
    x_2 = 'b00000001000000110001;
    x_3 = 'b00000001100111111001;
    x_4 = 'b11111111101111111000;
    x_5 = 'b11111101100111101000;
    x_6 = 'b11111101101101101001;
    x_7 = 'b00000000000101101001;
    x_8 = 'b00000000110101001101;
    x_9 = 'b00000000110011111101;
    x_10 = 'b00000001000000001100;
    x_11 = 'b00000000011101101110;
    x_12 = 'b11111110101011011101;
    x_13 = 'b11111101011110100001;
    x_14 = 'b00000001111001110100;
    x_15 = 'b00000001110111100111;

    h_0 = 'b00000001111010100110;
    h_1 = 'b00000000101110100110;
    h_2 = 'b00000001000000110001;
    h_3 = 'b00000001100111111001;
    h_4 = 'b11111111101111111000;
    h_5 = 'b11111101100111101000;
    h_6 = 'b11111101101101101001;
    h_7 = 'b00000000000101101001;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000010011101001000;
    x_1 = 'b00000001011010101001;
    x_2 = 'b00000001011001000011;
    x_3 = 'b00000001101100101110;
    x_4 = 'b00000000001001001001;
    x_5 = 'b11111101110010101110;
    x_6 = 'b11111100111011110111;
    x_7 = 'b00000001101011011100;
    x_8 = 'b00000001111101011010;
    x_9 = 'b00000010000100001000;
    x_10 = 'b00000010011000010000;
    x_11 = 'b00000010001000101111;
    x_12 = 'b11111111100101111111;
    x_13 = 'b11111110000000100110;
    x_14 = 'b00000010101001010010;
    x_15 = 'b00000011001000111111;

    h_0 = 'b00000010011101001000;
    h_1 = 'b00000001011010101001;
    h_2 = 'b00000001011001000011;
    h_3 = 'b00000001101100101110;
    h_4 = 'b00000000001001001001;
    h_5 = 'b11111101110010101110;
    h_6 = 'b11111100111011110111;
    h_7 = 'b00000001101011011100;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000011010011011000;
    x_1 = 'b00000011001011001110;
    x_2 = 'b00000011011100001010;
    x_3 = 'b00000011111101110000;
    x_4 = 'b00000011000100000100;
    x_5 = 'b00000000100100001110;
    x_6 = 'b11111111101010000111;
    x_7 = 'b00000010110111110010;
    x_8 = 'b00000011101001101101;
    x_9 = 'b00000011110010011000;
    x_10 = 'b00000100010111011101;
    x_11 = 'b00000100100001100111;
    x_12 = 'b00000010111000101101;
    x_13 = 'b00000001000110001101;
    x_14 = 'b00000100100111110110;
    x_15 = 'b00000100011111011011;

    h_0 = 'b00000011010011011000;
    h_1 = 'b00000011001011001110;
    h_2 = 'b00000011011100001010;
    h_3 = 'b00000011111101110000;
    h_4 = 'b00000011000100000100;
    h_5 = 'b00000000100100001110;
    h_6 = 'b11111111101010000111;
    h_7 = 'b00000010110111110010;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000000100110101111;
    x_1 = 'b00000000111000011001;
    x_2 = 'b11111100111111011010;
    x_3 = 'b11111101111111110111;
    x_4 = 'b11111101100111011110;
    x_5 = 'b11111101000110010110;
    x_6 = 'b11111110011111011100;
    x_7 = 'b00000010001001111111;
    x_8 = 'b00000000000110110011;
    x_9 = 'b11111110100010101000;
    x_10 = 'b11111101011111001000;
    x_11 = 'b11111011110110001011;
    x_12 = 'b11111100001101011011;
    x_13 = 'b11111100101110110101;
    x_14 = 'b00000011000011101001;
    x_15 = 'b00000001000100110000;

    h_0 = 'b00000000100110101111;
    h_1 = 'b00000000111000011001;
    h_2 = 'b11111100111111011010;
    h_3 = 'b11111101111111110111;
    h_4 = 'b11111101100111011110;
    h_5 = 'b11111101000110010110;
    h_6 = 'b11111110011111011100;
    h_7 = 'b00000010001001111111;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000010100110111111;
    x_1 = 'b00000011000001011011;
    x_2 = 'b00000000000001101001;
    x_3 = 'b00000000101001000011;
    x_4 = 'b11111111101010110101;
    x_5 = 'b11111111000101111011;
    x_6 = 'b11111111110000010110;
    x_7 = 'b00000100101100110110;
    x_8 = 'b00000010010010000010;
    x_9 = 'b00000000111000111110;
    x_10 = 'b00000000000000100101;
    x_11 = 'b11111110101101100111;
    x_12 = 'b11111111000010111000;
    x_13 = 'b11111111011001001011;
    x_14 = 'b00000011000011101001;
    x_15 = 'b00000010100000010011;

    h_0 = 'b00000010100110111111;
    h_1 = 'b00000011000001011011;
    h_2 = 'b00000000000001101001;
    h_3 = 'b00000000101001000011;
    h_4 = 'b11111111101010110101;
    h_5 = 'b11111111000101111011;
    h_6 = 'b11111111110000010110;
    h_7 = 'b00000100101100110110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000100100111001111;
    x_1 = 'b00000100001010110110;
    x_2 = 'b00000001001111010101;
    x_3 = 'b00000001011001011001;
    x_4 = 'b00000000000100000110;
    x_5 = 'b11111111100111001101;
    x_6 = 'b11111111101010000111;
    x_7 = 'b00000101010000011110;
    x_8 = 'b00000010100001100001;
    x_9 = 'b00000001100001000011;
    x_10 = 'b00000000011101111100;
    x_11 = 'b00000000000100010000;
    x_12 = 'b00000000001110111110;
    x_13 = 'b11111111011001001011;
    x_14 = 'b00000011100011010010;
    x_15 = 'b00000010101111100011;

    h_0 = 'b00000100100111001111;
    h_1 = 'b00000100001010110110;
    h_2 = 'b00000001001111010101;
    h_3 = 'b00000001011001011001;
    h_4 = 'b00000000000100000110;
    h_5 = 'b11111111100111001101;
    h_6 = 'b11111111101010000111;
    h_7 = 'b00000101010000011110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000111001010000001;
    x_1 = 'b00000110101100010111;
    x_2 = 'b00000011110100011100;
    x_3 = 'b00000011100000110000;
    x_4 = 'b00000010111001111101;
    x_5 = 'b00000010101110111010;
    x_6 = 'b00000001111111011111;
    x_7 = 'b00000111010100110100;
    x_8 = 'b00000101010000110111;
    x_9 = 'b00000100101001100000;
    x_10 = 'b00000100001000110010;
    x_11 = 'b00000011100100011110;
    x_12 = 'b00000100110011101000;
    x_13 = 'b00000011111110001100;
    x_14 = 'b00000110000110110001;
    x_15 = 'b00000101111010111110;

    h_0 = 'b00000111001010000001;
    h_1 = 'b00000110101100010111;
    h_2 = 'b00000011110100011100;
    h_3 = 'b00000011100000110000;
    h_4 = 'b00000010111001111101;
    h_5 = 'b00000010101110111010;
    h_6 = 'b00000001111111011111;
    h_7 = 'b00000111010100110100;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000010111010101110;
    x_1 = 'b00000011001011001110;
    x_2 = 'b00000001000000110001;
    x_3 = 'b00000001000110000011;
    x_4 = 'b00000001100100000101;
    x_5 = 'b00000001111100111111;
    x_6 = 'b00000010100100110100;
    x_7 = 'b00000011001100001001;
    x_8 = 'b00000010000010100100;
    x_9 = 'b00000001110000000110;
    x_10 = 'b00000001101100001110;
    x_11 = 'b00000001111110100011;
    x_12 = 'b00000100011100001101;
    x_13 = 'b00000100101101111001;
    x_14 = 'b00000011000011101001;
    x_15 = 'b00000010111001101110;

    h_0 = 'b00000010111010101110;
    h_1 = 'b00000011001011001110;
    h_2 = 'b00000001000000110001;
    h_3 = 'b00000001000110000011;
    h_4 = 'b00000001100100000101;
    h_5 = 'b00000001111100111111;
    h_6 = 'b00000010100100110100;
    h_7 = 'b00000011001100001001;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000000110000100110;
    x_1 = 'b00000001011010101001;
    x_2 = 'b11111111101001010111;
    x_3 = 'b00000000010000111000;
    x_4 = 'b00000001000101110001;
    x_5 = 'b00000001110001111001;
    x_6 = 'b00000010100100110100;
    x_7 = 'b00000010101101100111;
    x_8 = 'b00000000111010010111;
    x_9 = 'b00000001000010111111;
    x_10 = 'b00000001011000101001;
    x_11 = 'b00000010000011101001;
    x_12 = 'b00000011111001000110;
    x_13 = 'b00000100110100101101;
    x_14 = 'b00000010110011110101;
    x_15 = 'b00000010011011001101;

    h_0 = 'b00000000110000100110;
    h_1 = 'b00000001011010101001;
    h_2 = 'b11111111101001010111;
    h_3 = 'b00000000010000111000;
    h_4 = 'b00000001000101110001;
    h_5 = 'b00000001110001111001;
    h_6 = 'b00000010100100110100;
    h_7 = 'b00000010101101100111;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000100110001000111;
    x_1 = 'b00000100001010110110;
    x_2 = 'b00000001011001000011;
    x_3 = 'b00000010000100111001;
    x_4 = 'b00000001101001001000;
    x_5 = 'b00000001110001111001;
    x_6 = 'b00000010011110100110;
    x_7 = 'b00000110101100000110;
    x_8 = 'b00000011100100100011;
    x_9 = 'b00000010101100001110;
    x_10 = 'b00000010101011110100;
    x_11 = 'b00000010011000000010;
    x_12 = 'b00000011001010010001;
    x_13 = 'b00000011100010111100;
    x_14 = 'b00000110000110110001;
    x_15 = 'b00000100011111011011;

    h_0 = 'b00000100110001000111;
    h_1 = 'b00000100001010110110;
    h_2 = 'b00000001011001000011;
    h_3 = 'b00000010000100111001;
    h_4 = 'b00000001101001001000;
    h_5 = 'b00000001110001111001;
    h_6 = 'b00000010011110100110;
    h_7 = 'b00000110101100000110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000001000100010101;
    x_1 = 'b00000001101110001110;
    x_2 = 'b11111111110111111100;
    x_3 = 'b00000000110111100011;
    x_4 = 'b11111111111001111111;
    x_5 = 'b11111111100001101010;
    x_6 = 'b00000000011011111010;
    x_7 = 'b00000011001100001001;
    x_8 = 'b00000001011001010100;
    x_9 = 'b00000001011100000011;
    x_10 = 'b00000001100010011100;
    x_11 = 'b00000000001001010110;
    x_12 = 'b00000000111101110010;
    x_13 = 'b00000000010110100000;
    x_14 = 'b00000100011101010011;
    x_15 = 'b00000011000011111001;

    h_0 = 'b00000001000100010101;
    h_1 = 'b00000001101110001110;
    h_2 = 'b11111111110111111100;
    h_3 = 'b00000000110111100011;
    h_4 = 'b11111111111001111111;
    h_5 = 'b11111111100001101010;
    h_6 = 'b00000000011011111010;
    h_7 = 'b00000011001100001001;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000001001001010001;
    x_1 = 'b00000010010000011111;
    x_2 = 'b00000000011110110010;
    x_3 = 'b00000001001111101110;
    x_4 = 'b11111111111111000010;
    x_5 = 'b11111111000101111011;
    x_6 = 'b11111110101011111000;
    x_7 = 'b00000101010000011110;
    x_8 = 'b00000010110000111111;
    x_9 = 'b00000010101100001110;
    x_10 = 'b00000010100010000010;
    x_11 = 'b00000001010000101100;
    x_12 = 'b00000001011011000011;
    x_13 = 'b11111111110100011100;
    x_14 = 'b00000110000110110001;
    x_15 = 'b00000100111000110111;

    h_0 = 'b00000001001001010001;
    h_1 = 'b00000010010000011111;
    h_2 = 'b00000000011110110010;
    h_3 = 'b00000001001111101110;
    h_4 = 'b11111111111111000010;
    h_5 = 'b11111111000101111011;
    h_6 = 'b11111110101011111000;
    h_7 = 'b00000101010000011110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000001010011001000;
    x_1 = 'b00000011000110010100;
    x_2 = 'b00000001110001010101;
    x_3 = 'b00000010110000011010;
    x_4 = 'b00000001001111111000;
    x_5 = 'b00000000101111010100;
    x_6 = 'b00000000010101101011;
    x_7 = 'b00000100000100001000;
    x_8 = 'b00000010110110001001;
    x_9 = 'b00000010110110010000;
    x_10 = 'b00000010101011110100;
    x_11 = 'b00000001111001011101;
    x_12 = 'b00000010001001111000;
    x_13 = 'b00000000110001110001;
    x_14 = 'b00000100000010111011;
    x_15 = 'b00000011011000001111;

    h_0 = 'b00000001010011001000;
    h_1 = 'b00000011000110010100;
    h_2 = 'b00000001110001010101;
    h_3 = 'b00000010110000011010;
    h_4 = 'b00000001001111111000;
    h_5 = 'b00000000101111010100;
    h_6 = 'b00000000010101101011;
    h_7 = 'b00000100000100001000;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111111001101111101;
    x_1 = 'b00000000101110100110;
    x_2 = 'b00000000000110100000;
    x_3 = 'b00000001001010111001;
    x_4 = 'b11111111111111000010;
    x_5 = 'b11111111110010010011;
    x_6 = 'b00000000001001001111;
    x_7 = 'b00000000100100001100;
    x_8 = 'b11111111110111010100;
    x_9 = 'b00000000111101111110;
    x_10 = 'b00000001000101000101;
    x_11 = 'b00000000000100010000;
    x_12 = 'b00000000101100001111;
    x_13 = 'b00000000010110100000;
    x_14 = 'b00000000101010101110;
    x_15 = 'b00000001001001110110;

    h_0 = 'b11111111001101111101;
    h_1 = 'b00000000101110100110;
    h_2 = 'b00000000000110100000;
    h_3 = 'b00000001001010111001;
    h_4 = 'b11111111111111000010;
    h_5 = 'b11111111110010010011;
    h_6 = 'b00000000001001001111;
    h_7 = 'b00000000100100001100;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000001000100010101;
    x_1 = 'b00000001000111000100;
    x_2 = 'b11111111110011000101;
    x_3 = 'b00000000000111001110;
    x_4 = 'b11111110111101010111;
    x_5 = 'b11111110110101010010;
    x_6 = 'b11111111100011111001;
    x_7 = 'b00000011000001111110;
    x_8 = 'b00000000110000000011;
    x_9 = 'b00000001001000000000;
    x_10 = 'b00000001000101000101;
    x_11 = 'b11111111010110011001;
    x_12 = 'b11111111100101111111;
    x_13 = 'b11111111000100101111;
    x_14 = 'b00000010010100001100;
    x_15 = 'b00000010000110110111;

    h_0 = 'b00000001000100010101;
    h_1 = 'b00000001000111000100;
    h_2 = 'b11111111110011000101;
    h_3 = 'b00000000000111001110;
    h_4 = 'b11111110111101010111;
    h_5 = 'b11111110110101010010;
    h_6 = 'b11111111100011111001;
    h_7 = 'b00000011000001111110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000001010011001000;
    x_1 = 'b00000001010000110111;
    x_2 = 'b11111111011010110011;
    x_3 = 'b11111111100101011000;
    x_4 = 'b11111110000000101111;
    x_5 = 'b11111101000110010110;
    x_6 = 'b11111110000000010100;
    x_7 = 'b00000011011011011010;
    x_8 = 'b00000001101000110010;
    x_9 = 'b00000001000010111111;
    x_10 = 'b00000000011001000011;
    x_11 = 'b11111111001100001100;
    x_12 = 'b11111110000010011111;
    x_13 = 'b11111101010000111001;
    x_14 = 'b00000010110011110101;
    x_15 = 'b00000010000001110010;

    h_0 = 'b00000001010011001000;
    h_1 = 'b00000001010000110111;
    h_2 = 'b11111111011010110011;
    h_3 = 'b11111111100101011000;
    h_4 = 'b11111110000000101111;
    h_5 = 'b11111101000110010110;
    h_6 = 'b11111110000000010100;
    h_7 = 'b00000011011011011010;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000010111111101010;
    x_1 = 'b00000011100011101100;
    x_2 = 'b00000001100111100111;
    x_3 = 'b00000001111011001111;
    x_4 = 'b00000000110110100111;
    x_5 = 'b11111111100111001101;
    x_6 = 'b00000000101110100101;
    x_7 = 'b00000101100100110101;
    x_8 = 'b00000011101001101101;
    x_9 = 'b00000011001010010010;
    x_10 = 'b00000010101011110100;
    x_11 = 'b00000001001011100110;
    x_12 = 'b00000000000011010000;
    x_13 = 'b00000000111000100101;
    x_14 = 'b00000100001000001101;
    x_15 = 'b00000011100010011010;

    h_0 = 'b00000010111111101010;
    h_1 = 'b00000011100011101100;
    h_2 = 'b00000001100111100111;
    h_3 = 'b00000001111011001111;
    h_4 = 'b00000000110110100111;
    h_5 = 'b11111111100111001101;
    h_6 = 'b00000000101110100101;
    h_7 = 'b00000101100100110101;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000011111010110110;
    x_1 = 'b00000100000001000011;
    x_2 = 'b00000001110001010101;
    x_3 = 'b00000010110101001111;
    x_4 = 'b00000001010100111011;
    x_5 = 'b11111111111101011001;
    x_6 = 'b00000000000011000001;
    x_7 = 'b00000101000110010011;
    x_8 = 'b00000011000101100111;
    x_9 = 'b00000010101100001110;
    x_10 = 'b00000010001110011110;
    x_11 = 'b11111111110100111101;
    x_12 = 'b11111110110111001010;
    x_13 = 'b11111110001110001110;
    x_14 = 'b00000011101101110101;
    x_15 = 'b00000010011011001101;

    h_0 = 'b00000011111010110110;
    h_1 = 'b00000100000001000011;
    h_2 = 'b00000001110001010101;
    h_3 = 'b00000010110101001111;
    h_4 = 'b00000001010100111011;
    h_5 = 'b11111111111101011001;
    h_6 = 'b00000000000011000001;
    h_7 = 'b00000101000110010011;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000001100001111011;
    x_1 = 'b00000010100100000100;
    x_2 = 'b11111111110011000101;
    x_3 = 'b00000010010011011010;
    x_4 = 'b00000000110001100100;
    x_5 = 'b11111111000000011000;
    x_6 = 'b11111111010111011100;
    x_7 = 'b00000011100101100110;
    x_8 = 'b00000001110011000110;
    x_9 = 'b00000001100110000100;
    x_10 = 'b00000001000101000101;
    x_11 = 'b11111111010110011001;
    x_12 = 'b11111111000010111000;
    x_13 = 'b11111101100101010101;
    x_14 = 'b00000010110011110101;
    x_15 = 'b00000001010100000001;

    h_0 = 'b00000001100001111011;
    h_1 = 'b00000010100100000100;
    h_2 = 'b11111111110011000101;
    h_3 = 'b00000010010011011010;
    h_4 = 'b00000000110001100100;
    h_5 = 'b11111111000000011000;
    h_6 = 'b11111111010111011100;
    h_7 = 'b00000011100101100110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111110101011011011;
    x_1 = 'b11111110100101100100;
    x_2 = 'b11111110000011011001;
    x_3 = 'b11111110001001100010;
    x_4 = 'b11111101011101011000;
    x_5 = 'b11111011011100111101;
    x_6 = 'b11111010111111011001;
    x_7 = 'b11111111100111000111;
    x_8 = 'b11111110000101110111;
    x_9 = 'b11111101100110100000;
    x_10 = 'b11111101011111001000;
    x_11 = 'b11111100101001001000;
    x_12 = 'b11111011100100011101;
    x_13 = 'b11111001000000010101;
    x_14 = 'b11111111101011011100;
    x_15 = 'b11111110010111110111;

    h_0 = 'b11111110101011011011;
    h_1 = 'b11111110100101100100;
    h_2 = 'b11111110000011011001;
    h_3 = 'b11111110001001100010;
    h_4 = 'b11111101011101011000;
    h_5 = 'b11111011011100111101;
    h_6 = 'b11111010111111011001;
    h_7 = 'b11111111100111000111;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111100011100011000;
    x_1 = 'b11111100011100100001;
    x_2 = 'b11111011110110100101;
    x_3 = 'b11111011101010000000;
    x_4 = 'b11111011011010000001;
    x_5 = 'b11111001111001000110;
    x_6 = 'b11111001111010111011;
    x_7 = 'b11111110101010000010;
    x_8 = 'b11111100111101101010;
    x_9 = 'b11111100010001010100;
    x_10 = 'b11111100010000110111;
    x_11 = 'b11111100000000010111;
    x_12 = 'b11111011110000001010;
    x_13 = 'b11111010001011010010;
    x_14 = 'b11111110110001011011;
    x_15 = 'b11111101101111001011;

    h_0 = 'b11111100011100011000;
    h_1 = 'b11111100011100100001;
    h_2 = 'b11111011110110100101;
    h_3 = 'b11111011101010000000;
    h_4 = 'b11111011011010000001;
    h_5 = 'b11111001111001000110;
    h_6 = 'b11111001111010111011;
    h_7 = 'b11111110101010000010;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111100001101100100;
    x_1 = 'b11111100000100000011;
    x_2 = 'b11111011011001011100;
    x_3 = 'b11111011101010000000;
    x_4 = 'b11111011011010000001;
    x_5 = 'b11111010011010011001;
    x_6 = 'b11111001101110011111;
    x_7 = 'b11111110001011100000;
    x_8 = 'b11111101000010110100;
    x_9 = 'b11111100111001011001;
    x_10 = 'b11111101100100000010;
    x_11 = 'b11111101110101100100;
    x_12 = 'b11111101010011101010;
    x_13 = 'b11111100010011100100;
    x_14 = 'b11111101110010001001;
    x_15 = 'b11111110001000100110;

    h_0 = 'b11111100001101100100;
    h_1 = 'b11111100000100000011;
    h_2 = 'b11111011011001011100;
    h_3 = 'b11111011101010000000;
    h_4 = 'b11111011011010000001;
    h_5 = 'b11111010011010011001;
    h_6 = 'b11111001101110011111;
    h_7 = 'b11111110001011100000;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111101100110010111;
    x_1 = 'b11111110101010011101;
    x_2 = 'b11111110010110110100;
    x_3 = 'b11111110100001101101;
    x_4 = 'b11111110010100111100;
    x_5 = 'b11111101011100100010;
    x_6 = 'b11111100111011110111;
    x_7 = 'b00000000101001010010;
    x_8 = 'b11111111110010001010;
    x_9 = 'b11111111110010110100;
    x_10 = 'b00000000100010110101;
    x_11 = 'b00000000101101000001;
    x_12 = 'b11111111110111100011;
    x_13 = 'b11111110011011110110;
    x_14 = 'b00000000111111110100;
    x_15 = 'b00000000111111101011;

    h_0 = 'b11111101100110010111;
    h_1 = 'b11111110101010011101;
    h_2 = 'b11111110010110110100;
    h_3 = 'b11111110100001101101;
    h_4 = 'b11111110010100111100;
    h_5 = 'b11111101011100100010;
    h_6 = 'b11111100111011110111;
    h_7 = 'b00000000101001010010;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111111100001101011;
    x_1 = 'b00000000101110100110;
    x_2 = 'b11111111110111111100;
    x_3 = 'b11111111100000100011;
    x_4 = 'b11111111000010011010;
    x_5 = 'b11111110001000111010;
    x_6 = 'b11111101111010000110;
    x_7 = 'b00000010111100111000;
    x_8 = 'b00000001011001010100;
    x_9 = 'b00000001000010111111;
    x_10 = 'b00000001001110110111;
    x_11 = 'b00000000001110011100;
    x_12 = 'b11111111101011110110;
    x_13 = 'b11111100110101101001;
    x_14 = 'b00000010111001000110;
    x_15 = 'b00000010011011001101;

    h_0 = 'b11111111100001101011;
    h_1 = 'b00000000101110100110;
    h_2 = 'b11111111110111111100;
    h_3 = 'b11111111100000100011;
    h_4 = 'b11111111000010011010;
    h_5 = 'b11111110001000111010;
    h_6 = 'b11111101111010000110;
    h_7 = 'b00000010111100111000;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000000010011000000;
    x_1 = 'b00000000001100010110;
    x_2 = 'b11111111000111011000;
    x_3 = 'b11111110010011001100;
    x_4 = 'b11111101101100100010;
    x_5 = 'b11111101000000110011;
    x_6 = 'b11111101001000010011;
    x_7 = 'b00000011000111000100;
    x_8 = 'b00000001001110111111;
    x_9 = 'b00000000010101111001;
    x_10 = 'b11111111111011101100;
    x_11 = 'b11111110010100001001;
    x_12 = 'b11111110011001111001;
    x_13 = 'b11111100011010011000;
    x_14 = 'b00000011011110000001;
    x_15 = 'b00000010100101011000;

    h_0 = 'b00000000010011000000;
    h_1 = 'b00000000001100010110;
    h_2 = 'b11111111000111011000;
    h_3 = 'b11111110010011001100;
    h_4 = 'b11111101101100100010;
    h_5 = 'b11111101000000110011;
    h_6 = 'b11111101001000010011;
    h_7 = 'b00000011000111000100;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000010011000001100;
    x_1 = 'b00000010010000011111;
    x_2 = 'b00000000101101010110;
    x_3 = 'b11111111101010001101;
    x_4 = 'b11111110111101010111;
    x_5 = 'b11111101111000010001;
    x_6 = 'b11111101110011110111;
    x_7 = 'b00000101100100110101;
    x_8 = 'b00000011100100100011;
    x_9 = 'b00000010011000001011;
    x_10 = 'b00000001011000101001;
    x_11 = 'b11111111101010110001;
    x_12 = 'b11111111011010010010;
    x_13 = 'b11111101101100001010;
    x_14 = 'b00000101111100001110;
    x_15 = 'b00000100111101111100;

    h_0 = 'b00000010011000001100;
    h_1 = 'b00000010010000011111;
    h_2 = 'b00000000101101010110;
    h_3 = 'b11111111101010001101;
    h_4 = 'b11111110111101010111;
    h_5 = 'b11111101111000010001;
    h_6 = 'b11111101110011110111;
    h_7 = 'b00000101100100110101;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000001111010100110;
    x_1 = 'b00000010010101011000;
    x_2 = 'b00000000101101010110;
    x_3 = 'b00000000000111001110;
    x_4 = 'b11111111010110101000;
    x_5 = 'b11111110000011010111;
    x_6 = 'b11111110000000010100;
    x_7 = 'b00000101001011011001;
    x_8 = 'b00000011111110010110;
    x_9 = 'b00000010101100001110;
    x_10 = 'b00000010011101001001;
    x_11 = 'b00000000110010000111;
    x_12 = 'b00000000011010101011;
    x_13 = 'b11111110011011110110;
    x_14 = 'b00000101010111010011;
    x_15 = 'b00000101001101001101;

    h_0 = 'b00000001111010100110;
    h_1 = 'b00000010010101011000;
    h_2 = 'b00000000101101010110;
    h_3 = 'b00000000000111001110;
    h_4 = 'b11111111010110101000;
    h_5 = 'b11111110000011010111;
    h_6 = 'b11111110000000010100;
    h_7 = 'b00000101001011011001;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000000010111111100;
    x_1 = 'b00000001000111000100;
    x_2 = 'b00000000010000001101;
    x_3 = 'b11111111101010001101;
    x_4 = 'b11111111000111011110;
    x_5 = 'b11111101100111101000;
    x_6 = 'b11111101011010111110;
    x_7 = 'b00000011011011011010;
    x_8 = 'b00000011001010110001;
    x_9 = 'b00000010100010001101;
    x_10 = 'b00000010100110111011;
    x_11 = 'b00000001000110100000;
    x_12 = 'b11111111110001101101;
    x_13 = 'b11111100100001001100;
    x_14 = 'b00000100100111110110;
    x_15 = 'b00000100101110101100;

    h_0 = 'b00000000010111111100;
    h_1 = 'b00000001000111000100;
    h_2 = 'b00000000010000001101;
    h_3 = 'b11111111101010001101;
    h_4 = 'b11111111000111011110;
    h_5 = 'b11111101100111101000;
    h_6 = 'b11111101011010111110;
    h_7 = 'b00000011011011011010;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000010001001011001;
    x_1 = 'b00000011101000100101;
    x_2 = 'b00000010110101010100;
    x_3 = 'b00000010011000001111;
    x_4 = 'b00000001011001111110;
    x_5 = 'b11111111010110100100;
    x_6 = 'b11111101111010000110;
    x_7 = 'b00000110010010101001;
    x_8 = 'b00000101100000010101;
    x_9 = 'b00000100111000100010;
    x_10 = 'b00000100010010100100;
    x_11 = 'b00000010110110100111;
    x_12 = 'b00000000110010000101;
    x_13 = 'b11111100011010011000;
    x_14 = 'b00000111100000011010;
    x_15 = 'b00000110100011101010;

    h_0 = 'b00000010001001011001;
    h_1 = 'b00000011101000100101;
    h_2 = 'b00000010110101010100;
    h_3 = 'b00000010011000001111;
    h_4 = 'b00000001011001111110;
    h_5 = 'b11111111010110100100;
    h_6 = 'b11111101111010000110;
    h_7 = 'b00000110010010101001;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000010110000110111;
    x_1 = 'b00000011011001111001;
    x_2 = 'b00000010101011100110;
    x_3 = 'b00000010100110101111;
    x_4 = 'b00000001101110001100;
    x_5 = 'b00000000001000011111;
    x_6 = 'b11111111100011111001;
    x_7 = 'b00000100110111000010;
    x_8 = 'b00000100011000001000;
    x_9 = 'b00000100000001011010;
    x_10 = 'b00000011110101001101;
    x_11 = 'b00000011001010111111;
    x_12 = 'b00000001100110110001;
    x_13 = 'b11111110111101111011;
    x_14 = 'b00000101100001110110;
    x_15 = 'b00000101001000000111;

    h_0 = 'b00000010110000110111;
    h_1 = 'b00000011011001111001;
    h_2 = 'b00000010101011100110;
    h_3 = 'b00000010100110101111;
    h_4 = 'b00000001101110001100;
    h_5 = 'b00000000001000011111;
    h_6 = 'b11111111100011111001;
    h_7 = 'b00000100110111000010;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000010100010000011;
    x_1 = 'b00000010100100000100;
    x_2 = 'b00000001110001010101;
    x_3 = 'b00000001111011001111;
    x_4 = 'b00000001001010110100;
    x_5 = 'b11111111111101011001;
    x_6 = 'b00000001000001010000;
    x_7 = 'b00000011101111110001;
    x_8 = 'b00000011001111111011;
    x_9 = 'b00000010110110010000;
    x_10 = 'b00000011001001001011;
    x_11 = 'b00000011010000000101;
    x_12 = 'b00000010001111101111;
    x_13 = 'b00000001101000010010;
    x_14 = 'b00000011111000011000;
    x_15 = 'b00000011111011110101;

    h_0 = 'b00000010100010000011;
    h_1 = 'b00000010100100000100;
    h_2 = 'b00000001110001010101;
    h_3 = 'b00000001111011001111;
    h_4 = 'b00000001001010110100;
    h_5 = 'b11111111111101011001;
    h_6 = 'b00000001000001010000;
    h_7 = 'b00000011101111110001;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000011100010001100;
    x_1 = 'b00000011111100001010;
    x_2 = 'b00000011100001000001;
    x_3 = 'b00000011001101011010;
    x_4 = 'b00000010011011101001;
    x_5 = 'b00000001100001010000;
    x_6 = 'b00000010010010001010;
    x_7 = 'b00000101000110010011;
    x_8 = 'b00000100101100110000;
    x_9 = 'b00000100000110011011;
    x_10 = 'b00000100001000110010;
    x_11 = 'b00000011111000110110;
    x_12 = 'b00000011100001101011;
    x_13 = 'b00000010000011100010;
    x_14 = 'b00000100111100111100;
    x_15 = 'b00000100011111011011;

    h_0 = 'b00000011100010001100;
    h_1 = 'b00000011111100001010;
    h_2 = 'b00000011100001000001;
    h_3 = 'b00000011001101011010;
    h_4 = 'b00000010011011101001;
    h_5 = 'b00000001100001010000;
    h_6 = 'b00000010010010001010;
    h_7 = 'b00000101000110010011;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000011010011011000;
    x_1 = 'b00000100000101111101;
    x_2 = 'b00000011010010011100;
    x_3 = 'b00000010111010000101;
    x_4 = 'b00000001111101010110;
    x_5 = 'b00000001010000100110;
    x_6 = 'b00000001101100110100;
    x_7 = 'b00000101101001111011;
    x_8 = 'b00000100110111000100;
    x_9 = 'b00000100010101011101;
    x_10 = 'b00000100010111011101;
    x_11 = 'b00000011011010010010;
    x_12 = 'b00000011010000000111;
    x_13 = 'b00000001100001011110;
    x_14 = 'b00000101111100001110;
    x_15 = 'b00000100111101111100;

    h_0 = 'b00000011010011011000;
    h_1 = 'b00000100000101111101;
    h_2 = 'b00000011010010011100;
    h_3 = 'b00000010111010000101;
    h_4 = 'b00000001111101010110;
    h_5 = 'b00000001010000100110;
    h_6 = 'b00000001101100110100;
    h_7 = 'b00000101101001111011;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000100101100001011;
    x_1 = 'b00000101011110000011;
    x_2 = 'b00000100011011010010;
    x_3 = 'b00000100011111100101;
    x_4 = 'b00000011010011001110;
    x_5 = 'b00000001110001111001;
    x_6 = 'b00000001100110100101;
    x_7 = 'b00000110100001111010;
    x_8 = 'b00000101101010101001;
    x_9 = 'b00000110001000101101;
    x_10 = 'b00000110000011000101;
    x_11 = 'b00000101010100100101;
    x_12 = 'b00000100010000100000;
    x_13 = 'b00000010001010010110;
    x_14 = 'b00000101010111010011;
    x_15 = 'b00000101100110101000;

    h_0 = 'b00000100101100001011;
    h_1 = 'b00000101011110000011;
    h_2 = 'b00000100011011010010;
    h_3 = 'b00000100011111100101;
    h_4 = 'b00000011010011001110;
    h_5 = 'b00000001110001111001;
    h_6 = 'b00000001100110100101;
    h_7 = 'b00000110100001111010;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000010101011111011;
    x_1 = 'b00000011011110110011;
    x_2 = 'b00000011001000101111;
    x_3 = 'b00000011111101110000;
    x_4 = 'b00000011000100000100;
    x_5 = 'b00000001100001010000;
    x_6 = 'b00000001111001010000;
    x_7 = 'b00000010110111110010;
    x_8 = 'b00000011111110010110;
    x_9 = 'b00000100011111011111;
    x_10 = 'b00000100101111111010;
    x_11 = 'b00000100010010010101;
    x_12 = 'b00000100000100110011;
    x_13 = 'b00000010000011100010;
    x_14 = 'b00000011101000100100;
    x_15 = 'b00000100010000001011;

    h_0 = 'b00000010101011111011;
    h_1 = 'b00000011011110110011;
    h_2 = 'b00000011001000101111;
    h_3 = 'b00000011111101110000;
    h_4 = 'b00000011000100000100;
    h_5 = 'b00000001100001010000;
    h_6 = 'b00000001111001010000;
    h_7 = 'b00000010110111110010;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111100111001111110;
    x_1 = 'b11111010111111100001;
    x_2 = 'b11111000110100010110;
    x_3 = 'b11110110111110010011;
    x_4 = 'b11110111100010011110;
    x_5 = 'b11110111000010000011;
    x_6 = 'b11111000110000010000;
    x_7 = 'b11111101110111001001;
    x_8 = 'b11111000110001011110;
    x_9 = 'b11111000001100101111;
    x_10 = 'b11110111100110011011;
    x_11 = 'b11110110101010111100;
    x_12 = 'b11111000000000001011;
    x_13 = 'b11110110111000000010;
    x_14 = 'b11111010001111011000;
    x_15 = 'b11111001100001101001;

    h_0 = 'b11111100111001111110;
    h_1 = 'b11111010111111100001;
    h_2 = 'b11111000110100010110;
    h_3 = 'b11110110111110010011;
    h_4 = 'b11110111100010011110;
    h_5 = 'b11110111000010000011;
    h_6 = 'b11111000110000010000;
    h_7 = 'b11111101110111001001;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111010111001101110;
    x_1 = 'b11111001001110111101;
    x_2 = 'b11110110100111100010;
    x_3 = 'b11110100100011100111;
    x_4 = 'b11110100011101011100;
    x_5 = 'b11110011011110101000;
    x_6 = 'b11110110010100101010;
    x_7 = 'b11111011111100111111;
    x_8 = 'b11110111001010010101;
    x_9 = 'b11110110011110011111;
    x_10 = 'b11110101110001000000;
    x_11 = 'b11110101000101000001;
    x_12 = 'b11110101000100111000;
    x_13 = 'b11110101011000101001;
    x_14 = 'b11111001001010110101;
    x_15 = 'b11111000000110000111;

    h_0 = 'b11111010111001101110;
    h_1 = 'b11111001001110111101;
    h_2 = 'b11110110100111100010;
    h_3 = 'b11110100100011100111;
    h_4 = 'b11110100011101011100;
    h_5 = 'b11110011011110101000;
    h_6 = 'b11110110010100101010;
    h_7 = 'b11111011111100111111;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111011001000100001;
    x_1 = 'b11111001000101001010;
    x_2 = 'b11110111001001100001;
    x_3 = 'b11110101001111000111;
    x_4 = 'b11110101001010111010;
    x_5 = 'b11110100110001110101;
    x_6 = 'b11110111010010111001;
    x_7 = 'b11111100100101101101;
    x_8 = 'b11111000011100110110;
    x_9 = 'b11110111111000101100;
    x_10 = 'b11110111011100101000;
    x_11 = 'b11110110110101001000;
    x_12 = 'b11110101111111011010;
    x_13 = 'b11110110001111001010;
    x_14 = 'b11111010111110110110;
    x_15 = 'b11111001111011000101;

    h_0 = 'b11111011001000100001;
    h_1 = 'b11111001000101001010;
    h_2 = 'b11110111001001100001;
    h_3 = 'b11110101001111000111;
    h_4 = 'b11110101001010111010;
    h_5 = 'b11110100110001110101;
    h_6 = 'b11110111010010111001;
    h_7 = 'b11111100100101101101;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111101101011010011;
    x_1 = 'b11111100001000111100;
    x_2 = 'b11111001111101001100;
    x_3 = 'b11110111111101001001;
    x_4 = 'b11111000000000110010;
    x_5 = 'b11110111110011111110;
    x_6 = 'b11111010110010111100;
    x_7 = 'b00000000110011011101;
    x_8 = 'b11111011110101011101;
    x_9 = 'b11111011101110001111;
    x_10 = 'b11111011010001010000;
    x_11 = 'b11111001100010011001;
    x_12 = 'b11111001010111111110;
    x_13 = 'b11111001000111001001;
    x_14 = 'b11111110110001011011;
    x_15 = 'b11111101011010110101;

    h_0 = 'b11111101101011010011;
    h_1 = 'b11111100001000111100;
    h_2 = 'b11111001111101001100;
    h_3 = 'b11110111111101001001;
    h_4 = 'b11111000000000110010;
    h_5 = 'b11110111110011111110;
    h_6 = 'b11111010110010111100;
    h_7 = 'b00000000110011011101;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111111101011100011;
    x_1 = 'b11111110000011010011;
    x_2 = 'b11111100001010000000;
    x_3 = 'b11111010110000000000;
    x_4 = 'b11111010101100100011;
    x_5 = 'b11111010001111010011;
    x_6 = 'b11111101001000010011;
    x_7 = 'b00000001100110010110;
    x_8 = 'b11111100110011010110;
    x_9 = 'b11111101011100011110;
    x_10 = 'b11111101011111001000;
    x_11 = 'b11111011010111100110;
    x_12 = 'b11111011100100011101;
    x_13 = 'b11111011001000100111;
    x_14 = 'b11111101110010001001;
    x_15 = 'b11111101100101000000;

    h_0 = 'b11111111101011100011;
    h_1 = 'b11111110000011010011;
    h_2 = 'b11111100001010000000;
    h_3 = 'b11111010110000000000;
    h_4 = 'b11111010101100100011;
    h_5 = 'b11111010001111010011;
    h_6 = 'b11111101001000010011;
    h_7 = 'b00000001100110010110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111111010111110100;
    x_1 = 'b11111101111001100000;
    x_2 = 'b11111100010011101101;
    x_3 = 'b11111011001101000000;
    x_4 = 'b11111011000101110100;
    x_5 = 'b11111010011111111100;
    x_6 = 'b11111100101111011010;
    x_7 = 'b00000000111101101001;
    x_8 = 'b11111100011110101110;
    x_9 = 'b11111100111110011010;
    x_10 = 'b11111100110011000110;
    x_11 = 'b11111010101110110101;
    x_12 = 'b11111011011000110000;
    x_13 = 'b11111011100011110111;
    x_14 = 'b11111101100111100110;
    x_15 = 'b11111101000110011111;

    h_0 = 'b11111111010111110100;
    h_1 = 'b11111101111001100000;
    h_2 = 'b11111100010011101101;
    h_3 = 'b11111011001101000000;
    h_4 = 'b11111011000101110100;
    h_5 = 'b11111010011111111100;
    h_6 = 'b11111100101111011010;
    h_7 = 'b00000000111101101001;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111111001101111101;
    x_1 = 'b11111101100001000010;
    x_2 = 'b11111011011110010011;
    x_3 = 'b11111010000100011111;
    x_4 = 'b11111010000100001001;
    x_5 = 'b11111001101000011101;
    x_6 = 'b11111011101010111101;
    x_7 = 'b00000000111000100011;
    x_8 = 'b11111100101110001100;
    x_9 = 'b11111100001100010011;
    x_10 = 'b11111011011111111011;
    x_11 = 'b11111001010011000110;
    x_12 = 'b11111010011110001110;
    x_13 = 'b11111001111101101010;
    x_14 = 'b11111111000001001111;
    x_15 = 'b11111101000001011010;

    h_0 = 'b11111111001101111101;
    h_1 = 'b11111101100001000010;
    h_2 = 'b11111011011110010011;
    h_3 = 'b11111010000100011111;
    h_4 = 'b11111010000100001001;
    h_5 = 'b11111001101000011101;
    h_6 = 'b11111011101010111101;
    h_7 = 'b00000000111000100011;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111110111010001110;
    x_1 = 'b11111100110100111111;
    x_2 = 'b11111010101101101111;
    x_3 = 'b11111001101100010100;
    x_4 = 'b11111001100101110101;
    x_5 = 'b11111001001100101110;
    x_6 = 'b11111010011010000011;
    x_7 = 'b00000000000101101001;
    x_8 = 'b11111011111111110001;
    x_9 = 'b11111011011010001100;
    x_10 = 'b11111011000010100101;
    x_11 = 'b11111001001000111010;
    x_12 = 'b11111010000000111101;
    x_13 = 'b11111000000011000000;
    x_14 = 'b11111110010001110010;
    x_15 = 'b11111100011000101110;

    h_0 = 'b11111110111010001110;
    h_1 = 'b11111100110100111111;
    h_2 = 'b11111010101101101111;
    h_3 = 'b11111001101100010100;
    h_4 = 'b11111001100101110101;
    h_5 = 'b11111001001100101110;
    h_6 = 'b11111010011010000011;
    h_7 = 'b00000000000101101001;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111110110000010110;
    x_1 = 'b11111011111010010000;
    x_2 = 'b11111001111101001100;
    x_3 = 'b11111000110111001001;
    x_4 = 'b11111001000010011101;
    x_5 = 'b11111001010010010001;
    x_6 = 'b11111011000101100111;
    x_7 = 'b00000000000000100100;
    x_8 = 'b11111011010001010111;
    x_9 = 'b11111011000001001000;
    x_10 = 'b11111010100101001110;
    x_11 = 'b11111001001000111010;
    x_12 = 'b11111010010010100000;
    x_13 = 'b11111001100010011001;
    x_14 = 'b11111110000111001111;
    x_15 = 'b11111100100010111001;

    h_0 = 'b11111110110000010110;
    h_1 = 'b11111011111010010000;
    h_2 = 'b11111001111101001100;
    h_3 = 'b11111000110111001001;
    h_4 = 'b11111001000010011101;
    h_5 = 'b11111001010010010001;
    h_6 = 'b11111011000101100111;
    h_7 = 'b00000000000000100100;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111101110101001010;
    x_1 = 'b11111011011000000000;
    x_2 = 'b11111001100100111010;
    x_3 = 'b11111000011010001001;
    x_4 = 'b11111001000010011101;
    x_5 = 'b11111001000111001011;
    x_6 = 'b11111010111111011001;
    x_7 = 'b11111111010111110110;
    x_8 = 'b11111011001100001100;
    x_9 = 'b11111011000001001000;
    x_10 = 'b11111010111000110011;
    x_11 = 'b11111001011000001100;
    x_12 = 'b11111010101001111011;
    x_13 = 'b11111001111101101010;
    x_14 = 'b11111101111100101100;
    x_15 = 'b11111100111100010100;

    h_0 = 'b11111101110101001010;
    h_1 = 'b11111011011000000000;
    h_2 = 'b11111001100100111010;
    h_3 = 'b11111000011010001001;
    h_4 = 'b11111001000010011101;
    h_5 = 'b11111001000111001011;
    h_6 = 'b11111010111111011001;
    h_7 = 'b11111111010111110110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111101110000001110;
    x_1 = 'b11111011111111001001;
    x_2 = 'b11111001101001110001;
    x_3 = 'b11111000010101010100;
    x_4 = 'b11111000110011010011;
    x_5 = 'b11111000101011011100;
    x_6 = 'b11111001101000010000;
    x_7 = 'b11111111010010110000;
    x_8 = 'b11111011110101011101;
    x_9 = 'b11111011010101001011;
    x_10 = 'b11111011001100010111;
    x_11 = 'b11111001110001101011;
    x_12 = 'b11111010011000010111;
    x_13 = 'b11111000100101000100;
    x_14 = 'b11111110011100010101;
    x_15 = 'b11111101011111111011;

    h_0 = 'b11111101110000001110;
    h_1 = 'b11111011111111001001;
    h_2 = 'b11111001101001110001;
    h_3 = 'b11111000010101010100;
    h_4 = 'b11111000110011010011;
    h_5 = 'b11111000101011011100;
    h_6 = 'b11111001101000010000;
    h_7 = 'b11111111010010110000;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111111101011100011;
    x_1 = 'b11111101111110011010;
    x_2 = 'b11111011001111101111;
    x_3 = 'b11111001110101111111;
    x_4 = 'b11111001011011101110;
    x_5 = 'b11111001000111001011;
    x_6 = 'b11111010010011110100;
    x_7 = 'b00000001000010101110;
    x_8 = 'b11111101001101001000;
    x_9 = 'b11111100010001010100;
    x_10 = 'b11111011111000011001;
    x_11 = 'b11111010001011001010;
    x_12 = 'b11111011000111001100;
    x_13 = 'b11111001110110110101;
    x_14 = 'b00000000000000100010;
    x_15 = 'b11111110000011100001;

    h_0 = 'b11111111101011100011;
    h_1 = 'b11111101111110011010;
    h_2 = 'b11111011001111101111;
    h_3 = 'b11111001110101111111;
    h_4 = 'b11111001011011101110;
    h_5 = 'b11111001000111001011;
    h_6 = 'b11111010010011110100;
    h_7 = 'b00000001000010101110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111111100110100111;
    x_1 = 'b11111101010111010000;
    x_2 = 'b11111010110111011101;
    x_3 = 'b11111001001111010100;
    x_4 = 'b11111000101001001101;
    x_5 = 'b11111000001111101101;
    x_6 = 'b11111001000010111010;
    x_7 = 'b00000000110011011101;
    x_8 = 'b11111100101110001100;
    x_9 = 'b11111011111101010001;
    x_10 = 'b11111011111000011001;
    x_11 = 'b11111001100111011111;
    x_12 = 'b11111010111011011111;
    x_13 = 'b11111001111101101010;
    x_14 = 'b00000000000101110011;
    x_15 = 'b11111101101010000101;

    h_0 = 'b11111111100110100111;
    h_1 = 'b11111101010111010000;
    h_2 = 'b11111010110111011101;
    h_3 = 'b11111001001111010100;
    h_4 = 'b11111000101001001101;
    h_5 = 'b11111000001111101101;
    h_6 = 'b11111001000010111010;
    h_7 = 'b00000000110011011101;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000000100110101111;
    x_1 = 'b11111110010001111111;
    x_2 = 'b11111011011110010011;
    x_3 = 'b11111000101101011110;
    x_4 = 'b11111000011111000110;
    x_5 = 'b11111000001111101101;
    x_6 = 'b11111001110100101101;
    x_7 = 'b00000010101000100001;
    x_8 = 'b11111110011010011111;
    x_9 = 'b11111101100110100000;
    x_10 = 'b11111101010000011101;
    x_11 = 'b11111010011111100010;
    x_12 = 'b11111011011000110000;
    x_13 = 'b11111011101010101011;
    x_14 = 'b00000010011001011101;
    x_15 = 'b00000000001100110100;

    h_0 = 'b00000000100110101111;
    h_1 = 'b11111110010001111111;
    h_2 = 'b11111011011110010011;
    h_3 = 'b11111000101101011110;
    h_4 = 'b11111000011111000110;
    h_5 = 'b11111000001111101101;
    h_6 = 'b11111001110100101101;
    h_7 = 'b00000010101000100001;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000000000100001101;
    x_1 = 'b11111110110100001111;
    x_2 = 'b11111100000101001001;
    x_3 = 'b11111001010100001001;
    x_4 = 'b11111000000101110101;
    x_5 = 'b11110111001101001001;
    x_6 = 'b11111001001111010111;
    x_7 = 'b00000010100011011011;
    x_8 = 'b11111110101001111101;
    x_9 = 'b11111110010011100110;
    x_10 = 'b11111101010101010110;
    x_11 = 'b11111001100010011001;
    x_12 = 'b11111001010111111110;
    x_13 = 'b11111001111101101010;
    x_14 = 'b00000011011110000001;
    x_15 = 'b00000000101011010101;

    h_0 = 'b00000000000100001101;
    h_1 = 'b11111110110100001111;
    h_2 = 'b11111100000101001001;
    h_3 = 'b11111001010100001001;
    h_4 = 'b11111000000101110101;
    h_5 = 'b11110111001101001001;
    h_6 = 'b11111001001111010111;
    h_7 = 'b00000010100011011011;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000000111010011110;
    x_1 = 'b11111111010110100000;
    x_2 = 'b11111100011101011011;
    x_3 = 'b11111001110101111111;
    x_4 = 'b11111000111000010111;
    x_5 = 'b11110111101000111000;
    x_6 = 'b11111001011011110100;
    x_7 = 'b00000010110111110010;
    x_8 = 'b11111110101111000111;
    x_9 = 'b11111110000100100100;
    x_10 = 'b11111100101001010100;
    x_11 = 'b11111001100010011001;
    x_12 = 'b11111000110100110111;
    x_13 = 'b11111001111101101010;
    x_14 = 'b00000010111001000110;
    x_15 = 'b00000000010110111111;

    h_0 = 'b00000000111010011110;
    h_1 = 'b11111111010110100000;
    h_2 = 'b11111100011101011011;
    h_3 = 'b11111001110101111111;
    h_4 = 'b11111000111000010111;
    h_5 = 'b11110111101000111000;
    h_6 = 'b11111001011011110100;
    h_7 = 'b00000010110111110010;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111001001101001100;
    x_1 = 'b11111011110000011110;
    x_2 = 'b11111100001010000000;
    x_3 = 'b11111110100110100010;
    x_4 = 'b11111111000111011110;
    x_5 = 'b11111111000000011000;
    x_6 = 'b11111101000010000101;
    x_7 = 'b11111011011001010111;
    x_8 = 'b11111101100001110000;
    x_9 = 'b11111110011000100111;
    x_10 = 'b11111111011001011100;
    x_11 = 'b11111111111111001010;
    x_12 = 'b00000000011010101011;
    x_13 = 'b11111111001011100011;
    x_14 = 'b11111101100010010100;
    x_15 = 'b11111110100010000010;

    h_0 = 'b11111001001101001100;
    h_1 = 'b11111011110000011110;
    h_2 = 'b11111100001010000000;
    h_3 = 'b11111110100110100010;
    h_4 = 'b11111111000111011110;
    h_5 = 'b11111111000000011000;
    h_6 = 'b11111101000010000101;
    h_7 = 'b11111011011001010111;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111001101111101110;
    x_1 = 'b11111100100001011010;
    x_2 = 'b11111100111010100100;
    x_3 = 'b11111110101011010111;
    x_4 = 'b11111111010110101000;
    x_5 = 'b11111111110010010011;
    x_6 = 'b11111110111110100011;
    x_7 = 'b11111100010001010110;
    x_8 = 'b11111110001011000001;
    x_9 = 'b11111110100010101000;
    x_10 = 'b11111110101101011010;
    x_11 = 'b11111111111010000100;
    x_12 = 'b00000000100110011000;
    x_13 = 'b00000000101010111101;
    x_14 = 'b11111101010111110001;
    x_15 = 'b11111110010111110111;

    h_0 = 'b11111001101111101110;
    h_1 = 'b11111100100001011010;
    h_2 = 'b11111100111010100100;
    h_3 = 'b11111110101011010111;
    h_4 = 'b11111111010110101000;
    h_5 = 'b11111111110010010011;
    h_6 = 'b11111110111110100011;
    h_7 = 'b11111100010001010110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111010100101111111;
    x_1 = 'b11111101010111010000;
    x_2 = 'b11111101010111101100;
    x_3 = 'b11111110100001101101;
    x_4 = 'b11111111000111011110;
    x_5 = 'b11111111110010010011;
    x_6 = 'b00000000000011000001;
    x_7 = 'b11111101011000100110;
    x_8 = 'b11111110110100010001;
    x_9 = 'b11111110001110100110;
    x_10 = 'b11111101110111100110;
    x_11 = 'b11111111000010000000;
    x_12 = 'b00000000001110111110;
    x_13 = 'b00000001010011110101;
    x_14 = 'b11111101111100101100;
    x_15 = 'b11111110111011011101;

    h_0 = 'b11111010100101111111;
    h_1 = 'b11111101010111010000;
    h_2 = 'b11111101010111101100;
    h_3 = 'b11111110100001101101;
    h_4 = 'b11111111000111011110;
    h_5 = 'b11111111110010010011;
    h_6 = 'b00000000000011000001;
    h_7 = 'b11111101011000100110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111100001101100100;
    x_1 = 'b11111110010001111111;
    x_2 = 'b11111101111001101100;
    x_3 = 'b11111110100110100010;
    x_4 = 'b11111110111101010111;
    x_5 = 'b11111111010001000001;
    x_6 = 'b11111110111110100011;
    x_7 = 'b11111110101010000010;
    x_8 = 'b11111111011000011000;
    x_9 = 'b11111110100111101001;
    x_10 = 'b11111110011110101111;
    x_11 = 'b11111110011110010101;
    x_12 = 'b11111110111101000001;
    x_13 = 'b11111110010101000010;
    x_14 = 'b11111111000110100001;
    x_15 = 'b11111111001111110011;

    h_0 = 'b11111100001101100100;
    h_1 = 'b11111110010001111111;
    h_2 = 'b11111101111001101100;
    h_3 = 'b11111110100110100010;
    h_4 = 'b11111110111101010111;
    h_5 = 'b11111111010001000001;
    h_6 = 'b11111110111110100011;
    h_7 = 'b11111110101010000010;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111011111001110110;
    x_1 = 'b11111101111001100000;
    x_2 = 'b11111101101111111110;
    x_3 = 'b11111110100110100010;
    x_4 = 'b11111110111000010100;
    x_5 = 'b11111110111010110101;
    x_6 = 'b11111101101101101001;
    x_7 = 'b11111101100010110010;
    x_8 = 'b11111110111001011100;
    x_9 = 'b11111110110110101011;
    x_10 = 'b11111111001010110001;
    x_11 = 'b11111111100000100101;
    x_12 = 'b11111110110001010100;
    x_13 = 'b11111101111001110010;
    x_14 = 'b11111101001101001110;
    x_15 = 'b11111110010111110111;

    h_0 = 'b11111011111001110110;
    h_1 = 'b11111101111001100000;
    h_2 = 'b11111101101111111110;
    h_3 = 'b11111110100110100010;
    h_4 = 'b11111110111000010100;
    h_5 = 'b11111110111010110101;
    h_6 = 'b11111101101101101001;
    h_7 = 'b11111101100010110010;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111011111110110001;
    x_1 = 'b11111110000011010011;
    x_2 = 'b11111110100000100010;
    x_3 = 'b11111111110011111000;
    x_4 = 'b00000000010011010000;
    x_5 = 'b00000000011110101011;
    x_6 = 'b11111111101010000111;
    x_7 = 'b11111110010000100101;
    x_8 = 'b11111111100010101100;
    x_9 = 'b11111111101101110011;
    x_10 = 'b00000000000000100101;
    x_11 = 'b00000000100010110101;
    x_12 = 'b00000000111101110010;
    x_13 = 'b00000000100100001001;
    x_14 = 'b11111100111101011010;
    x_15 = 'b11111110101100001101;

    h_0 = 'b11111011111110110001;
    h_1 = 'b11111110000011010011;
    h_2 = 'b11111110100000100010;
    h_3 = 'b11111111110011111000;
    h_4 = 'b00000000010011010000;
    h_5 = 'b00000000011110101011;
    h_6 = 'b11111111101010000111;
    h_7 = 'b11111110010000100101;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111010001000011001;
    x_1 = 'b11111100011100100001;
    x_2 = 'b11111100110101101101;
    x_3 = 'b11111110110101000010;
    x_4 = 'b11111111011011101011;
    x_5 = 'b11111111011100000111;
    x_6 = 'b11111110001100110001;
    x_7 = 'b11111011110111111001;
    x_8 = 'b11111101110001001111;
    x_9 = 'b11111101110101100010;
    x_10 = 'b11111110011110101111;
    x_11 = 'b11111111110100111101;
    x_12 = 'b00000000100110011000;
    x_13 = 'b11111111000100101111;
    x_14 = 'b11111011111000110110;
    x_15 = 'b11111100111100010100;

    h_0 = 'b11111010001000011001;
    h_1 = 'b11111100011100100001;
    h_2 = 'b11111100110101101101;
    h_3 = 'b11111110110101000010;
    h_4 = 'b11111111011011101011;
    h_5 = 'b11111111011100000111;
    h_6 = 'b11111110001100110001;
    h_7 = 'b11111011110111111001;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111010101010111011;
    x_1 = 'b11111101001101011101;
    x_2 = 'b11111101001101111111;
    x_3 = 'b11111111010110111000;
    x_4 = 'b00000000011101010110;
    x_5 = 'b00000001000101100000;
    x_6 = 'b11111111010001001110;
    x_7 = 'b11111101011000100110;
    x_8 = 'b11111110010000001011;
    x_9 = 'b11111110011101101000;
    x_10 = 'b11111111011110010101;
    x_11 = 'b00000001010101110010;
    x_12 = 'b00000010011011011100;
    x_13 = 'b00000001000110001101;
    x_14 = 'b11111100111101011010;
    x_15 = 'b11111101010101110000;

    h_0 = 'b11111010101010111011;
    h_1 = 'b11111101001101011101;
    h_2 = 'b11111101001101111111;
    h_3 = 'b11111111010110111000;
    h_4 = 'b00000000011101010110;
    h_5 = 'b00000001000101100000;
    h_6 = 'b11111111010001001110;
    h_7 = 'b11111101011000100110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111100011100011000;
    x_1 = 'b11111110001101000101;
    x_2 = 'b11111110000011011001;
    x_3 = 'b00000000000010011000;
    x_4 = 'b00000000110001100100;
    x_5 = 'b00000000111010011010;
    x_6 = 'b11111111011101101011;
    x_7 = 'b11111101101100111101;
    x_8 = 'b11111110010000001011;
    x_9 = 'b11111110110110101011;
    x_10 = 'b11111111110110110011;
    x_11 = 'b00000001000110100000;
    x_12 = 'b00000001101100100111;
    x_13 = 'b00000000001000111000;
    x_14 = 'b11111100001000101011;
    x_15 = 'b11111101010000101010;

    h_0 = 'b11111100011100011000;
    h_1 = 'b11111110001101000101;
    h_2 = 'b11111110000011011001;
    h_3 = 'b00000000000010011000;
    h_4 = 'b00000000110001100100;
    h_5 = 'b00000000111010011010;
    h_6 = 'b11111111011101101011;
    h_7 = 'b11111101101100111101;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111100110101000010;
    x_1 = 'b11111110111110000010;
    x_2 = 'b11111110011011101011;
    x_3 = 'b00000000010000111000;
    x_4 = 'b00000000010011010000;
    x_5 = 'b00000000001000011111;
    x_6 = 'b11111110111110100011;
    x_7 = 'b11111110011010110001;
    x_8 = 'b11111110111001011100;
    x_9 = 'b11111111011110110001;
    x_10 = 'b00000000001111010001;
    x_11 = 'b00000001000110100000;
    x_12 = 'b00000001001001100000;
    x_13 = 'b11111111110100011100;
    x_14 = 'b11111101011101000011;
    x_15 = 'b11111110100010000010;

    h_0 = 'b11111100110101000010;
    h_1 = 'b11111110111110000010;
    h_2 = 'b11111110011011101011;
    h_3 = 'b00000000010000111000;
    h_4 = 'b00000000010011010000;
    h_5 = 'b00000000001000011111;
    h_6 = 'b11111110111110100011;
    h_7 = 'b11111110011010110001;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111100100001010011;
    x_1 = 'b11111111010001100111;
    x_2 = 'b11111110100000100010;
    x_3 = 'b00000000001100000011;
    x_4 = 'b00000000001001001001;
    x_5 = 'b00000000011110101011;
    x_6 = 'b11111111010001001110;
    x_7 = 'b11111111011100111100;
    x_8 = 'b00000000000001101000;
    x_9 = 'b11111111110010110100;
    x_10 = 'b11111111110110110011;
    x_11 = 'b00000001000110100000;
    x_12 = 'b00000000110010000101;
    x_13 = 'b00000000001000111000;
    x_14 = 'b11111110111011111110;
    x_15 = 'b11111111100100001001;

    h_0 = 'b11111100100001010011;
    h_1 = 'b11111111010001100111;
    h_2 = 'b11111110100000100010;
    h_3 = 'b00000000001100000011;
    h_4 = 'b00000000001001001001;
    h_5 = 'b00000000011110101011;
    h_6 = 'b11111111010001001110;
    h_7 = 'b11111111011100111100;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111011101011000011;
    x_1 = 'b11111100111110110010;
    x_2 = 'b11111100110101101101;
    x_3 = 'b11111110111001110111;
    x_4 = 'b11111110101110001101;
    x_5 = 'b11111110010100000000;
    x_6 = 'b11111101010100110000;
    x_7 = 'b11111101100010110010;
    x_8 = 'b11111110000101110111;
    x_9 = 'b11111101110000100001;
    x_10 = 'b11111101110111100110;
    x_11 = 'b11111111010001010010;
    x_12 = 'b11111110011001111001;
    x_13 = 'b11111101001010000101;
    x_14 = 'b11111101110010001001;
    x_15 = 'b11111101111110011011;

    h_0 = 'b11111011101011000011;
    h_1 = 'b11111100111110110010;
    h_2 = 'b11111100110101101101;
    h_3 = 'b11111110111001110111;
    h_4 = 'b11111110101110001101;
    h_5 = 'b11111110010100000000;
    h_6 = 'b11111101010100110000;
    h_7 = 'b11111101100010110010;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111110001000111001;
    x_1 = 'b11111111010110100000;
    x_2 = 'b11111111000010100001;
    x_3 = 'b00000000110111100011;
    x_4 = 'b00000000110001100100;
    x_5 = 'b00000000001000011111;
    x_6 = 'b11111110101011111000;
    x_7 = 'b00000001010111000101;
    x_8 = 'b00000000110000000011;
    x_9 = 'b00000000000001110110;
    x_10 = 'b00000000001010011000;
    x_11 = 'b00000001101010001011;
    x_12 = 'b00000000100000100001;
    x_13 = 'b11111111001011100011;
    x_14 = 'b00000000010101101000;
    x_15 = 'b00000000100110010000;

    h_0 = 'b11111110001000111001;
    h_1 = 'b11111111010110100000;
    h_2 = 'b11111111000010100001;
    h_3 = 'b00000000110111100011;
    h_4 = 'b00000000110001100100;
    h_5 = 'b00000000001000011111;
    h_6 = 'b11111110101011111000;
    h_7 = 'b00000001010111000101;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111110100110011111;
    x_1 = 'b11111111010110100000;
    x_2 = 'b11111110100000100010;
    x_3 = 'b11111111111000101101;
    x_4 = 'b11111111100101110010;
    x_5 = 'b11111111001011011110;
    x_6 = 'b11111101110011110111;
    x_7 = 'b00000000011111000110;
    x_8 = 'b11111111110111010100;
    x_9 = 'b11111111000101101101;
    x_10 = 'b11111110110111001101;
    x_11 = 'b11111111101010110001;
    x_12 = 'b11111110001000010110;
    x_13 = 'b11111101001010000101;
    x_14 = 'b11111110100001100110;
    x_15 = 'b11111111000000100010;

    h_0 = 'b11111110100110011111;
    h_1 = 'b11111111010110100000;
    h_2 = 'b11111110100000100010;
    h_3 = 'b11111111111000101101;
    h_4 = 'b11111111100101110010;
    h_5 = 'b11111111001011011110;
    h_6 = 'b11111101110011110111;
    h_7 = 'b00000000011111000110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111101001000110001;
    x_1 = 'b11111110010001111111;
    x_2 = 'b11111101100110010001;
    x_3 = 'b11111110100001101101;
    x_4 = 'b11111110101001001010;
    x_5 = 'b11111110011001100011;
    x_6 = 'b11111101110011110111;
    x_7 = 'b11111101111100001111;
    x_8 = 'b11111110000101110111;
    x_9 = 'b11111101111010100011;
    x_10 = 'b11111101101000111011;
    x_11 = 'b11111110110111110100;
    x_12 = 'b11111101011111010111;
    x_13 = 'b11111101001010000101;
    x_14 = 'b11111100111000001000;
    x_15 = 'b11111101001011100101;

    h_0 = 'b11111101001000110001;
    h_1 = 'b11111110010001111111;
    h_2 = 'b11111101100110010001;
    h_3 = 'b11111110100001101101;
    h_4 = 'b11111110101001001010;
    h_5 = 'b11111110011001100011;
    h_6 = 'b11111101110011110111;
    h_7 = 'b11111101111100001111;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111101010111100100;
    x_1 = 'b11111110101111010110;
    x_2 = 'b11111110100000100010;
    x_3 = 'b11111111101010001101;
    x_4 = 'b11111111110100111100;
    x_5 = 'b00000000000010111100;
    x_6 = 'b11111110101011111000;
    x_7 = 'b11111110111110011001;
    x_8 = 'b11111110100100110011;
    x_9 = 'b11111110100010101000;
    x_10 = 'b11111110101000100001;
    x_11 = 'b00000000001001010110;
    x_12 = 'b11111111010100011011;
    x_13 = 'b11111110111101111011;
    x_14 = 'b11111101010111110001;
    x_15 = 'b11111101100101000000;

    h_0 = 'b11111101010111100100;
    h_1 = 'b11111110101111010110;
    h_2 = 'b11111110100000100010;
    h_3 = 'b11111111101010001101;
    h_4 = 'b11111111110100111100;
    h_5 = 'b00000000000010111100;
    h_6 = 'b11111110101011111000;
    h_7 = 'b11111110111110011001;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000001110000101111;
    x_1 = 'b00000001110011000111;
    x_2 = 'b00000000101101010110;
    x_3 = 'b00000001100011000100;
    x_4 = 'b00000001111101010110;
    x_5 = 'b00000000111010011010;
    x_6 = 'b00000000111011000001;
    x_7 = 'b00000000011010000000;
    x_8 = 'b00000001001110111111;
    x_9 = 'b00000001100001000011;
    x_10 = 'b00000010001001100101;
    x_11 = 'b00000000001110011100;
    x_12 = 'b00000001011011000011;
    x_13 = 'b00000010000011100010;
    x_14 = 'b00000001011010001011;
    x_15 = 'b00000001011110001100;

    h_0 = 'b00000001110000101111;
    h_1 = 'b00000001110011000111;
    h_2 = 'b00000000101101010110;
    h_3 = 'b00000001100011000100;
    h_4 = 'b00000001111101010110;
    h_5 = 'b00000000111010011010;
    h_6 = 'b00000000111011000001;
    h_7 = 'b00000000011010000000;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000000100110101111;
    x_1 = 'b00000000110011011111;
    x_2 = 'b00000000000110100000;
    x_3 = 'b00000001001111101110;
    x_4 = 'b00000001100100000101;
    x_5 = 'b00000000000010111100;
    x_6 = 'b11111111110000010110;
    x_7 = 'b11111111010111110110;
    x_8 = 'b00000000011011011011;
    x_9 = 'b00000001001000000000;
    x_10 = 'b00000001100111010101;
    x_11 = 'b00000000011000101000;
    x_12 = 'b00000000110010000101;
    x_13 = 'b00000000111000100101;
    x_14 = 'b00000000101111111111;
    x_15 = 'b00000000011100000101;

    h_0 = 'b00000000100110101111;
    h_1 = 'b00000000110011011111;
    h_2 = 'b00000000000110100000;
    h_3 = 'b00000001001111101110;
    h_4 = 'b00000001100100000101;
    h_5 = 'b00000000000010111100;
    h_6 = 'b11111111110000010110;
    h_7 = 'b11111111010111110110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111111010111110100;
    x_1 = 'b00000000000010100011;
    x_2 = 'b00000000000001101001;
    x_3 = 'b00000001100011000100;
    x_4 = 'b00000001101110001100;
    x_5 = 'b00000000000010111100;
    x_6 = 'b11111111010001001110;
    x_7 = 'b11111101110111001001;
    x_8 = 'b11111111001110000100;
    x_9 = 'b00000000101001111100;
    x_10 = 'b00000001111010111001;
    x_11 = 'b11111111111111001010;
    x_12 = 'b00000000011010101011;
    x_13 = 'b00000000110001110001;
    x_14 = 'b11111110110110101100;
    x_15 = 'b11111111110011011001;

    h_0 = 'b11111111010111110100;
    h_1 = 'b00000000000010100011;
    h_2 = 'b00000000000001101001;
    h_3 = 'b00000001100011000100;
    h_4 = 'b00000001101110001100;
    h_5 = 'b00000000000010111100;
    h_6 = 'b11111111010001001110;
    h_7 = 'b11111101110111001001;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111101101011010011;
    x_1 = 'b11111110011011110001;
    x_2 = 'b11111110001101000111;
    x_3 = 'b11111111100000100011;
    x_4 = 'b11111111101111111000;
    x_5 = 'b11111110000011010111;
    x_6 = 'b11111101001000010011;
    x_7 = 'b11111100000111001011;
    x_8 = 'b11111110000000101101;
    x_9 = 'b11111111001111101111;
    x_10 = 'b00000000011101111100;
    x_11 = 'b11111101110000011110;
    x_12 = 'b11111110100101100111;
    x_13 = 'b11111111101101101000;
    x_14 = 'b11111110110110101100;
    x_15 = 'b11111111100100001001;

    h_0 = 'b11111101101011010011;
    h_1 = 'b11111110011011110001;
    h_2 = 'b11111110001101000111;
    h_3 = 'b11111111100000100011;
    h_4 = 'b11111111101111111000;
    h_5 = 'b11111110000011010111;
    h_6 = 'b11111101001000010011;
    h_7 = 'b11111100000111001011;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111110100110011111;
    x_1 = 'b11111111001100101101;
    x_2 = 'b11111110000011011001;
    x_3 = 'b11111110110000001101;
    x_4 = 'b11111110110011010000;
    x_5 = 'b11111101010110111111;
    x_6 = 'b11111101010100110000;
    x_7 = 'b11111101011101101100;
    x_8 = 'b11111110100100110011;
    x_9 = 'b11111110111011101100;
    x_10 = 'b11111111011110010101;
    x_11 = 'b11111101000010100111;
    x_12 = 'b11111101011001100001;
    x_13 = 'b11111111001011100011;
    x_14 = 'b11111111010110010110;
    x_15 = 'b11111111101001001110;

    h_0 = 'b11111110100110011111;
    h_1 = 'b11111111001100101101;
    h_2 = 'b11111110000011011001;
    h_3 = 'b11111110110000001101;
    h_4 = 'b11111110110011010000;
    h_5 = 'b11111101010110111111;
    h_6 = 'b11111101010100110000;
    h_7 = 'b11111101011101101100;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111110100110011111;
    x_1 = 'b11111111010001100111;
    x_2 = 'b11111110010110110100;
    x_3 = 'b11111110101011010111;
    x_4 = 'b11111111001100100001;
    x_5 = 'b11111110000011010111;
    x_6 = 'b11111101100111011011;
    x_7 = 'b11111110010101101011;
    x_8 = 'b11111111010011001110;
    x_9 = 'b11111111011110110001;
    x_10 = 'b11111111101101000001;
    x_11 = 'b11111101100110010010;
    x_12 = 'b11111101111100101000;
    x_13 = 'b11111111001011100011;
    x_14 = 'b00000000010000010110;
    x_15 = 'b00000000011100000101;

    h_0 = 'b11111110100110011111;
    h_1 = 'b11111111010001100111;
    h_2 = 'b11111110010110110100;
    h_3 = 'b11111110101011010111;
    h_4 = 'b11111111001100100001;
    h_5 = 'b11111110000011010111;
    h_6 = 'b11111101100111011011;
    h_7 = 'b11111110010101101011;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000000001001001001;
    x_1 = 'b00000000010110001000;
    x_2 = 'b11111111010001000101;
    x_3 = 'b11111111010110111000;
    x_4 = 'b00000000001110001100;
    x_5 = 'b11111111101100110000;
    x_6 = 'b11111111110110100100;
    x_7 = 'b11111111010111110110;
    x_8 = 'b00000000000001101000;
    x_9 = 'b00000000010000111000;
    x_10 = 'b00000000100010110101;
    x_11 = 'b11111110011110010101;
    x_12 = 'b11111111110111100011;
    x_13 = 'b00000001000110001101;
    x_14 = 'b00000001001010010111;
    x_15 = 'b00000000110101100000;

    h_0 = 'b00000000001001001001;
    h_1 = 'b00000000010110001000;
    h_2 = 'b11111111010001000101;
    h_3 = 'b11111111010110111000;
    h_4 = 'b00000000001110001100;
    h_5 = 'b11111111101100110000;
    h_6 = 'b11111111110110100100;
    h_7 = 'b11111111010111110110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000000111111011010;
    x_1 = 'b00000001000010001011;
    x_2 = 'b11111111110111111100;
    x_3 = 'b11111111111101100011;
    x_4 = 'b00000000100010011010;
    x_5 = 'b00000000000010111100;
    x_6 = 'b00000000000011000001;
    x_7 = 'b00000000011111000110;
    x_8 = 'b00000000111010010111;
    x_9 = 'b00000001001101000001;
    x_10 = 'b00000010000100101011;
    x_11 = 'b11111111010110011001;
    x_12 = 'b00000000110111111100;
    x_13 = 'b00000001101111000110;
    x_14 = 'b00000010100100000000;
    x_15 = 'b00000001111100101101;

    h_0 = 'b00000000111111011010;
    h_1 = 'b00000001000010001011;
    h_2 = 'b11111111110111111100;
    h_3 = 'b11111111111101100011;
    h_4 = 'b00000000100010011010;
    h_5 = 'b00000000000010111100;
    h_6 = 'b00000000000011000001;
    h_7 = 'b00000000011111000110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000001011000000100;
    x_1 = 'b00000001000111000100;
    x_2 = 'b00000000001011010111;
    x_3 = 'b00000000101101111001;
    x_4 = 'b00000001001010110100;
    x_5 = 'b11111111111101011001;
    x_6 = 'b11111110100101101010;
    x_7 = 'b00000001000010101110;
    x_8 = 'b00000000110101001101;
    x_9 = 'b00000001011100000011;
    x_10 = 'b00000010101011110100;
    x_11 = 'b11111111111111001010;
    x_12 = 'b00000001010101001101;
    x_13 = 'b00000001110101111010;
    x_14 = 'b00000010110011110101;
    x_15 = 'b00000001110111100111;

    h_0 = 'b00000001011000000100;
    h_1 = 'b00000001000111000100;
    h_2 = 'b00000000001011010111;
    h_3 = 'b00000000101101111001;
    h_4 = 'b00000001001010110100;
    h_5 = 'b11111111111101011001;
    h_6 = 'b11111110100101101010;
    h_7 = 'b00000001000010101110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000001110000101111;
    x_1 = 'b00000001101110001110;
    x_2 = 'b00000001001010011111;
    x_3 = 'b00000001111011001111;
    x_4 = 'b00000010100101110000;
    x_5 = 'b00000001011011101101;
    x_6 = 'b00000000000011000001;
    x_7 = 'b00000000000000100100;
    x_8 = 'b00000000100101101111;
    x_9 = 'b00000001111010000111;
    x_10 = 'b00000011011100101111;
    x_11 = 'b00000001100101000100;
    x_12 = 'b00000001110010011110;
    x_13 = 'b00000001101111000110;
    x_14 = 'b00000000100000001011;
    x_15 = 'b00000000111010100110;

    h_0 = 'b00000001110000101111;
    h_1 = 'b00000001101110001110;
    h_2 = 'b00000001001010011111;
    h_3 = 'b00000001111011001111;
    h_4 = 'b00000010100101110000;
    h_5 = 'b00000001011011101101;
    h_6 = 'b00000000000011000001;
    h_7 = 'b00000000000000100100;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000001000100010101;
    x_1 = 'b00000010010000011111;
    x_2 = 'b00000010101011100110;
    x_3 = 'b00000011100101100101;
    x_4 = 'b00000011100111011011;
    x_5 = 'b00000010001000000101;
    x_6 = 'b00000001011010001001;
    x_7 = 'b00000000000000100100;
    x_8 = 'b00000000111111100001;
    x_9 = 'b00000011000000010001;
    x_10 = 'b00000100101111111010;
    x_11 = 'b00000001111001011101;
    x_12 = 'b00000001100000111010;
    x_13 = 'b00000001010011110101;
    x_14 = 'b11111111010110010110;
    x_15 = 'b00000000111111101011;

    h_0 = 'b00000001000100010101;
    h_1 = 'b00000010010000011111;
    h_2 = 'b00000010101011100110;
    h_3 = 'b00000011100101100101;
    h_4 = 'b00000011100111011011;
    h_5 = 'b00000010001000000101;
    h_6 = 'b00000001011010001001;
    h_7 = 'b00000000000000100100;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000001110000101111;
    x_1 = 'b00000011010101000000;
    x_2 = 'b00000011110100011100;
    x_3 = 'b00000100100100011011;
    x_4 = 'b00000100001010110011;
    x_5 = 'b00000010011110010001;
    x_6 = 'b00000001011010001001;
    x_7 = 'b00000000001010101111;
    x_8 = 'b00000010101011110101;
    x_9 = 'b00000100101110100001;
    x_10 = 'b00000110001100111000;
    x_11 = 'b00000010011000000010;
    x_12 = 'b00000010000100000010;
    x_13 = 'b00000010101100011011;
    x_14 = 'b00000000110101010001;
    x_15 = 'b00000010101111100011;

    h_0 = 'b00000001110000101111;
    h_1 = 'b00000011010101000000;
    h_2 = 'b00000011110100011100;
    h_3 = 'b00000100100100011011;
    h_4 = 'b00000100001010110011;
    h_5 = 'b00000010011110010001;
    h_6 = 'b00000001011010001001;
    h_7 = 'b00000000001010101111;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000011010011011000;
    x_1 = 'b00000100101101000110;
    x_2 = 'b00000100111000011010;
    x_3 = 'b00000101011001100110;
    x_4 = 'b00000100111000010001;
    x_5 = 'b00000011011011010010;
    x_6 = 'b00000010010010001010;
    x_7 = 'b00000010101101100111;
    x_8 = 'b00000100110111000100;
    x_9 = 'b00000110101011110010;
    x_10 = 'b00001000001100000101;
    x_11 = 'b00000100110000111010;
    x_12 = 'b00000011100111100010;
    x_13 = 'b00000011100010111100;
    x_14 = 'b00000011111101101010;
    x_15 = 'b00000101101011101101;

    h_0 = 'b00000011010011011000;
    h_1 = 'b00000100101101000110;
    h_2 = 'b00000100111000011010;
    h_3 = 'b00000101011001100110;
    h_4 = 'b00000100111000010001;
    h_5 = 'b00000011011011010010;
    h_6 = 'b00000010010010001010;
    h_7 = 'b00000010101101100111;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000100100010010100;
    x_1 = 'b00000101111011011010;
    x_2 = 'b00000101110111100010;
    x_3 = 'b00000110000101000110;
    x_4 = 'b00000101101111110101;
    x_5 = 'b00000100001101001101;
    x_6 = 'b00000011000011111100;
    x_7 = 'b00000100001001001110;
    x_8 = 'b00000101111111010001;
    x_9 = 'b00000111000100110110;
    x_10 = 'b00001000000111001100;
    x_11 = 'b00000101101110000011;
    x_12 = 'b00000100111111010101;
    x_13 = 'b00000100110100101101;
    x_14 = 'b00000100111100111100;
    x_15 = 'b00000110001010001110;

    h_0 = 'b00000100100010010100;
    h_1 = 'b00000101111011011010;
    h_2 = 'b00000101110111100010;
    h_3 = 'b00000110000101000110;
    h_4 = 'b00000101101111110101;
    h_5 = 'b00000100001101001101;
    h_6 = 'b00000011000011111100;
    h_7 = 'b00000100001001001110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000010001110010101;
    x_1 = 'b00000011010000000111;
    x_2 = 'b00000010110000011101;
    x_3 = 'b00000010100110101111;
    x_4 = 'b00000010000111011100;
    x_5 = 'b00000000011001001000;
    x_6 = 'b11111110011111011100;
    x_7 = 'b00000001111010101101;
    x_8 = 'b00000011101001101101;
    x_9 = 'b00000011111100011010;
    x_10 = 'b00000100111001101101;
    x_11 = 'b00000010101100011010;
    x_12 = 'b00000010100001010011;
    x_13 = 'b00000001101000010010;
    x_14 = 'b00000010111110011000;
    x_15 = 'b00000100000110000000;

    h_0 = 'b00000010001110010101;
    h_1 = 'b00000011010000000111;
    h_2 = 'b00000010110000011101;
    h_3 = 'b00000010100110101111;
    h_4 = 'b00000010000111011100;
    h_5 = 'b00000000011001001000;
    h_6 = 'b11111110011111011100;
    h_7 = 'b00000001111010101101;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000001000100010101;
    x_1 = 'b00000001111100111010;
    x_2 = 'b00000001011001000011;
    x_3 = 'b00000001010100100100;
    x_4 = 'b00000000110001100100;
    x_5 = 'b11111111001011011110;
    x_6 = 'b11111101101101101001;
    x_7 = 'b00000001000111110100;
    x_8 = 'b00000010011100010110;
    x_9 = 'b00000011001111010011;
    x_10 = 'b00000100011100010110;
    x_11 = 'b00000010011000000010;
    x_12 = 'b00000010001111101111;
    x_13 = 'b00000001010011110101;
    x_14 = 'b00000010100100000000;
    x_15 = 'b00000011101100100101;

    h_0 = 'b00000001000100010101;
    h_1 = 'b00000001111100111010;
    h_2 = 'b00000001011001000011;
    h_3 = 'b00000001010100100100;
    h_4 = 'b00000000110001100100;
    h_5 = 'b11111111001011011110;
    h_6 = 'b11111101101101101001;
    h_7 = 'b00000001000111110100;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111111000100000101;
    x_1 = 'b11111111000111110100;
    x_2 = 'b11111101111001101100;
    x_3 = 'b11111110100110100010;
    x_4 = 'b11111110111101010111;
    x_5 = 'b11111110011111000110;
    x_6 = 'b11111111001011000000;
    x_7 = 'b11111111111011011110;
    x_8 = 'b11111110010000001011;
    x_9 = 'b11111101010111011110;
    x_10 = 'b11111101101101110100;
    x_11 = 'b11111101100110010010;
    x_12 = 'b11111110111101000001;
    x_13 = 'b00000000101010111101;
    x_14 = 'b11111110010001110010;
    x_15 = 'b11111110010111110111;

    h_0 = 'b11111111000100000101;
    h_1 = 'b11111111000111110100;
    h_2 = 'b11111101111001101100;
    h_3 = 'b11111110100110100010;
    h_4 = 'b11111110111101010111;
    h_5 = 'b11111110011111000110;
    h_6 = 'b11111111001011000000;
    h_7 = 'b11111111111011011110;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b00000000000100001101;
    x_1 = 'b11111111111101101010;
    x_2 = 'b11111110101010001111;
    x_3 = 'b11111111100101011000;
    x_4 = 'b11111111100000101110;
    x_5 = 'b11111110111010110101;
    x_6 = 'b11111111010001001110;
    x_7 = 'b00000000011010000000;
    x_8 = 'b11111110011111101001;
    x_9 = 'b11111101110000100001;
    x_10 = 'b11111110011001110110;
    x_11 = 'b11111110011001001111;
    x_12 = 'b11111111001110100101;
    x_13 = 'b00000001011010101010;
    x_14 = 'b11111110010111000011;
    x_15 = 'b11111110000011100001;

    h_0 = 'b00000000000100001101;
    h_1 = 'b11111111111101101010;
    h_2 = 'b11111110101010001111;
    h_3 = 'b11111111100101011000;
    h_4 = 'b11111111100000101110;
    h_5 = 'b11111110111010110101;
    h_6 = 'b11111111010001001110;
    h_7 = 'b00000000011010000000;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111110111010001110;
    x_1 = 'b11111110100101100100;
    x_2 = 'b11111101011100100011;
    x_3 = 'b11111110011100110111;
    x_4 = 'b11111110010100111100;
    x_5 = 'b11111101101101001011;
    x_6 = 'b11111101101101101001;
    x_7 = 'b11111110101010000010;
    x_8 = 'b11111100101001000010;
    x_9 = 'b11111100000010010010;
    x_10 = 'b11111100101110001101;
    x_11 = 'b11111100011110111100;
    x_12 = 'b11111100111100010000;
    x_13 = 'b11111110001110001110;
    x_14 = 'b11111100101101100101;
    x_15 = 'b11111011111010001101;

    h_0 = 'b11111110111010001110;
    h_1 = 'b11111110100101100100;
    h_2 = 'b11111101011100100011;
    h_3 = 'b11111110011100110111;
    h_4 = 'b11111110010100111100;
    h_5 = 'b11111101101101001011;
    h_6 = 'b11111101101101101001;
    h_7 = 'b11111110101010000010;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    x_0 = 'b11111110111010001110;
    x_1 = 'b11111110010001111111;
    x_2 = 'b11111100101011111111;
    x_3 = 'b11111101110110001100;
    x_4 = 'b11111101110110101000;
    x_5 = 'b11111101001011111001;
    x_6 = 'b11111101100001001101;
    x_7 = 'b11111111001000100101;
    x_8 = 'b11111011110101011101;
    x_9 = 'b11111011000001001000;
    x_10 = 'b11111011010110001001;
    x_11 = 'b11111011000011001101;
    x_12 = 'b11111011000111001100;
    x_13 = 'b11111100010011100100;
    x_14 = 'b11111100111000001000;
    x_15 = 'b11111011010110100111;

    h_0 = 'b11111110111010001110;
    h_1 = 'b11111110010001111111;
    h_2 = 'b11111100101011111111;
    h_3 = 'b11111101110110001100;
    h_4 = 'b11111101110110101000;
    h_5 = 'b11111101001011111001;
    h_6 = 'b11111101100001001101;
    h_7 = 'b11111111001000100101;
    #20;
    $fdisplay(fd, "%020b %020b %020b %020b %020b %020b %020b %020b", y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7);

    $fclose(fd);    
$finish;
    end
endmodule