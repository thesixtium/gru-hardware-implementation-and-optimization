`timescale 1ns / 1ps

module gru_tb;

// Parameters
parameter int INT_WIDTH  = 4;
parameter int FRAC_WIDTH = 5;
parameter int WIDTH      = INT_WIDTH + FRAC_WIDTH;
parameter real CLK_PERIOD = 10.0;

// Clock and reset
logic clk;
logic reset;

// Inputs
logic signed [WIDTH-1:0] x_0 = 0;
logic signed [WIDTH-1:0] x_1 = 0;
logic signed [WIDTH-1:0] x_2 = 0;
logic signed [WIDTH-1:0] x_3 = 0;
logic signed [WIDTH-1:0] x_4 = 0;

logic signed [WIDTH-1:0] h_0 = 0;
logic signed [WIDTH-1:0] h_1 = 0;
logic signed [WIDTH-1:0] h_2 = 0;

// Input weights (h×d for each gate)
logic signed [WIDTH-1:0] w_ir_0_0 = 'b000000011;
logic signed [WIDTH-1:0] w_ir_0_1 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_0_2 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_3 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_0_4 = 'b111111110;
logic signed [WIDTH-1:0] w_ir_1_0 = 'b111111011;
logic signed [WIDTH-1:0] w_ir_1_1 = 'b000000100;
logic signed [WIDTH-1:0] w_ir_1_2 = 'b000000010;
logic signed [WIDTH-1:0] w_ir_1_3 = 'b111111001;
logic signed [WIDTH-1:0] w_ir_1_4 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_0 = 'b000001000;
logic signed [WIDTH-1:0] w_ir_2_1 = 'b000000000;
logic signed [WIDTH-1:0] w_ir_2_2 = 'b000000101;
logic signed [WIDTH-1:0] w_ir_2_3 = 'b000000001;
logic signed [WIDTH-1:0] w_ir_2_4 = 'b000000001;

logic signed [WIDTH-1:0] w_iz_0_0 = 'b000000110;
logic signed [WIDTH-1:0] w_iz_0_1 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_2 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_0_3 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_0_4 = 'b000000101;
logic signed [WIDTH-1:0] w_iz_1_0 = 'b111111111;
logic signed [WIDTH-1:0] w_iz_1_1 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_1_2 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_1_3 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_1_4 = 'b111111011;
logic signed [WIDTH-1:0] w_iz_2_0 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_2_1 = 'b000000100;
logic signed [WIDTH-1:0] w_iz_2_2 = 'b000000011;
logic signed [WIDTH-1:0] w_iz_2_3 = 'b000000111;
logic signed [WIDTH-1:0] w_iz_2_4 = 'b111111001;

logic signed [WIDTH-1:0] w_in_0_0 = 'b111111110;
logic signed [WIDTH-1:0] w_in_0_1 = 'b000000011;
logic signed [WIDTH-1:0] w_in_0_2 = 'b000000010;
logic signed [WIDTH-1:0] w_in_0_3 = 'b000000100;
logic signed [WIDTH-1:0] w_in_0_4 = 'b000000100;
logic signed [WIDTH-1:0] w_in_1_0 = 'b000000001;
logic signed [WIDTH-1:0] w_in_1_1 = 'b000001000;
logic signed [WIDTH-1:0] w_in_1_2 = 'b000000011;
logic signed [WIDTH-1:0] w_in_1_3 = 'b111111110;
logic signed [WIDTH-1:0] w_in_1_4 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_0 = 'b000000101;
logic signed [WIDTH-1:0] w_in_2_1 = 'b111111010;
logic signed [WIDTH-1:0] w_in_2_2 = 'b000000010;
logic signed [WIDTH-1:0] w_in_2_3 = 'b111111101;
logic signed [WIDTH-1:0] w_in_2_4 = 'b000000000;

// Recurrent weights (h×h for each gate)
logic signed [WIDTH-1:0] w_hr_0_0 = 'b000000000;
logic signed [WIDTH-1:0] w_hr_0_1 = 'b000000001;
logic signed [WIDTH-1:0] w_hr_0_2 = 'b000000010;
logic signed [WIDTH-1:0] w_hr_1_0 = 'b111111011;
logic signed [WIDTH-1:0] w_hr_1_1 = 'b000001001;
logic signed [WIDTH-1:0] w_hr_1_2 = 'b000001001;
logic signed [WIDTH-1:0] w_hr_2_0 = 'b000001001;
logic signed [WIDTH-1:0] w_hr_2_1 = 'b111110111;
logic signed [WIDTH-1:0] w_hr_2_2 = 'b000001000;

logic signed [WIDTH-1:0] w_hz_0_0 = 'b000001001;
logic signed [WIDTH-1:0] w_hz_0_1 = 'b111111100;
logic signed [WIDTH-1:0] w_hz_0_2 = 'b111111011;
logic signed [WIDTH-1:0] w_hz_1_0 = 'b000000100;
logic signed [WIDTH-1:0] w_hz_1_1 = 'b000000101;
logic signed [WIDTH-1:0] w_hz_1_2 = 'b000001011;
logic signed [WIDTH-1:0] w_hz_2_0 = 'b111111000;
logic signed [WIDTH-1:0] w_hz_2_1 = 'b000000111;
logic signed [WIDTH-1:0] w_hz_2_2 = 'b000000100;

logic signed [WIDTH-1:0] w_hn_0_0 = 'b111111101;
logic signed [WIDTH-1:0] w_hn_0_1 = 'b000000100;
logic signed [WIDTH-1:0] w_hn_0_2 = 'b000001101;
logic signed [WIDTH-1:0] w_hn_1_0 = 'b111110100;
logic signed [WIDTH-1:0] w_hn_1_1 = 'b000000000;
logic signed [WIDTH-1:0] w_hn_1_2 = 'b000001001;
logic signed [WIDTH-1:0] w_hn_2_0 = 'b000000111;
logic signed [WIDTH-1:0] w_hn_2_1 = 'b000000000;
logic signed [WIDTH-1:0] w_hn_2_2 = 'b111110000;

// Biases (h for each gate type)
logic signed [WIDTH-1:0] b_ir_0 = 'b000000001;
logic signed [WIDTH-1:0] b_ir_1 = 'b000001000;
logic signed [WIDTH-1:0] b_ir_2 = 'b000001111;

logic signed [WIDTH-1:0] b_iz_0 = 'b000000101;
logic signed [WIDTH-1:0] b_iz_1 = 'b000000110;
logic signed [WIDTH-1:0] b_iz_2 = 'b000000100;

logic signed [WIDTH-1:0] b_in_0 = 'b000010000;
logic signed [WIDTH-1:0] b_in_1 = 'b000000000;
logic signed [WIDTH-1:0] b_in_2 = 'b000001011;

logic signed [WIDTH-1:0] b_hr_0 = 'b000000010;
logic signed [WIDTH-1:0] b_hr_1 = 'b000001110;
logic signed [WIDTH-1:0] b_hr_2 = 'b000000010;

logic signed [WIDTH-1:0] b_hz_0 = 'b000000010;
logic signed [WIDTH-1:0] b_hz_1 = 'b000001010;
logic signed [WIDTH-1:0] b_hz_2 = 'b000000111;

logic signed [WIDTH-1:0] b_hn_0 = 'b000001101;
logic signed [WIDTH-1:0] b_hn_1 = 'b000000111;
logic signed [WIDTH-1:0] b_hn_2 = 'b000001001;

// Outputs (h=3)
logic signed [WIDTH-1:0]  y_0 = 0;
logic signed [WIDTH-1:0]  y_1 = 0;
logic signed [WIDTH-1:0]  y_2 = 0;

gru #(
        .INT_WIDTH(INT_WIDTH),
        .FRAC_WIDTH(FRAC_WIDTH)
    ) gru_inst (
        .clk(clk),
        .reset(reset),
        // Input features (d=64)
        	
.x_0(x_0), .x_1(x_1), .x_2(x_2), .x_3(x_3), .x_4(x_4), 	
.h_0(h_0), .h_1(h_1), .h_2(h_2), 	
.w_ir_0_0(w_ir_0_0), .w_ir_0_1(w_ir_0_1), .w_ir_0_2(w_ir_0_2), .w_ir_0_3(w_ir_0_3), .w_ir_0_4(w_ir_0_4), .w_ir_1_0(w_ir_1_0), .w_ir_1_1(w_ir_1_1), .w_ir_1_2(w_ir_1_2), .w_ir_1_3(w_ir_1_3), .w_ir_1_4(w_ir_1_4), .w_ir_2_0(w_ir_2_0), .w_ir_2_1(w_ir_2_1), .w_ir_2_2(w_ir_2_2), .w_ir_2_3(w_ir_2_3), .w_ir_2_4(w_ir_2_4), 	
.w_iz_0_0(w_iz_0_0), .w_iz_0_1(w_iz_0_1), .w_iz_0_2(w_iz_0_2), .w_iz_0_3(w_iz_0_3), .w_iz_0_4(w_iz_0_4), .w_iz_1_0(w_iz_1_0), .w_iz_1_1(w_iz_1_1), .w_iz_1_2(w_iz_1_2), .w_iz_1_3(w_iz_1_3), .w_iz_1_4(w_iz_1_4), .w_iz_2_0(w_iz_2_0), .w_iz_2_1(w_iz_2_1), .w_iz_2_2(w_iz_2_2), .w_iz_2_3(w_iz_2_3), .w_iz_2_4(w_iz_2_4), 
.w_in_0_0(w_in_0_0), .w_in_0_1(w_in_0_1), .w_in_0_2(w_in_0_2), .w_in_0_3(w_in_0_3), .w_in_0_4(w_in_0_4), .w_in_1_0(w_in_1_0), .w_in_1_1(w_in_1_1), .w_in_1_2(w_in_1_2), .w_in_1_3(w_in_1_3), .w_in_1_4(w_in_1_4), .w_in_2_0(w_in_2_0), .w_in_2_1(w_in_2_1), .w_in_2_2(w_in_2_2), .w_in_2_3(w_in_2_3), .w_in_2_4(w_in_2_4), 
.w_hr_0_0(w_hr_0_0), .w_hr_0_1(w_hr_0_1), .w_hr_0_2(w_hr_0_2), .w_hr_1_0(w_hr_1_0), .w_hr_1_1(w_hr_1_1), .w_hr_1_2(w_hr_1_2), .w_hr_2_0(w_hr_2_0), .w_hr_2_1(w_hr_2_1), .w_hr_2_2(w_hr_2_2), 
.w_hz_0_0(w_hz_0_0), .w_hz_0_1(w_hz_0_1), .w_hz_0_2(w_hz_0_2), .w_hz_1_0(w_hz_1_0), .w_hz_1_1(w_hz_1_1), .w_hz_1_2(w_hz_1_2), .w_hz_2_0(w_hz_2_0), .w_hz_2_1(w_hz_2_1), .w_hz_2_2(w_hz_2_2), 
.w_hn_0_0(w_hn_0_0), .w_hn_0_1(w_hn_0_1), .w_hn_0_2(w_hn_0_2), .w_hn_1_0(w_hn_1_0), .w_hn_1_1(w_hn_1_1), .w_hn_1_2(w_hn_1_2), .w_hn_2_0(w_hn_2_0), .w_hn_2_1(w_hn_2_1), .w_hn_2_2(w_hn_2_2), 
.b_ir_0(b_ir_0), .b_ir_1(b_ir_1), .b_ir_2(b_ir_2), 
.b_iz_0(b_iz_0), .b_iz_1(b_iz_1), .b_iz_2(b_iz_2), 
.b_in_0(b_in_0), .b_in_1(b_in_1), .b_in_2(b_in_2), 
.b_hr_0(b_hr_0), .b_hr_1(b_hr_1), .b_hr_2(b_hr_2), 
.b_hz_0(b_hz_0), .b_hz_1(b_hz_1), .b_hz_2(b_hz_2), 
.b_hn_0(b_hn_0), .b_hn_1(b_hn_1), .b_hn_2(b_hn_2), 
.y_0(y_0), .y_1(y_1), .y_2(y_2)
);

    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end
    
    initial begin
        // Open file for writing (overwrite existing)
        integer fd;
        fd = $fopen("../../../../../output_d5_h3_int4_frac5.txt", "w+");
        if (fd == 0) begin
            $display("ERROR: Failed to open file!");
            $finish;
        end
        x_0 = 'b000100100;
    x_1 = 'b000110111;
    x_2 = 'b001000001;
    x_3 = 'b001001001;
    x_4 = 'b000111011;

    h_0 = 'b000100100;
    h_1 = 'b000110111;
    h_2 = 'b001000001;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000101110;
    x_1 = 'b001001001;
    x_2 = 'b001010010;
    x_3 = 'b001010101;
    x_4 = 'b001001111;

    h_0 = 'b000101110;
    h_1 = 'b001001001;
    h_2 = 'b001010010;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000111111;
    x_1 = 'b001000011;
    x_2 = 'b001000001;
    x_3 = 'b001000000;
    x_4 = 'b000110111;

    h_0 = 'b000111111;
    h_1 = 'b001000011;
    h_2 = 'b001000001;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000101101;
    x_1 = 'b000101111;
    x_2 = 'b000110100;
    x_3 = 'b000111010;
    x_4 = 'b000110001;

    h_0 = 'b000101101;
    h_1 = 'b000101111;
    h_2 = 'b000110100;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000011100;
    x_1 = 'b000100110;
    x_2 = 'b000101001;
    x_3 = 'b000110001;
    x_4 = 'b000101100;

    h_0 = 'b000011100;
    h_1 = 'b000100110;
    h_2 = 'b000101001;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000010011;
    x_1 = 'b000011111;
    x_2 = 'b000100100;
    x_3 = 'b000101100;
    x_4 = 'b000100101;

    h_0 = 'b000010011;
    h_1 = 'b000011111;
    h_2 = 'b000100100;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000011001;
    x_1 = 'b000100101;
    x_2 = 'b000101100;
    x_3 = 'b000110101;
    x_4 = 'b000101111;

    h_0 = 'b000011001;
    h_1 = 'b000100101;
    h_2 = 'b000101100;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000011001;
    x_1 = 'b000100011;
    x_2 = 'b000101001;
    x_3 = 'b000110101;
    x_4 = 'b000110001;

    h_0 = 'b000011001;
    h_1 = 'b000100011;
    h_2 = 'b000101001;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000010111;
    x_1 = 'b000011110;
    x_2 = 'b000100110;
    x_3 = 'b000101111;
    x_4 = 'b000101011;

    h_0 = 'b000010111;
    h_1 = 'b000011110;
    h_2 = 'b000100110;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000010001;
    x_1 = 'b000010011;
    x_2 = 'b000011010;
    x_3 = 'b000100010;
    x_4 = 'b000011111;

    h_0 = 'b000010001;
    h_1 = 'b000010011;
    h_2 = 'b000011010;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000000110;
    x_1 = 'b000000111;
    x_2 = 'b000001011;
    x_3 = 'b000010001;
    x_4 = 'b000001101;

    h_0 = 'b000000110;
    h_1 = 'b000000111;
    h_2 = 'b000001011;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000010101;
    x_1 = 'b000010000;
    x_2 = 'b000010000;
    x_3 = 'b000010001;
    x_4 = 'b000001101;

    h_0 = 'b000010101;
    h_1 = 'b000010000;
    h_2 = 'b000010000;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000010101;
    x_1 = 'b000010010;
    x_2 = 'b000010001;
    x_3 = 'b000010010;
    x_4 = 'b000001010;

    h_0 = 'b000010101;
    h_1 = 'b000010010;
    h_2 = 'b000010001;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000001111;
    x_1 = 'b000000110;
    x_2 = 'b000001000;
    x_3 = 'b000001101;
    x_4 = 'b111111110;

    h_0 = 'b000001111;
    h_1 = 'b000000110;
    h_2 = 'b000001000;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000010100;
    x_1 = 'b000001011;
    x_2 = 'b000001011;
    x_3 = 'b000001110;
    x_4 = 'b000000001;

    h_0 = 'b000010100;
    h_1 = 'b000001011;
    h_2 = 'b000001011;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000011010;
    x_1 = 'b000011001;
    x_2 = 'b000011100;
    x_3 = 'b000100000;
    x_4 = 'b000011001;

    h_0 = 'b000011010;
    h_1 = 'b000011001;
    h_2 = 'b000011100;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000000101;
    x_1 = 'b000000111;
    x_2 = 'b111101000;
    x_3 = 'b111110000;
    x_4 = 'b111101101;

    h_0 = 'b000000101;
    h_1 = 'b000000111;
    h_2 = 'b111101000;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000010101;
    x_1 = 'b000011000;
    x_2 = 'b000000000;
    x_3 = 'b000000101;
    x_4 = 'b111111101;

    h_0 = 'b000010101;
    h_1 = 'b000011000;
    h_2 = 'b000000000;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000100101;
    x_1 = 'b000100001;
    x_2 = 'b000001010;
    x_3 = 'b000001011;
    x_4 = 'b000000001;

    h_0 = 'b000100101;
    h_1 = 'b000100001;
    h_2 = 'b000001010;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000111001;
    x_1 = 'b000110110;
    x_2 = 'b000011111;
    x_3 = 'b000011100;
    x_4 = 'b000010111;

    h_0 = 'b000111001;
    h_1 = 'b000110110;
    h_2 = 'b000011111;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000010111;
    x_1 = 'b000011001;
    x_2 = 'b000001000;
    x_3 = 'b000001001;
    x_4 = 'b000001101;

    h_0 = 'b000010111;
    h_1 = 'b000011001;
    h_2 = 'b000001000;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000000110;
    x_1 = 'b000001011;
    x_2 = 'b111111101;
    x_3 = 'b000000010;
    x_4 = 'b000001001;

    h_0 = 'b000000110;
    h_1 = 'b000001011;
    h_2 = 'b111111101;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000100110;
    x_1 = 'b000100001;
    x_2 = 'b000001011;
    x_3 = 'b000010001;
    x_4 = 'b000001101;

    h_0 = 'b000100110;
    h_1 = 'b000100001;
    h_2 = 'b000001011;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000001001;
    x_1 = 'b000001110;
    x_2 = 'b111111111;
    x_3 = 'b000000111;
    x_4 = 'b111111111;

    h_0 = 'b000001001;
    h_1 = 'b000001110;
    h_2 = 'b111111111;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000001001;
    x_1 = 'b000010010;
    x_2 = 'b000000100;
    x_3 = 'b000001010;
    x_4 = 'b000000000;

    h_0 = 'b000001001;
    h_1 = 'b000010010;
    h_2 = 'b000000100;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000001010;
    x_1 = 'b000011001;
    x_2 = 'b000001110;
    x_3 = 'b000010110;
    x_4 = 'b000001010;

    h_0 = 'b000001010;
    h_1 = 'b000011001;
    h_2 = 'b000001110;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111111010;
    x_1 = 'b000000110;
    x_2 = 'b000000001;
    x_3 = 'b000001001;
    x_4 = 'b000000000;

    h_0 = 'b111111010;
    h_1 = 'b000000110;
    h_2 = 'b000000001;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000001001;
    x_1 = 'b000001001;
    x_2 = 'b111111110;
    x_3 = 'b000000001;
    x_4 = 'b111111000;

    h_0 = 'b000001001;
    h_1 = 'b000001001;
    h_2 = 'b111111110;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000001010;
    x_1 = 'b000001010;
    x_2 = 'b111111011;
    x_3 = 'b111111101;
    x_4 = 'b111110000;

    h_0 = 'b000001010;
    h_1 = 'b000001010;
    h_2 = 'b111111011;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000011000;
    x_1 = 'b000011100;
    x_2 = 'b000001101;
    x_3 = 'b000001111;
    x_4 = 'b000000111;

    h_0 = 'b000011000;
    h_1 = 'b000011100;
    h_2 = 'b000001101;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000011111;
    x_1 = 'b000100000;
    x_2 = 'b000001110;
    x_3 = 'b000010111;
    x_4 = 'b000001011;

    h_0 = 'b000011111;
    h_1 = 'b000100000;
    h_2 = 'b000001110;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000001100;
    x_1 = 'b000010101;
    x_2 = 'b111111110;
    x_3 = 'b000010010;
    x_4 = 'b000000110;

    h_0 = 'b000001100;
    h_1 = 'b000010101;
    h_2 = 'b111111110;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111110101;
    x_1 = 'b111110101;
    x_2 = 'b111110000;
    x_3 = 'b111110001;
    x_4 = 'b111101100;

    h_0 = 'b111110101;
    h_1 = 'b111110101;
    h_2 = 'b111110000;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111100100;
    x_1 = 'b111100100;
    x_2 = 'b111011111;
    x_3 = 'b111011101;
    x_4 = 'b111011011;

    h_0 = 'b111100100;
    h_1 = 'b111100100;
    h_2 = 'b111011111;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111100010;
    x_1 = 'b111100001;
    x_2 = 'b111011011;
    x_3 = 'b111011101;
    x_4 = 'b111011011;

    h_0 = 'b111100010;
    h_1 = 'b111100001;
    h_2 = 'b111011011;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111101101;
    x_1 = 'b111110101;
    x_2 = 'b111110011;
    x_3 = 'b111110100;
    x_4 = 'b111110011;

    h_0 = 'b111101101;
    h_1 = 'b111110101;
    h_2 = 'b111110011;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111111100;
    x_1 = 'b000000110;
    x_2 = 'b111111111;
    x_3 = 'b111111100;
    x_4 = 'b111111000;

    h_0 = 'b111111100;
    h_1 = 'b000000110;
    h_2 = 'b111111111;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000000010;
    x_1 = 'b000000010;
    x_2 = 'b111111001;
    x_3 = 'b111110010;
    x_4 = 'b111101110;

    h_0 = 'b000000010;
    h_1 = 'b000000010;
    h_2 = 'b111111001;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000010011;
    x_1 = 'b000010010;
    x_2 = 'b000000110;
    x_3 = 'b111111101;
    x_4 = 'b111111000;

    h_0 = 'b000010011;
    h_1 = 'b000010010;
    h_2 = 'b000000110;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000001111;
    x_1 = 'b000010011;
    x_2 = 'b000000110;
    x_3 = 'b000000001;
    x_4 = 'b111111011;

    h_0 = 'b000001111;
    h_1 = 'b000010011;
    h_2 = 'b000000110;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000000011;
    x_1 = 'b000001001;
    x_2 = 'b000000010;
    x_3 = 'b111111101;
    x_4 = 'b111111001;

    h_0 = 'b000000011;
    h_1 = 'b000001001;
    h_2 = 'b000000010;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000010001;
    x_1 = 'b000011101;
    x_2 = 'b000010111;
    x_3 = 'b000010011;
    x_4 = 'b000001011;

    h_0 = 'b000010001;
    h_1 = 'b000011101;
    h_2 = 'b000010111;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000010110;
    x_1 = 'b000011011;
    x_2 = 'b000010101;
    x_3 = 'b000010101;
    x_4 = 'b000001110;

    h_0 = 'b000010110;
    h_1 = 'b000011011;
    h_2 = 'b000010101;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000010100;
    x_1 = 'b000010101;
    x_2 = 'b000001110;
    x_3 = 'b000001111;
    x_4 = 'b000001001;

    h_0 = 'b000010100;
    h_1 = 'b000010101;
    h_2 = 'b000001110;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000011100;
    x_1 = 'b000100000;
    x_2 = 'b000011100;
    x_3 = 'b000011010;
    x_4 = 'b000010011;

    h_0 = 'b000011100;
    h_1 = 'b000100000;
    h_2 = 'b000011100;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000011010;
    x_1 = 'b000100001;
    x_2 = 'b000011010;
    x_3 = 'b000010111;
    x_4 = 'b000010000;

    h_0 = 'b000011010;
    h_1 = 'b000100001;
    h_2 = 'b000011010;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000100110;
    x_1 = 'b000101100;
    x_2 = 'b000100011;
    x_3 = 'b000100100;
    x_4 = 'b000011010;

    h_0 = 'b000100110;
    h_1 = 'b000101100;
    h_2 = 'b000100011;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000010101;
    x_1 = 'b000011100;
    x_2 = 'b000011001;
    x_3 = 'b000100000;
    x_4 = 'b000011001;

    h_0 = 'b000010101;
    h_1 = 'b000011100;
    h_2 = 'b000011001;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111100111;
    x_1 = 'b111011000;
    x_2 = 'b111000111;
    x_3 = 'b110111000;
    x_4 = 'b110111100;

    h_0 = 'b111100111;
    h_1 = 'b111011000;
    h_2 = 'b111000111;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111010111;
    x_1 = 'b111001010;
    x_2 = 'b110110101;
    x_3 = 'b110100100;
    x_4 = 'b110100100;

    h_0 = 'b111010111;
    h_1 = 'b111001010;
    h_2 = 'b110110101;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111011001;
    x_1 = 'b111001001;
    x_2 = 'b110111001;
    x_3 = 'b110101010;
    x_4 = 'b110101001;

    h_0 = 'b111011001;
    h_1 = 'b111001001;
    h_2 = 'b110111001;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111101101;
    x_1 = 'b111100001;
    x_2 = 'b111010000;
    x_3 = 'b111000000;
    x_4 = 'b111000000;

    h_0 = 'b111101101;
    h_1 = 'b111100001;
    h_2 = 'b111010000;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111111101;
    x_1 = 'b111110000;
    x_2 = 'b111100001;
    x_3 = 'b111010110;
    x_4 = 'b111010110;

    h_0 = 'b111111101;
    h_1 = 'b111110000;
    h_2 = 'b111100001;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111111011;
    x_1 = 'b111101111;
    x_2 = 'b111100010;
    x_3 = 'b111011010;
    x_4 = 'b111011001;

    h_0 = 'b111111011;
    h_1 = 'b111101111;
    h_2 = 'b111100010;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111111010;
    x_1 = 'b111101100;
    x_2 = 'b111011100;
    x_3 = 'b111010001;
    x_4 = 'b111010001;

    h_0 = 'b111111010;
    h_1 = 'b111101100;
    h_2 = 'b111011100;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111110111;
    x_1 = 'b111100111;
    x_2 = 'b111010110;
    x_3 = 'b111001110;
    x_4 = 'b111001101;

    h_0 = 'b111110111;
    h_1 = 'b111100111;
    h_2 = 'b111010110;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111110110;
    x_1 = 'b111011111;
    x_2 = 'b111010000;
    x_3 = 'b111000111;
    x_4 = 'b111001000;

    h_0 = 'b111110110;
    h_1 = 'b111011111;
    h_2 = 'b111010000;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111101111;
    x_1 = 'b111011011;
    x_2 = 'b111001101;
    x_3 = 'b111000011;
    x_4 = 'b111001000;

    h_0 = 'b111101111;
    h_1 = 'b111011011;
    h_2 = 'b111001101;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111101110;
    x_1 = 'b111100000;
    x_2 = 'b111001101;
    x_3 = 'b111000011;
    x_4 = 'b111000110;

    h_0 = 'b111101110;
    h_1 = 'b111100000;
    h_2 = 'b111001101;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111111101;
    x_1 = 'b111110000;
    x_2 = 'b111011010;
    x_3 = 'b111001111;
    x_4 = 'b111001011;

    h_0 = 'b111111101;
    h_1 = 'b111110000;
    h_2 = 'b111011010;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111111101;
    x_1 = 'b111101011;
    x_2 = 'b111010111;
    x_3 = 'b111001010;
    x_4 = 'b111000101;

    h_0 = 'b111111101;
    h_1 = 'b111101011;
    h_2 = 'b111010111;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000000101;
    x_1 = 'b111110010;
    x_2 = 'b111011100;
    x_3 = 'b111000110;
    x_4 = 'b111000100;

    h_0 = 'b000000101;
    h_1 = 'b111110010;
    h_2 = 'b111011100;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000000001;
    x_1 = 'b111110111;
    x_2 = 'b111100001;
    x_3 = 'b111001011;
    x_4 = 'b111000001;

    h_0 = 'b000000001;
    h_1 = 'b111110111;
    h_2 = 'b111100001;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000000111;
    x_1 = 'b111111011;
    x_2 = 'b111100100;
    x_3 = 'b111001111;
    x_4 = 'b111000111;

    h_0 = 'b000000111;
    h_1 = 'b111111011;
    h_2 = 'b111100100;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111001010;
    x_1 = 'b111011110;
    x_2 = 'b111100001;
    x_3 = 'b111110101;
    x_4 = 'b111111001;

    h_0 = 'b111001010;
    h_1 = 'b111011110;
    h_2 = 'b111100001;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111001110;
    x_1 = 'b111100100;
    x_2 = 'b111100111;
    x_3 = 'b111110101;
    x_4 = 'b111111011;

    h_0 = 'b111001110;
    h_1 = 'b111100100;
    h_2 = 'b111100111;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111010101;
    x_1 = 'b111101011;
    x_2 = 'b111101011;
    x_3 = 'b111110100;
    x_4 = 'b111111001;

    h_0 = 'b111010101;
    h_1 = 'b111101011;
    h_2 = 'b111101011;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111100010;
    x_1 = 'b111110010;
    x_2 = 'b111101111;
    x_3 = 'b111110101;
    x_4 = 'b111111000;

    h_0 = 'b111100010;
    h_1 = 'b111110010;
    h_2 = 'b111101111;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111011111;
    x_1 = 'b111101111;
    x_2 = 'b111101110;
    x_3 = 'b111110101;
    x_4 = 'b111110111;

    h_0 = 'b111011111;
    h_1 = 'b111101111;
    h_2 = 'b111101110;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111100000;
    x_1 = 'b111110000;
    x_2 = 'b111110100;
    x_3 = 'b111111110;
    x_4 = 'b000000010;

    h_0 = 'b111100000;
    h_1 = 'b111110000;
    h_2 = 'b111110100;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111010001;
    x_1 = 'b111100100;
    x_2 = 'b111100111;
    x_3 = 'b111110111;
    x_4 = 'b111111011;

    h_0 = 'b111010001;
    h_1 = 'b111100100;
    h_2 = 'b111100111;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111010101;
    x_1 = 'b111101010;
    x_2 = 'b111101010;
    x_3 = 'b111111011;
    x_4 = 'b000000100;

    h_0 = 'b111010101;
    h_1 = 'b111101010;
    h_2 = 'b111101010;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111100100;
    x_1 = 'b111110010;
    x_2 = 'b111110000;
    x_3 = 'b000000000;
    x_4 = 'b000000110;

    h_0 = 'b111100100;
    h_1 = 'b111110010;
    h_2 = 'b111110000;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111100111;
    x_1 = 'b111111000;
    x_2 = 'b111110011;
    x_3 = 'b000000010;
    x_4 = 'b000000010;

    h_0 = 'b111100111;
    h_1 = 'b111111000;
    h_2 = 'b111110011;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111100100;
    x_1 = 'b111111010;
    x_2 = 'b111110100;
    x_3 = 'b000000010;
    x_4 = 'b000000001;

    h_0 = 'b111100100;
    h_1 = 'b111111010;
    h_2 = 'b111110100;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111011101;
    x_1 = 'b111101000;
    x_2 = 'b111100111;
    x_3 = 'b111110111;
    x_4 = 'b111110110;

    h_0 = 'b111011101;
    h_1 = 'b111101000;
    h_2 = 'b111100111;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111110001;
    x_1 = 'b111111011;
    x_2 = 'b111111000;
    x_3 = 'b000000111;
    x_4 = 'b000000110;

    h_0 = 'b111110001;
    h_1 = 'b111111011;
    h_2 = 'b111111000;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111110101;
    x_1 = 'b111111011;
    x_2 = 'b111110100;
    x_3 = 'b111111111;
    x_4 = 'b111111101;

    h_0 = 'b111110101;
    h_1 = 'b111111011;
    h_2 = 'b111110100;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111101001;
    x_1 = 'b111110010;
    x_2 = 'b111101101;
    x_3 = 'b111110100;
    x_4 = 'b111110101;

    h_0 = 'b111101001;
    h_1 = 'b111110010;
    h_2 = 'b111101101;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111101011;
    x_1 = 'b111110110;
    x_2 = 'b111110100;
    x_3 = 'b111111101;
    x_4 = 'b111111111;

    h_0 = 'b111101011;
    h_1 = 'b111110110;
    h_2 = 'b111110100;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000001110;
    x_1 = 'b000001110;
    x_2 = 'b000000110;
    x_3 = 'b000001100;
    x_4 = 'b000010000;

    h_0 = 'b000001110;
    h_1 = 'b000001110;
    h_2 = 'b000000110;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000000101;
    x_1 = 'b000000110;
    x_2 = 'b000000001;
    x_3 = 'b000001010;
    x_4 = 'b000001101;

    h_0 = 'b000000101;
    h_1 = 'b000000110;
    h_2 = 'b000000001;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111111011;
    x_1 = 'b000000000;
    x_2 = 'b000000000;
    x_3 = 'b000001100;
    x_4 = 'b000001110;

    h_0 = 'b111111011;
    h_1 = 'b000000000;
    h_2 = 'b000000000;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111101101;
    x_1 = 'b111110011;
    x_2 = 'b111110010;
    x_3 = 'b111111100;
    x_4 = 'b111111110;

    h_0 = 'b111101101;
    h_1 = 'b111110011;
    h_2 = 'b111110010;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111110101;
    x_1 = 'b111111010;
    x_2 = 'b111110000;
    x_3 = 'b111110110;
    x_4 = 'b111110110;

    h_0 = 'b111110101;
    h_1 = 'b111111010;
    h_2 = 'b111110000;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111110101;
    x_1 = 'b111111010;
    x_2 = 'b111110011;
    x_3 = 'b111110101;
    x_4 = 'b111111010;

    h_0 = 'b111110101;
    h_1 = 'b111111010;
    h_2 = 'b111110011;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000000001;
    x_1 = 'b000000011;
    x_2 = 'b111111010;
    x_3 = 'b111111011;
    x_4 = 'b000000010;

    h_0 = 'b000000001;
    h_1 = 'b000000011;
    h_2 = 'b111111010;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000001000;
    x_1 = 'b000001000;
    x_2 = 'b111111111;
    x_3 = 'b000000000;
    x_4 = 'b000000100;

    h_0 = 'b000001000;
    h_1 = 'b000001000;
    h_2 = 'b111111111;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000001011;
    x_1 = 'b000001001;
    x_2 = 'b000000001;
    x_3 = 'b000000110;
    x_4 = 'b000001001;

    h_0 = 'b000001011;
    h_1 = 'b000001001;
    h_2 = 'b000000001;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000001110;
    x_1 = 'b000001110;
    x_2 = 'b000001001;
    x_3 = 'b000001111;
    x_4 = 'b000010101;

    h_0 = 'b000001110;
    h_1 = 'b000001110;
    h_2 = 'b000001001;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000001001;
    x_1 = 'b000010010;
    x_2 = 'b000010101;
    x_3 = 'b000011101;
    x_4 = 'b000011101;

    h_0 = 'b000001001;
    h_1 = 'b000010010;
    h_2 = 'b000010101;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000001110;
    x_1 = 'b000011011;
    x_2 = 'b000011111;
    x_3 = 'b000100101;
    x_4 = 'b000100001;

    h_0 = 'b000001110;
    h_1 = 'b000011011;
    h_2 = 'b000011111;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000011010;
    x_1 = 'b000100110;
    x_2 = 'b000100111;
    x_3 = 'b000101011;
    x_4 = 'b000100111;

    h_0 = 'b000011010;
    h_1 = 'b000100110;
    h_2 = 'b000100111;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000100100;
    x_1 = 'b000101111;
    x_2 = 'b000101111;
    x_3 = 'b000110001;
    x_4 = 'b000101110;

    h_0 = 'b000100100;
    h_1 = 'b000101111;
    h_2 = 'b000101111;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000010010;
    x_1 = 'b000011010;
    x_2 = 'b000010110;
    x_3 = 'b000010101;
    x_4 = 'b000010001;

    h_0 = 'b000010010;
    h_1 = 'b000011010;
    h_2 = 'b000010110;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000001001;
    x_1 = 'b000010000;
    x_2 = 'b000001011;
    x_3 = 'b000001011;
    x_4 = 'b000000110;

    h_0 = 'b000001001;
    h_1 = 'b000010000;
    h_2 = 'b000001011;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111111001;
    x_1 = 'b111111001;
    x_2 = 'b111101111;
    x_3 = 'b111110101;
    x_4 = 'b111111000;

    h_0 = 'b111111001;
    h_1 = 'b111111001;
    h_2 = 'b111101111;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b000000001;
    x_1 = 'b000000000;
    x_2 = 'b111110101;
    x_3 = 'b111111101;
    x_4 = 'b111111100;

    h_0 = 'b000000001;
    h_1 = 'b000000000;
    h_2 = 'b111110101;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111110111;
    x_1 = 'b111110101;
    x_2 = 'b111101100;
    x_3 = 'b111110100;
    x_4 = 'b111110011;

    h_0 = 'b111110111;
    h_1 = 'b111110101;
    h_2 = 'b111101100;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    x_0 = 'b111110111;
    x_1 = 'b111110010;
    x_2 = 'b111100101;
    x_3 = 'b111101111;
    x_4 = 'b111101111;

    h_0 = 'b111110111;
    h_1 = 'b111110010;
    h_2 = 'b111100101;
    #20;
    $fdisplay(fd, "%09b %09b %09b", y_0, y_1, y_2);

    $fclose(fd);    
$finish;
    end
endmodule